module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70,
        output wire [0:0] dst71);
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    reg [161:0] src16;
    reg [161:0] src17;
    reg [161:0] src18;
    reg [161:0] src19;
    reg [161:0] src20;
    reg [161:0] src21;
    reg [161:0] src22;
    reg [161:0] src23;
    reg [161:0] src24;
    reg [161:0] src25;
    reg [161:0] src26;
    reg [161:0] src27;
    reg [161:0] src28;
    reg [161:0] src29;
    reg [161:0] src30;
    reg [161:0] src31;
    reg [161:0] src32;
    reg [161:0] src33;
    reg [161:0] src34;
    reg [161:0] src35;
    reg [161:0] src36;
    reg [161:0] src37;
    reg [161:0] src38;
    reg [161:0] src39;
    reg [161:0] src40;
    reg [161:0] src41;
    reg [161:0] src42;
    reg [161:0] src43;
    reg [161:0] src44;
    reg [161:0] src45;
    reg [161:0] src46;
    reg [161:0] src47;
    reg [161:0] src48;
    reg [161:0] src49;
    reg [161:0] src50;
    reg [161:0] src51;
    reg [161:0] src52;
    reg [161:0] src53;
    reg [161:0] src54;
    reg [161:0] src55;
    reg [161:0] src56;
    reg [161:0] src57;
    reg [161:0] src58;
    reg [161:0] src59;
    reg [161:0] src60;
    reg [161:0] src61;
    reg [161:0] src62;
    reg [161:0] src63;
    compressor_CLA162_64 compressor_CLA162_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70),
            .dst71(dst71));
    initial begin
        src0 <= 162'h0;
        src1 <= 162'h0;
        src2 <= 162'h0;
        src3 <= 162'h0;
        src4 <= 162'h0;
        src5 <= 162'h0;
        src6 <= 162'h0;
        src7 <= 162'h0;
        src8 <= 162'h0;
        src9 <= 162'h0;
        src10 <= 162'h0;
        src11 <= 162'h0;
        src12 <= 162'h0;
        src13 <= 162'h0;
        src14 <= 162'h0;
        src15 <= 162'h0;
        src16 <= 162'h0;
        src17 <= 162'h0;
        src18 <= 162'h0;
        src19 <= 162'h0;
        src20 <= 162'h0;
        src21 <= 162'h0;
        src22 <= 162'h0;
        src23 <= 162'h0;
        src24 <= 162'h0;
        src25 <= 162'h0;
        src26 <= 162'h0;
        src27 <= 162'h0;
        src28 <= 162'h0;
        src29 <= 162'h0;
        src30 <= 162'h0;
        src31 <= 162'h0;
        src32 <= 162'h0;
        src33 <= 162'h0;
        src34 <= 162'h0;
        src35 <= 162'h0;
        src36 <= 162'h0;
        src37 <= 162'h0;
        src38 <= 162'h0;
        src39 <= 162'h0;
        src40 <= 162'h0;
        src41 <= 162'h0;
        src42 <= 162'h0;
        src43 <= 162'h0;
        src44 <= 162'h0;
        src45 <= 162'h0;
        src46 <= 162'h0;
        src47 <= 162'h0;
        src48 <= 162'h0;
        src49 <= 162'h0;
        src50 <= 162'h0;
        src51 <= 162'h0;
        src52 <= 162'h0;
        src53 <= 162'h0;
        src54 <= 162'h0;
        src55 <= 162'h0;
        src56 <= 162'h0;
        src57 <= 162'h0;
        src58 <= 162'h0;
        src59 <= 162'h0;
        src60 <= 162'h0;
        src61 <= 162'h0;
        src62 <= 162'h0;
        src63 <= 162'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA162_64(
    input [161:0]src0,
    input [161:0]src1,
    input [161:0]src2,
    input [161:0]src3,
    input [161:0]src4,
    input [161:0]src5,
    input [161:0]src6,
    input [161:0]src7,
    input [161:0]src8,
    input [161:0]src9,
    input [161:0]src10,
    input [161:0]src11,
    input [161:0]src12,
    input [161:0]src13,
    input [161:0]src14,
    input [161:0]src15,
    input [161:0]src16,
    input [161:0]src17,
    input [161:0]src18,
    input [161:0]src19,
    input [161:0]src20,
    input [161:0]src21,
    input [161:0]src22,
    input [161:0]src23,
    input [161:0]src24,
    input [161:0]src25,
    input [161:0]src26,
    input [161:0]src27,
    input [161:0]src28,
    input [161:0]src29,
    input [161:0]src30,
    input [161:0]src31,
    input [161:0]src32,
    input [161:0]src33,
    input [161:0]src34,
    input [161:0]src35,
    input [161:0]src36,
    input [161:0]src37,
    input [161:0]src38,
    input [161:0]src39,
    input [161:0]src40,
    input [161:0]src41,
    input [161:0]src42,
    input [161:0]src43,
    input [161:0]src44,
    input [161:0]src45,
    input [161:0]src46,
    input [161:0]src47,
    input [161:0]src48,
    input [161:0]src49,
    input [161:0]src50,
    input [161:0]src51,
    input [161:0]src52,
    input [161:0]src53,
    input [161:0]src54,
    input [161:0]src55,
    input [161:0]src56,
    input [161:0]src57,
    input [161:0]src58,
    input [161:0]src59,
    input [161:0]src60,
    input [161:0]src61,
    input [161:0]src62,
    input [161:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70,
    output dst71);

    wire [1:0] comp_out0;
    wire [0:0] comp_out1;
    wire [0:0] comp_out2;
    wire [0:0] comp_out3;
    wire [1:0] comp_out4;
    wire [0:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [0:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [0:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [0:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [1:0] comp_out69;
    wire [0:0] comp_out70;
    wire [0:0] comp_out71;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70),
        .dst71(comp_out71)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out71[0], comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out69[1], comp_out68[1], comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], 1'h0, comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], 1'h0, comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], 1'h0, comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], 1'h0, comp_out4[1], 1'h0, 1'h0, 1'h0, comp_out0[1]}),
        .dst({dst71, dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      input wire [161:0] src12,
      input wire [161:0] src13,
      input wire [161:0] src14,
      input wire [161:0] src15,
      input wire [161:0] src16,
      input wire [161:0] src17,
      input wire [161:0] src18,
      input wire [161:0] src19,
      input wire [161:0] src20,
      input wire [161:0] src21,
      input wire [161:0] src22,
      input wire [161:0] src23,
      input wire [161:0] src24,
      input wire [161:0] src25,
      input wire [161:0] src26,
      input wire [161:0] src27,
      input wire [161:0] src28,
      input wire [161:0] src29,
      input wire [161:0] src30,
      input wire [161:0] src31,
      input wire [161:0] src32,
      input wire [161:0] src33,
      input wire [161:0] src34,
      input wire [161:0] src35,
      input wire [161:0] src36,
      input wire [161:0] src37,
      input wire [161:0] src38,
      input wire [161:0] src39,
      input wire [161:0] src40,
      input wire [161:0] src41,
      input wire [161:0] src42,
      input wire [161:0] src43,
      input wire [161:0] src44,
      input wire [161:0] src45,
      input wire [161:0] src46,
      input wire [161:0] src47,
      input wire [161:0] src48,
      input wire [161:0] src49,
      input wire [161:0] src50,
      input wire [161:0] src51,
      input wire [161:0] src52,
      input wire [161:0] src53,
      input wire [161:0] src54,
      input wire [161:0] src55,
      input wire [161:0] src56,
      input wire [161:0] src57,
      input wire [161:0] src58,
      input wire [161:0] src59,
      input wire [161:0] src60,
      input wire [161:0] src61,
      input wire [161:0] src62,
      input wire [161:0] src63,
      output wire [1:0] dst0,
      output wire [0:0] dst1,
      output wire [0:0] dst2,
      output wire [0:0] dst3,
      output wire [1:0] dst4,
      output wire [0:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [0:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [0:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [0:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [1:0] dst69,
      output wire [0:0] dst70,
      output wire [0:0] dst71);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [161:0] stage0_12;
   wire [161:0] stage0_13;
   wire [161:0] stage0_14;
   wire [161:0] stage0_15;
   wire [161:0] stage0_16;
   wire [161:0] stage0_17;
   wire [161:0] stage0_18;
   wire [161:0] stage0_19;
   wire [161:0] stage0_20;
   wire [161:0] stage0_21;
   wire [161:0] stage0_22;
   wire [161:0] stage0_23;
   wire [161:0] stage0_24;
   wire [161:0] stage0_25;
   wire [161:0] stage0_26;
   wire [161:0] stage0_27;
   wire [161:0] stage0_28;
   wire [161:0] stage0_29;
   wire [161:0] stage0_30;
   wire [161:0] stage0_31;
   wire [161:0] stage0_32;
   wire [161:0] stage0_33;
   wire [161:0] stage0_34;
   wire [161:0] stage0_35;
   wire [161:0] stage0_36;
   wire [161:0] stage0_37;
   wire [161:0] stage0_38;
   wire [161:0] stage0_39;
   wire [161:0] stage0_40;
   wire [161:0] stage0_41;
   wire [161:0] stage0_42;
   wire [161:0] stage0_43;
   wire [161:0] stage0_44;
   wire [161:0] stage0_45;
   wire [161:0] stage0_46;
   wire [161:0] stage0_47;
   wire [161:0] stage0_48;
   wire [161:0] stage0_49;
   wire [161:0] stage0_50;
   wire [161:0] stage0_51;
   wire [161:0] stage0_52;
   wire [161:0] stage0_53;
   wire [161:0] stage0_54;
   wire [161:0] stage0_55;
   wire [161:0] stage0_56;
   wire [161:0] stage0_57;
   wire [161:0] stage0_58;
   wire [161:0] stage0_59;
   wire [161:0] stage0_60;
   wire [161:0] stage0_61;
   wire [161:0] stage0_62;
   wire [161:0] stage0_63;
   wire [33:0] stage1_0;
   wire [46:0] stage1_1;
   wire [54:0] stage1_2;
   wire [83:0] stage1_3;
   wire [82:0] stage1_4;
   wire [114:0] stage1_5;
   wire [57:0] stage1_6;
   wire [70:0] stage1_7;
   wire [80:0] stage1_8;
   wire [57:0] stage1_9;
   wire [94:0] stage1_10;
   wire [80:0] stage1_11;
   wire [66:0] stage1_12;
   wire [86:0] stage1_13;
   wire [61:0] stage1_14;
   wire [97:0] stage1_15;
   wire [67:0] stage1_16;
   wire [113:0] stage1_17;
   wire [62:0] stage1_18;
   wire [70:0] stage1_19;
   wire [67:0] stage1_20;
   wire [70:0] stage1_21;
   wire [66:0] stage1_22;
   wire [142:0] stage1_23;
   wire [82:0] stage1_24;
   wire [84:0] stage1_25;
   wire [71:0] stage1_26;
   wire [73:0] stage1_27;
   wire [76:0] stage1_28;
   wire [80:0] stage1_29;
   wire [106:0] stage1_30;
   wire [96:0] stage1_31;
   wire [86:0] stage1_32;
   wire [89:0] stage1_33;
   wire [55:0] stage1_34;
   wire [59:0] stage1_35;
   wire [82:0] stage1_36;
   wire [127:0] stage1_37;
   wire [65:0] stage1_38;
   wire [67:0] stage1_39;
   wire [81:0] stage1_40;
   wire [73:0] stage1_41;
   wire [95:0] stage1_42;
   wire [137:0] stage1_43;
   wire [45:0] stage1_44;
   wire [92:0] stage1_45;
   wire [63:0] stage1_46;
   wire [57:0] stage1_47;
   wire [71:0] stage1_48;
   wire [86:0] stage1_49;
   wire [57:0] stage1_50;
   wire [93:0] stage1_51;
   wire [76:0] stage1_52;
   wire [65:0] stage1_53;
   wire [57:0] stage1_54;
   wire [97:0] stage1_55;
   wire [79:0] stage1_56;
   wire [71:0] stage1_57;
   wire [73:0] stage1_58;
   wire [79:0] stage1_59;
   wire [66:0] stage1_60;
   wire [90:0] stage1_61;
   wire [86:0] stage1_62;
   wire [62:0] stage1_63;
   wire [44:0] stage1_64;
   wire [23:0] stage1_65;
   wire [9:0] stage2_0;
   wire [18:0] stage2_1;
   wire [37:0] stage2_2;
   wire [22:0] stage2_3;
   wire [47:0] stage2_4;
   wire [35:0] stage2_5;
   wire [28:0] stage2_6;
   wire [40:0] stage2_7;
   wire [60:0] stage2_8;
   wire [25:0] stage2_9;
   wire [40:0] stage2_10;
   wire [38:0] stage2_11;
   wire [30:0] stage2_12;
   wire [44:0] stage2_13;
   wire [73:0] stage2_14;
   wire [36:0] stage2_15;
   wire [46:0] stage2_16;
   wire [39:0] stage2_17;
   wire [42:0] stage2_18;
   wire [50:0] stage2_19;
   wire [57:0] stage2_20;
   wire [39:0] stage2_21;
   wire [30:0] stage2_22;
   wire [46:0] stage2_23;
   wire [45:0] stage2_24;
   wire [36:0] stage2_25;
   wire [52:0] stage2_26;
   wire [49:0] stage2_27;
   wire [34:0] stage2_28;
   wire [49:0] stage2_29;
   wire [49:0] stage2_30;
   wire [38:0] stage2_31;
   wire [55:0] stage2_32;
   wire [27:0] stage2_33;
   wire [34:0] stage2_34;
   wire [44:0] stage2_35;
   wire [36:0] stage2_36;
   wire [41:0] stage2_37;
   wire [32:0] stage2_38;
   wire [33:0] stage2_39;
   wire [40:0] stage2_40;
   wire [55:0] stage2_41;
   wire [61:0] stage2_42;
   wire [51:0] stage2_43;
   wire [65:0] stage2_44;
   wire [25:0] stage2_45;
   wire [32:0] stage2_46;
   wire [45:0] stage2_47;
   wire [23:0] stage2_48;
   wire [36:0] stage2_49;
   wire [40:0] stage2_50;
   wire [24:0] stage2_51;
   wire [33:0] stage2_52;
   wire [50:0] stage2_53;
   wire [27:0] stage2_54;
   wire [37:0] stage2_55;
   wire [52:0] stage2_56;
   wire [29:0] stage2_57;
   wire [32:0] stage2_58;
   wire [80:0] stage2_59;
   wire [21:0] stage2_60;
   wire [66:0] stage2_61;
   wire [34:0] stage2_62;
   wire [37:0] stage2_63;
   wire [45:0] stage2_64;
   wire [12:0] stage2_65;
   wire [9:0] stage2_66;
   wire [1:0] stage2_67;
   wire [7:0] stage3_0;
   wire [13:0] stage3_1;
   wire [10:0] stage3_2;
   wire [13:0] stage3_3;
   wire [13:0] stage3_4;
   wire [17:0] stage3_5;
   wire [19:0] stage3_6;
   wire [16:0] stage3_7;
   wire [16:0] stage3_8;
   wire [20:0] stage3_9;
   wire [14:0] stage3_10;
   wire [17:0] stage3_11;
   wire [23:0] stage3_12;
   wire [19:0] stage3_13;
   wire [35:0] stage3_14;
   wire [36:0] stage3_15;
   wire [21:0] stage3_16;
   wire [16:0] stage3_17;
   wire [22:0] stage3_18;
   wire [26:0] stage3_19;
   wire [22:0] stage3_20;
   wire [24:0] stage3_21;
   wire [26:0] stage3_22;
   wire [11:0] stage3_23;
   wire [25:0] stage3_24;
   wire [21:0] stage3_25;
   wire [15:0] stage3_26;
   wire [18:0] stage3_27;
   wire [19:0] stage3_28;
   wire [23:0] stage3_29;
   wire [25:0] stage3_30;
   wire [20:0] stage3_31;
   wire [34:0] stage3_32;
   wire [14:0] stage3_33;
   wire [22:0] stage3_34;
   wire [25:0] stage3_35;
   wire [16:0] stage3_36;
   wire [11:0] stage3_37;
   wire [13:0] stage3_38;
   wire [23:0] stage3_39;
   wire [23:0] stage3_40;
   wire [24:0] stage3_41;
   wire [25:0] stage3_42;
   wire [20:0] stage3_43;
   wire [30:0] stage3_44;
   wire [17:0] stage3_45;
   wire [16:0] stage3_46;
   wire [23:0] stage3_47;
   wire [15:0] stage3_48;
   wire [13:0] stage3_49;
   wire [31:0] stage3_50;
   wire [13:0] stage3_51;
   wire [23:0] stage3_52;
   wire [15:0] stage3_53;
   wire [15:0] stage3_54;
   wire [17:0] stage3_55;
   wire [30:0] stage3_56;
   wire [12:0] stage3_57;
   wire [32:0] stage3_58;
   wire [27:0] stage3_59;
   wire [14:0] stage3_60;
   wire [24:0] stage3_61;
   wire [20:0] stage3_62;
   wire [17:0] stage3_63;
   wire [28:0] stage3_64;
   wire [13:0] stage3_65;
   wire [8:0] stage3_66;
   wire [4:0] stage3_67;
   wire [1:0] stage3_68;
   wire [3:0] stage4_0;
   wire [3:0] stage4_1;
   wire [6:0] stage4_2;
   wire [4:0] stage4_3;
   wire [8:0] stage4_4;
   wire [8:0] stage4_5;
   wire [13:0] stage4_6;
   wire [7:0] stage4_7;
   wire [9:0] stage4_8;
   wire [6:0] stage4_9;
   wire [8:0] stage4_10;
   wire [6:0] stage4_11;
   wire [8:0] stage4_12;
   wire [9:0] stage4_13;
   wire [10:0] stage4_14;
   wire [16:0] stage4_15;
   wire [12:0] stage4_16;
   wire [16:0] stage4_17;
   wire [5:0] stage4_18;
   wire [15:0] stage4_19;
   wire [10:0] stage4_20;
   wire [7:0] stage4_21;
   wire [13:0] stage4_22;
   wire [9:0] stage4_23;
   wire [17:0] stage4_24;
   wire [5:0] stage4_25;
   wire [7:0] stage4_26;
   wire [6:0] stage4_27;
   wire [11:0] stage4_28;
   wire [9:0] stage4_29;
   wire [15:0] stage4_30;
   wire [8:0] stage4_31;
   wire [19:0] stage4_32;
   wire [11:0] stage4_33;
   wire [10:0] stage4_34;
   wire [10:0] stage4_35;
   wire [9:0] stage4_36;
   wire [5:0] stage4_37;
   wire [5:0] stage4_38;
   wire [9:0] stage4_39;
   wire [13:0] stage4_40;
   wire [16:0] stage4_41;
   wire [16:0] stage4_42;
   wire [6:0] stage4_43;
   wire [12:0] stage4_44;
   wire [8:0] stage4_45;
   wire [17:0] stage4_46;
   wire [15:0] stage4_47;
   wire [11:0] stage4_48;
   wire [12:0] stage4_49;
   wire [6:0] stage4_50;
   wire [8:0] stage4_51;
   wire [8:0] stage4_52;
   wire [14:0] stage4_53;
   wire [9:0] stage4_54;
   wire [16:0] stage4_55;
   wire [12:0] stage4_56;
   wire [5:0] stage4_57;
   wire [20:0] stage4_58;
   wire [16:0] stage4_59;
   wire [15:0] stage4_60;
   wire [16:0] stage4_61;
   wire [7:0] stage4_62;
   wire [12:0] stage4_63;
   wire [21:0] stage4_64;
   wire [5:0] stage4_65;
   wire [12:0] stage4_66;
   wire [6:0] stage4_67;
   wire [1:0] stage4_68;
   wire [1:0] stage5_0;
   wire [0:0] stage5_1;
   wire [4:0] stage5_2;
   wire [4:0] stage5_3;
   wire [4:0] stage5_4;
   wire [4:0] stage5_5;
   wire [9:0] stage5_6;
   wire [3:0] stage5_7;
   wire [7:0] stage5_8;
   wire [2:0] stage5_9;
   wire [4:0] stage5_10;
   wire [2:0] stage5_11;
   wire [10:0] stage5_12;
   wire [5:0] stage5_13;
   wire [7:0] stage5_14;
   wire [7:0] stage5_15;
   wire [8:0] stage5_16;
   wire [4:0] stage5_17;
   wire [5:0] stage5_18;
   wire [6:0] stage5_19;
   wire [3:0] stage5_20;
   wire [5:0] stage5_21;
   wire [10:0] stage5_22;
   wire [6:0] stage5_23;
   wire [9:0] stage5_24;
   wire [2:0] stage5_25;
   wire [2:0] stage5_26;
   wire [3:0] stage5_27;
   wire [4:0] stage5_28;
   wire [3:0] stage5_29;
   wire [4:0] stage5_30;
   wire [5:0] stage5_31;
   wire [11:0] stage5_32;
   wire [4:0] stage5_33;
   wire [7:0] stage5_34;
   wire [3:0] stage5_35;
   wire [4:0] stage5_36;
   wire [3:0] stage5_37;
   wire [1:0] stage5_38;
   wire [5:0] stage5_39;
   wire [5:0] stage5_40;
   wire [12:0] stage5_41;
   wire [4:0] stage5_42;
   wire [3:0] stage5_43;
   wire [5:0] stage5_44;
   wire [4:0] stage5_45;
   wire [5:0] stage5_46;
   wire [12:0] stage5_47;
   wire [3:0] stage5_48;
   wire [6:0] stage5_49;
   wire [4:0] stage5_50;
   wire [3:0] stage5_51;
   wire [5:0] stage5_52;
   wire [6:0] stage5_53;
   wire [8:0] stage5_54;
   wire [6:0] stage5_55;
   wire [4:0] stage5_56;
   wire [5:0] stage5_57;
   wire [5:0] stage5_58;
   wire [5:0] stage5_59;
   wire [8:0] stage5_60;
   wire [10:0] stage5_61;
   wire [5:0] stage5_62;
   wire [11:0] stage5_63;
   wire [10:0] stage5_64;
   wire [3:0] stage5_65;
   wire [4:0] stage5_66;
   wire [3:0] stage5_67;
   wire [4:0] stage5_68;
   wire [0:0] stage5_69;
   wire [1:0] stage6_0;
   wire [0:0] stage6_1;
   wire [4:0] stage6_2;
   wire [0:0] stage6_3;
   wire [4:0] stage6_4;
   wire [0:0] stage6_5;
   wire [2:0] stage6_6;
   wire [4:0] stage6_7;
   wire [1:0] stage6_8;
   wire [2:0] stage6_9;
   wire [6:0] stage6_10;
   wire [2:0] stage6_11;
   wire [5:0] stage6_12;
   wire [1:0] stage6_13;
   wire [3:0] stage6_14;
   wire [3:0] stage6_15;
   wire [5:0] stage6_16;
   wire [6:0] stage6_17;
   wire [0:0] stage6_18;
   wire [3:0] stage6_19;
   wire [2:0] stage6_20;
   wire [5:0] stage6_21;
   wire [3:0] stage6_22;
   wire [2:0] stage6_23;
   wire [2:0] stage6_24;
   wire [2:0] stage6_25;
   wire [2:0] stage6_26;
   wire [1:0] stage6_27;
   wire [2:0] stage6_28;
   wire [1:0] stage6_29;
   wire [1:0] stage6_30;
   wire [1:0] stage6_31;
   wire [8:0] stage6_32;
   wire [2:0] stage6_33;
   wire [2:0] stage6_34;
   wire [1:0] stage6_35;
   wire [6:0] stage6_36;
   wire [4:0] stage6_37;
   wire [0:0] stage6_38;
   wire [1:0] stage6_39;
   wire [1:0] stage6_40;
   wire [3:0] stage6_41;
   wire [7:0] stage6_42;
   wire [1:0] stage6_43;
   wire [1:0] stage6_44;
   wire [2:0] stage6_45;
   wire [1:0] stage6_46;
   wire [4:0] stage6_47;
   wire [5:0] stage6_48;
   wire [2:0] stage6_49;
   wire [3:0] stage6_50;
   wire [1:0] stage6_51;
   wire [3:0] stage6_52;
   wire [4:0] stage6_53;
   wire [2:0] stage6_54;
   wire [2:0] stage6_55;
   wire [4:0] stage6_56;
   wire [1:0] stage6_57;
   wire [1:0] stage6_58;
   wire [2:0] stage6_59;
   wire [4:0] stage6_60;
   wire [2:0] stage6_61;
   wire [3:0] stage6_62;
   wire [3:0] stage6_63;
   wire [3:0] stage6_64;
   wire [3:0] stage6_65;
   wire [2:0] stage6_66;
   wire [5:0] stage6_67;
   wire [5:0] stage6_68;
   wire [0:0] stage6_69;
   wire [1:0] stage7_0;
   wire [0:0] stage7_1;
   wire [0:0] stage7_2;
   wire [0:0] stage7_3;
   wire [1:0] stage7_4;
   wire [0:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [1:0] stage7_19;
   wire [1:0] stage7_20;
   wire [1:0] stage7_21;
   wire [1:0] stage7_22;
   wire [1:0] stage7_23;
   wire [1:0] stage7_24;
   wire [1:0] stage7_25;
   wire [0:0] stage7_26;
   wire [1:0] stage7_27;
   wire [1:0] stage7_28;
   wire [1:0] stage7_29;
   wire [1:0] stage7_30;
   wire [1:0] stage7_31;
   wire [1:0] stage7_32;
   wire [1:0] stage7_33;
   wire [1:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [1:0] stage7_37;
   wire [1:0] stage7_38;
   wire [1:0] stage7_39;
   wire [0:0] stage7_40;
   wire [1:0] stage7_41;
   wire [1:0] stage7_42;
   wire [1:0] stage7_43;
   wire [1:0] stage7_44;
   wire [1:0] stage7_45;
   wire [1:0] stage7_46;
   wire [1:0] stage7_47;
   wire [1:0] stage7_48;
   wire [1:0] stage7_49;
   wire [1:0] stage7_50;
   wire [1:0] stage7_51;
   wire [1:0] stage7_52;
   wire [1:0] stage7_53;
   wire [1:0] stage7_54;
   wire [1:0] stage7_55;
   wire [1:0] stage7_56;
   wire [1:0] stage7_57;
   wire [1:0] stage7_58;
   wire [1:0] stage7_59;
   wire [1:0] stage7_60;
   wire [0:0] stage7_61;
   wire [1:0] stage7_62;
   wire [1:0] stage7_63;
   wire [1:0] stage7_64;
   wire [1:0] stage7_65;
   wire [1:0] stage7_66;
   wire [1:0] stage7_67;
   wire [1:0] stage7_68;
   wire [1:0] stage7_69;
   wire [0:0] stage7_70;
   wire [0:0] stage7_71;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;
   assign dst21 = stage7_21;
   assign dst22 = stage7_22;
   assign dst23 = stage7_23;
   assign dst24 = stage7_24;
   assign dst25 = stage7_25;
   assign dst26 = stage7_26;
   assign dst27 = stage7_27;
   assign dst28 = stage7_28;
   assign dst29 = stage7_29;
   assign dst30 = stage7_30;
   assign dst31 = stage7_31;
   assign dst32 = stage7_32;
   assign dst33 = stage7_33;
   assign dst34 = stage7_34;
   assign dst35 = stage7_35;
   assign dst36 = stage7_36;
   assign dst37 = stage7_37;
   assign dst38 = stage7_38;
   assign dst39 = stage7_39;
   assign dst40 = stage7_40;
   assign dst41 = stage7_41;
   assign dst42 = stage7_42;
   assign dst43 = stage7_43;
   assign dst44 = stage7_44;
   assign dst45 = stage7_45;
   assign dst46 = stage7_46;
   assign dst47 = stage7_47;
   assign dst48 = stage7_48;
   assign dst49 = stage7_49;
   assign dst50 = stage7_50;
   assign dst51 = stage7_51;
   assign dst52 = stage7_52;
   assign dst53 = stage7_53;
   assign dst54 = stage7_54;
   assign dst55 = stage7_55;
   assign dst56 = stage7_56;
   assign dst57 = stage7_57;
   assign dst58 = stage7_58;
   assign dst59 = stage7_59;
   assign dst60 = stage7_60;
   assign dst61 = stage7_61;
   assign dst62 = stage7_62;
   assign dst63 = stage7_63;
   assign dst64 = stage7_64;
   assign dst65 = stage7_65;
   assign dst66 = stage7_66;
   assign dst67 = stage7_67;
   assign dst68 = stage7_68;
   assign dst69 = stage7_69;
   assign dst70 = stage7_70;
   assign dst71 = stage7_71;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7]},
      {stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[1]},
      {stage0_3[2]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[8], stage0_0[9], stage0_0[10]},
      {stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[2]},
      {stage0_3[3]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[3]},
      {stage0_3[4]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[4]},
      {stage0_3[5]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[5]},
      {stage0_3[6]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc1163_5 gpc6 (
      {stage0_0[20], stage0_0[21], stage0_0[22]},
      {stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_2[6]},
      {stage0_3[7]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc1163_5 gpc7 (
      {stage0_0[23], stage0_0[24], stage0_0[25]},
      {stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_2[7]},
      {stage0_3[8]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1163_5 gpc8 (
      {stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_2[8]},
      {stage0_3[9]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc1163_5 gpc9 (
      {stage0_0[29], stage0_0[30], stage0_0[31]},
      {stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56]},
      {stage0_2[9]},
      {stage0_3[10]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62]},
      {stage0_2[10]},
      {stage0_3[11]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68]},
      {stage0_2[11]},
      {stage0_3[12]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[38], stage0_0[39], stage0_0[40]},
      {stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74]},
      {stage0_2[12]},
      {stage0_3[13]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[41], stage0_0[42], stage0_0[43]},
      {stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80]},
      {stage0_2[13]},
      {stage0_3[14]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc207_4 gpc14 (
      {stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[14], stage0_2[15]},
      {stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21]},
      {stage1_4[14],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27]},
      {stage1_4[15],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33]},
      {stage1_4[16],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39]},
      {stage1_4[17],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45]},
      {stage1_4[18],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51]},
      {stage1_4[19],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57]},
      {stage1_4[20],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63]},
      {stage1_4[21],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69]},
      {stage1_4[22],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75]},
      {stage1_4[23],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81]},
      {stage1_4[24],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121], stage0_0[122]},
      {stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87]},
      {stage1_4[25],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127], stage0_0[128]},
      {stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93]},
      {stage1_4[26],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134]},
      {stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99]},
      {stage1_4[27],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140]},
      {stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105]},
      {stage1_4[28],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146]},
      {stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111]},
      {stage1_4[29],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc615_5 gpc31 (
      {stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151]},
      {stage0_1[81]},
      {stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117]},
      {stage1_4[30],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc615_5 gpc32 (
      {stage0_0[152], stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_1[82]},
      {stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123]},
      {stage1_4[31],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc615_5 gpc33 (
      {stage0_0[157], stage0_0[158], stage0_0[159], stage0_0[160], stage0_0[161]},
      {stage0_1[83]},
      {stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129]},
      {stage1_4[32],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[0],stage1_4[33],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[1],stage1_4[34],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[2],stage1_4[35],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[3],stage1_4[36],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[4],stage1_4[37],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[5],stage1_4[38],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[6],stage1_4[39],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[7],stage1_4[40],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[8],stage1_4[41],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[9],stage1_4[42],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[10],stage1_4[43],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[11],stage1_4[44],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[12],stage1_4[45],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc615_5 gpc47 (
      {stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage0_3[93]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[13],stage1_4[46],stage1_3[47],stage1_2[47]}
   );
   gpc615_5 gpc48 (
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139]},
      {stage0_3[94]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[14],stage1_4[47],stage1_3[48],stage1_2[48]}
   );
   gpc615_5 gpc49 (
      {stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage0_3[95]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[15],stage1_4[48],stage1_3[49],stage1_2[49]}
   );
   gpc615_5 gpc50 (
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149]},
      {stage0_3[96]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[16],stage1_4[49],stage1_3[50],stage1_2[50]}
   );
   gpc615_5 gpc51 (
      {stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154]},
      {stage0_3[97]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[17],stage1_4[50],stage1_3[51],stage1_2[51]}
   );
   gpc615_5 gpc52 (
      {stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158], stage0_2[159]},
      {stage0_3[98]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[18],stage1_4[51],stage1_3[52],stage1_2[52]}
   );
   gpc615_5 gpc53 (
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103]},
      {stage0_4[36]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[6],stage1_5[19],stage1_4[52],stage1_3[53]}
   );
   gpc615_5 gpc54 (
      {stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108]},
      {stage0_4[37]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[7],stage1_5[20],stage1_4[53],stage1_3[54]}
   );
   gpc615_5 gpc55 (
      {stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113]},
      {stage0_4[38]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[8],stage1_5[21],stage1_4[54],stage1_3[55]}
   );
   gpc615_5 gpc56 (
      {stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118]},
      {stage0_4[39]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[9],stage1_5[22],stage1_4[55],stage1_3[56]}
   );
   gpc615_5 gpc57 (
      {stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage0_4[40]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[10],stage1_5[23],stage1_4[56],stage1_3[57]}
   );
   gpc615_5 gpc58 (
      {stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128]},
      {stage0_4[41]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[11],stage1_5[24],stage1_4[57],stage1_3[58]}
   );
   gpc615_5 gpc59 (
      {stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133]},
      {stage0_4[42]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[12],stage1_5[25],stage1_4[58],stage1_3[59]}
   );
   gpc615_5 gpc60 (
      {stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138]},
      {stage0_4[43]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[13],stage1_5[26],stage1_4[59],stage1_3[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[8],stage1_6[14],stage1_5[27],stage1_4[60]}
   );
   gpc606_5 gpc62 (
      {stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[9],stage1_6[15],stage1_5[28],stage1_4[61]}
   );
   gpc606_5 gpc63 (
      {stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[10],stage1_6[16],stage1_5[29],stage1_4[62]}
   );
   gpc606_5 gpc64 (
      {stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[11],stage1_6[17],stage1_5[30],stage1_4[63]}
   );
   gpc606_5 gpc65 (
      {stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[12],stage1_6[18],stage1_5[31],stage1_4[64]}
   );
   gpc606_5 gpc66 (
      {stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[13],stage1_6[19],stage1_5[32],stage1_4[65]}
   );
   gpc606_5 gpc67 (
      {stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[14],stage1_6[20],stage1_5[33],stage1_4[66]}
   );
   gpc606_5 gpc68 (
      {stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[15],stage1_6[21],stage1_5[34],stage1_4[67]}
   );
   gpc606_5 gpc69 (
      {stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[16],stage1_6[22],stage1_5[35],stage1_4[68]}
   );
   gpc606_5 gpc70 (
      {stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[17],stage1_6[23],stage1_5[36],stage1_4[69]}
   );
   gpc606_5 gpc71 (
      {stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[18],stage1_6[24],stage1_5[37],stage1_4[70]}
   );
   gpc606_5 gpc72 (
      {stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[19],stage1_6[25],stage1_5[38],stage1_4[71]}
   );
   gpc606_5 gpc73 (
      {stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[20],stage1_6[26],stage1_5[39],stage1_4[72]}
   );
   gpc606_5 gpc74 (
      {stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[21],stage1_6[27],stage1_5[40],stage1_4[73]}
   );
   gpc606_5 gpc75 (
      {stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[22],stage1_6[28],stage1_5[41],stage1_4[74]}
   );
   gpc606_5 gpc76 (
      {stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[23],stage1_6[29],stage1_5[42],stage1_4[75]}
   );
   gpc606_5 gpc77 (
      {stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[24],stage1_6[30],stage1_5[43],stage1_4[76]}
   );
   gpc606_5 gpc78 (
      {stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[25],stage1_6[31],stage1_5[44],stage1_4[77]}
   );
   gpc606_5 gpc79 (
      {stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[26],stage1_6[32],stage1_5[45],stage1_4[78]}
   );
   gpc606_5 gpc80 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[19],stage1_7[27],stage1_6[33],stage1_5[46]}
   );
   gpc606_5 gpc81 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[20],stage1_7[28],stage1_6[34],stage1_5[47]}
   );
   gpc606_5 gpc82 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[21],stage1_7[29],stage1_6[35],stage1_5[48]}
   );
   gpc606_5 gpc83 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[22],stage1_7[30],stage1_6[36],stage1_5[49]}
   );
   gpc606_5 gpc84 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[23],stage1_7[31],stage1_6[37],stage1_5[50]}
   );
   gpc606_5 gpc85 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[24],stage1_7[32],stage1_6[38],stage1_5[51]}
   );
   gpc606_5 gpc86 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[25],stage1_7[33],stage1_6[39],stage1_5[52]}
   );
   gpc606_5 gpc87 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[26],stage1_7[34],stage1_6[40],stage1_5[53]}
   );
   gpc606_5 gpc88 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[27],stage1_7[35],stage1_6[41],stage1_5[54]}
   );
   gpc615_5 gpc89 (
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118]},
      {stage0_7[54]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[9],stage1_8[28],stage1_7[36],stage1_6[42]}
   );
   gpc615_5 gpc90 (
      {stage0_6[119], stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123]},
      {stage0_7[55]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[10],stage1_8[29],stage1_7[37],stage1_6[43]}
   );
   gpc615_5 gpc91 (
      {stage0_6[124], stage0_6[125], stage0_6[126], stage0_6[127], stage0_6[128]},
      {stage0_7[56]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[11],stage1_8[30],stage1_7[38],stage1_6[44]}
   );
   gpc615_5 gpc92 (
      {stage0_6[129], stage0_6[130], stage0_6[131], stage0_6[132], stage0_6[133]},
      {stage0_7[57]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[12],stage1_8[31],stage1_7[39],stage1_6[45]}
   );
   gpc615_5 gpc93 (
      {stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137], stage0_6[138]},
      {stage0_7[58]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[13],stage1_8[32],stage1_7[40],stage1_6[46]}
   );
   gpc615_5 gpc94 (
      {stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage0_7[59]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[14],stage1_8[33],stage1_7[41],stage1_6[47]}
   );
   gpc615_5 gpc95 (
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148]},
      {stage0_7[60]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[15],stage1_8[34],stage1_7[42],stage1_6[48]}
   );
   gpc615_5 gpc96 (
      {stage0_6[149], stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153]},
      {stage0_7[61]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[16],stage1_8[35],stage1_7[43],stage1_6[49]}
   );
   gpc606_5 gpc97 (
      {stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65], stage0_7[66], stage0_7[67]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[8],stage1_9[17],stage1_8[36],stage1_7[44]}
   );
   gpc615_5 gpc98 (
      {stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71], stage0_7[72]},
      {stage0_8[48]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[9],stage1_9[18],stage1_8[37],stage1_7[45]}
   );
   gpc615_5 gpc99 (
      {stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage0_8[49]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[10],stage1_9[19],stage1_8[38],stage1_7[46]}
   );
   gpc615_5 gpc100 (
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82]},
      {stage0_8[50]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[11],stage1_9[20],stage1_8[39],stage1_7[47]}
   );
   gpc615_5 gpc101 (
      {stage0_7[83], stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87]},
      {stage0_8[51]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[12],stage1_9[21],stage1_8[40],stage1_7[48]}
   );
   gpc615_5 gpc102 (
      {stage0_7[88], stage0_7[89], stage0_7[90], stage0_7[91], stage0_7[92]},
      {stage0_8[52]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[13],stage1_9[22],stage1_8[41],stage1_7[49]}
   );
   gpc615_5 gpc103 (
      {stage0_7[93], stage0_7[94], stage0_7[95], stage0_7[96], stage0_7[97]},
      {stage0_8[53]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[14],stage1_9[23],stage1_8[42],stage1_7[50]}
   );
   gpc615_5 gpc104 (
      {stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101], stage0_7[102]},
      {stage0_8[54]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[15],stage1_9[24],stage1_8[43],stage1_7[51]}
   );
   gpc615_5 gpc105 (
      {stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage0_8[55]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[16],stage1_9[25],stage1_8[44],stage1_7[52]}
   );
   gpc615_5 gpc106 (
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112]},
      {stage0_8[56]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[17],stage1_9[26],stage1_8[45],stage1_7[53]}
   );
   gpc615_5 gpc107 (
      {stage0_7[113], stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117]},
      {stage0_8[57]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[18],stage1_9[27],stage1_8[46],stage1_7[54]}
   );
   gpc615_5 gpc108 (
      {stage0_7[118], stage0_7[119], stage0_7[120], stage0_7[121], stage0_7[122]},
      {stage0_8[58]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[19],stage1_9[28],stage1_8[47],stage1_7[55]}
   );
   gpc615_5 gpc109 (
      {stage0_7[123], stage0_7[124], stage0_7[125], stage0_7[126], stage0_7[127]},
      {stage0_8[59]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[20],stage1_9[29],stage1_8[48],stage1_7[56]}
   );
   gpc615_5 gpc110 (
      {stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131], stage0_7[132]},
      {stage0_8[60]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[21],stage1_9[30],stage1_8[49],stage1_7[57]}
   );
   gpc615_5 gpc111 (
      {stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage0_8[61]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[22],stage1_9[31],stage1_8[50],stage1_7[58]}
   );
   gpc615_5 gpc112 (
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142]},
      {stage0_8[62]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[23],stage1_9[32],stage1_8[51],stage1_7[59]}
   );
   gpc615_5 gpc113 (
      {stage0_7[143], stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147]},
      {stage0_8[63]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[24],stage1_9[33],stage1_8[52],stage1_7[60]}
   );
   gpc615_5 gpc114 (
      {stage0_7[148], stage0_7[149], stage0_7[150], stage0_7[151], stage0_7[152]},
      {stage0_8[64]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[25],stage1_9[34],stage1_8[53],stage1_7[61]}
   );
   gpc606_5 gpc115 (
      {stage0_8[65], stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[18],stage1_10[26],stage1_9[35],stage1_8[54]}
   );
   gpc606_5 gpc116 (
      {stage0_8[71], stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[19],stage1_10[27],stage1_9[36],stage1_8[55]}
   );
   gpc606_5 gpc117 (
      {stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[20],stage1_10[28],stage1_9[37],stage1_8[56]}
   );
   gpc606_5 gpc118 (
      {stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[21],stage1_10[29],stage1_9[38],stage1_8[57]}
   );
   gpc606_5 gpc119 (
      {stage0_8[89], stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[22],stage1_10[30],stage1_9[39],stage1_8[58]}
   );
   gpc606_5 gpc120 (
      {stage0_8[95], stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[23],stage1_10[31],stage1_9[40],stage1_8[59]}
   );
   gpc606_5 gpc121 (
      {stage0_8[101], stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[24],stage1_10[32],stage1_9[41],stage1_8[60]}
   );
   gpc606_5 gpc122 (
      {stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[25],stage1_10[33],stage1_9[42],stage1_8[61]}
   );
   gpc606_5 gpc123 (
      {stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[26],stage1_10[34],stage1_9[43],stage1_8[62]}
   );
   gpc606_5 gpc124 (
      {stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[27],stage1_10[35],stage1_9[44],stage1_8[63]}
   );
   gpc606_5 gpc125 (
      {stage0_8[125], stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[28],stage1_10[36],stage1_9[45],stage1_8[64]}
   );
   gpc606_5 gpc126 (
      {stage0_8[131], stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[29],stage1_10[37],stage1_9[46],stage1_8[65]}
   );
   gpc606_5 gpc127 (
      {stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[30],stage1_10[38],stage1_9[47],stage1_8[66]}
   );
   gpc606_5 gpc128 (
      {stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[31],stage1_10[39],stage1_9[48],stage1_8[67]}
   );
   gpc606_5 gpc129 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[14],stage1_11[32],stage1_10[40],stage1_9[49]}
   );
   gpc606_5 gpc130 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[15],stage1_11[33],stage1_10[41],stage1_9[50]}
   );
   gpc606_5 gpc131 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[16],stage1_11[34],stage1_10[42],stage1_9[51]}
   );
   gpc606_5 gpc132 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[17],stage1_11[35],stage1_10[43],stage1_9[52]}
   );
   gpc606_5 gpc133 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[18],stage1_11[36],stage1_10[44],stage1_9[53]}
   );
   gpc606_5 gpc134 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[19],stage1_11[37],stage1_10[45],stage1_9[54]}
   );
   gpc606_5 gpc135 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[20],stage1_11[38],stage1_10[46],stage1_9[55]}
   );
   gpc606_5 gpc136 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[21],stage1_11[39],stage1_10[47],stage1_9[56]}
   );
   gpc606_5 gpc137 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160], stage0_9[161]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[22],stage1_11[40],stage1_10[48],stage1_9[57]}
   );
   gpc615_5 gpc138 (
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88]},
      {stage0_11[54]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[9],stage1_12[23],stage1_11[41],stage1_10[49]}
   );
   gpc615_5 gpc139 (
      {stage0_10[89], stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93]},
      {stage0_11[55]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[10],stage1_12[24],stage1_11[42],stage1_10[50]}
   );
   gpc615_5 gpc140 (
      {stage0_10[94], stage0_10[95], stage0_10[96], stage0_10[97], stage0_10[98]},
      {stage0_11[56]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[11],stage1_12[25],stage1_11[43],stage1_10[51]}
   );
   gpc615_5 gpc141 (
      {stage0_10[99], stage0_10[100], stage0_10[101], stage0_10[102], stage0_10[103]},
      {stage0_11[57]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[12],stage1_12[26],stage1_11[44],stage1_10[52]}
   );
   gpc615_5 gpc142 (
      {stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107], stage0_10[108]},
      {stage0_11[58]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[13],stage1_12[27],stage1_11[45],stage1_10[53]}
   );
   gpc615_5 gpc143 (
      {stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage0_11[59]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[14],stage1_12[28],stage1_11[46],stage1_10[54]}
   );
   gpc615_5 gpc144 (
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118]},
      {stage0_11[60]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[15],stage1_12[29],stage1_11[47],stage1_10[55]}
   );
   gpc615_5 gpc145 (
      {stage0_10[119], stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123]},
      {stage0_11[61]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[16],stage1_12[30],stage1_11[48],stage1_10[56]}
   );
   gpc606_5 gpc146 (
      {stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65], stage0_11[66], stage0_11[67]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[8],stage1_13[17],stage1_12[31],stage1_11[49]}
   );
   gpc606_5 gpc147 (
      {stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71], stage0_11[72], stage0_11[73]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[9],stage1_13[18],stage1_12[32],stage1_11[50]}
   );
   gpc606_5 gpc148 (
      {stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77], stage0_11[78], stage0_11[79]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[10],stage1_13[19],stage1_12[33],stage1_11[51]}
   );
   gpc606_5 gpc149 (
      {stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83], stage0_11[84], stage0_11[85]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[11],stage1_13[20],stage1_12[34],stage1_11[52]}
   );
   gpc606_5 gpc150 (
      {stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89], stage0_11[90], stage0_11[91]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[12],stage1_13[21],stage1_12[35],stage1_11[53]}
   );
   gpc606_5 gpc151 (
      {stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95], stage0_11[96], stage0_11[97]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[13],stage1_13[22],stage1_12[36],stage1_11[54]}
   );
   gpc606_5 gpc152 (
      {stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101], stage0_11[102], stage0_11[103]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[14],stage1_13[23],stage1_12[37],stage1_11[55]}
   );
   gpc606_5 gpc153 (
      {stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107], stage0_11[108], stage0_11[109]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[15],stage1_13[24],stage1_12[38],stage1_11[56]}
   );
   gpc606_5 gpc154 (
      {stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113], stage0_11[114], stage0_11[115]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[16],stage1_13[25],stage1_12[39],stage1_11[57]}
   );
   gpc606_5 gpc155 (
      {stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119], stage0_11[120], stage0_11[121]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[17],stage1_13[26],stage1_12[40],stage1_11[58]}
   );
   gpc606_5 gpc156 (
      {stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125], stage0_11[126], stage0_11[127]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[18],stage1_13[27],stage1_12[41],stage1_11[59]}
   );
   gpc606_5 gpc157 (
      {stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131], stage0_11[132], stage0_11[133]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[19],stage1_13[28],stage1_12[42],stage1_11[60]}
   );
   gpc615_5 gpc158 (
      {stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137], stage0_11[138]},
      {stage0_12[48]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[20],stage1_13[29],stage1_12[43],stage1_11[61]}
   );
   gpc615_5 gpc159 (
      {stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage0_12[49]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[21],stage1_13[30],stage1_12[44],stage1_11[62]}
   );
   gpc606_5 gpc160 (
      {stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[14],stage1_14[22],stage1_13[31],stage1_12[45]}
   );
   gpc606_5 gpc161 (
      {stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[15],stage1_14[23],stage1_13[32],stage1_12[46]}
   );
   gpc606_5 gpc162 (
      {stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65], stage0_12[66], stage0_12[67]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[16],stage1_14[24],stage1_13[33],stage1_12[47]}
   );
   gpc606_5 gpc163 (
      {stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71], stage0_12[72], stage0_12[73]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[17],stage1_14[25],stage1_13[34],stage1_12[48]}
   );
   gpc606_5 gpc164 (
      {stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77], stage0_12[78], stage0_12[79]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[18],stage1_14[26],stage1_13[35],stage1_12[49]}
   );
   gpc606_5 gpc165 (
      {stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83], stage0_12[84], stage0_12[85]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[19],stage1_14[27],stage1_13[36],stage1_12[50]}
   );
   gpc606_5 gpc166 (
      {stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89], stage0_12[90], stage0_12[91]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[20],stage1_14[28],stage1_13[37],stage1_12[51]}
   );
   gpc606_5 gpc167 (
      {stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95], stage0_12[96], stage0_12[97]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[21],stage1_14[29],stage1_13[38],stage1_12[52]}
   );
   gpc606_5 gpc168 (
      {stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[22],stage1_14[30],stage1_13[39],stage1_12[53]}
   );
   gpc606_5 gpc169 (
      {stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[23],stage1_14[31],stage1_13[40],stage1_12[54]}
   );
   gpc606_5 gpc170 (
      {stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[24],stage1_14[32],stage1_13[41],stage1_12[55]}
   );
   gpc606_5 gpc171 (
      {stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[25],stage1_14[33],stage1_13[42],stage1_12[56]}
   );
   gpc606_5 gpc172 (
      {stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[26],stage1_14[34],stage1_13[43],stage1_12[57]}
   );
   gpc606_5 gpc173 (
      {stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[27],stage1_14[35],stage1_13[44],stage1_12[58]}
   );
   gpc606_5 gpc174 (
      {stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[28],stage1_14[36],stage1_13[45],stage1_12[59]}
   );
   gpc606_5 gpc175 (
      {stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[29],stage1_14[37],stage1_13[46],stage1_12[60]}
   );
   gpc606_5 gpc176 (
      {stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[30],stage1_14[38],stage1_13[47],stage1_12[61]}
   );
   gpc606_5 gpc177 (
      {stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155], stage0_12[156], stage0_12[157]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[31],stage1_14[39],stage1_13[48],stage1_12[62]}
   );
   gpc606_5 gpc178 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[18],stage1_15[32],stage1_14[40],stage1_13[49]}
   );
   gpc606_5 gpc179 (
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[19],stage1_15[33],stage1_14[41],stage1_13[50]}
   );
   gpc606_5 gpc180 (
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[20],stage1_15[34],stage1_14[42],stage1_13[51]}
   );
   gpc606_5 gpc181 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[21],stage1_15[35],stage1_14[43],stage1_13[52]}
   );
   gpc606_5 gpc182 (
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[22],stage1_15[36],stage1_14[44],stage1_13[53]}
   );
   gpc606_5 gpc183 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[23],stage1_15[37],stage1_14[45],stage1_13[54]}
   );
   gpc606_5 gpc184 (
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[24],stage1_15[38],stage1_14[46],stage1_13[55]}
   );
   gpc606_5 gpc185 (
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[25],stage1_15[39],stage1_14[47],stage1_13[56]}
   );
   gpc615_5 gpc186 (
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112]},
      {stage0_15[48]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[8],stage1_16[26],stage1_15[40],stage1_14[48]}
   );
   gpc615_5 gpc187 (
      {stage0_14[113], stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117]},
      {stage0_15[49]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[9],stage1_16[27],stage1_15[41],stage1_14[49]}
   );
   gpc615_5 gpc188 (
      {stage0_14[118], stage0_14[119], stage0_14[120], stage0_14[121], stage0_14[122]},
      {stage0_15[50]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[10],stage1_16[28],stage1_15[42],stage1_14[50]}
   );
   gpc615_5 gpc189 (
      {stage0_14[123], stage0_14[124], stage0_14[125], stage0_14[126], stage0_14[127]},
      {stage0_15[51]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[11],stage1_16[29],stage1_15[43],stage1_14[51]}
   );
   gpc615_5 gpc190 (
      {stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132]},
      {stage0_15[52]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[12],stage1_16[30],stage1_15[44],stage1_14[52]}
   );
   gpc615_5 gpc191 (
      {stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage0_15[53]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[13],stage1_16[31],stage1_15[45],stage1_14[53]}
   );
   gpc615_5 gpc192 (
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142]},
      {stage0_15[54]},
      {stage0_16[36], stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41]},
      {stage1_18[6],stage1_17[14],stage1_16[32],stage1_15[46],stage1_14[54]}
   );
   gpc615_5 gpc193 (
      {stage0_14[143], stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147]},
      {stage0_15[55]},
      {stage0_16[42], stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47]},
      {stage1_18[7],stage1_17[15],stage1_16[33],stage1_15[47],stage1_14[55]}
   );
   gpc615_5 gpc194 (
      {stage0_14[148], stage0_14[149], stage0_14[150], stage0_14[151], stage0_14[152]},
      {stage0_15[56]},
      {stage0_16[48], stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53]},
      {stage1_18[8],stage1_17[16],stage1_16[34],stage1_15[48],stage1_14[56]}
   );
   gpc615_5 gpc195 (
      {stage0_14[153], stage0_14[154], stage0_14[155], stage0_14[156], stage0_14[157]},
      {stage0_15[57]},
      {stage0_16[54], stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59]},
      {stage1_18[9],stage1_17[17],stage1_16[35],stage1_15[49],stage1_14[57]}
   );
   gpc615_5 gpc196 (
      {stage0_15[58], stage0_15[59], stage0_15[60], stage0_15[61], stage0_15[62]},
      {stage0_16[60]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[10],stage1_17[18],stage1_16[36],stage1_15[50]}
   );
   gpc615_5 gpc197 (
      {stage0_15[63], stage0_15[64], stage0_15[65], stage0_15[66], stage0_15[67]},
      {stage0_16[61]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[11],stage1_17[19],stage1_16[37],stage1_15[51]}
   );
   gpc615_5 gpc198 (
      {stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71], stage0_15[72]},
      {stage0_16[62]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[12],stage1_17[20],stage1_16[38],stage1_15[52]}
   );
   gpc615_5 gpc199 (
      {stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage0_16[63]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[13],stage1_17[21],stage1_16[39],stage1_15[53]}
   );
   gpc615_5 gpc200 (
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82]},
      {stage0_16[64]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[14],stage1_17[22],stage1_16[40],stage1_15[54]}
   );
   gpc615_5 gpc201 (
      {stage0_15[83], stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87]},
      {stage0_16[65]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[15],stage1_17[23],stage1_16[41],stage1_15[55]}
   );
   gpc615_5 gpc202 (
      {stage0_15[88], stage0_15[89], stage0_15[90], stage0_15[91], stage0_15[92]},
      {stage0_16[66]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[16],stage1_17[24],stage1_16[42],stage1_15[56]}
   );
   gpc615_5 gpc203 (
      {stage0_15[93], stage0_15[94], stage0_15[95], stage0_15[96], stage0_15[97]},
      {stage0_16[67]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[17],stage1_17[25],stage1_16[43],stage1_15[57]}
   );
   gpc615_5 gpc204 (
      {stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101], stage0_15[102]},
      {stage0_16[68]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[18],stage1_17[26],stage1_16[44],stage1_15[58]}
   );
   gpc615_5 gpc205 (
      {stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage0_16[69]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[19],stage1_17[27],stage1_16[45],stage1_15[59]}
   );
   gpc615_5 gpc206 (
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112]},
      {stage0_16[70]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[20],stage1_17[28],stage1_16[46],stage1_15[60]}
   );
   gpc615_5 gpc207 (
      {stage0_15[113], stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117]},
      {stage0_16[71]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[21],stage1_17[29],stage1_16[47],stage1_15[61]}
   );
   gpc615_5 gpc208 (
      {stage0_15[118], stage0_15[119], stage0_15[120], stage0_15[121], stage0_15[122]},
      {stage0_16[72]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[22],stage1_17[30],stage1_16[48],stage1_15[62]}
   );
   gpc615_5 gpc209 (
      {stage0_15[123], stage0_15[124], stage0_15[125], stage0_15[126], stage0_15[127]},
      {stage0_16[73]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[23],stage1_17[31],stage1_16[49],stage1_15[63]}
   );
   gpc606_5 gpc210 (
      {stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77], stage0_16[78], stage0_16[79]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[14],stage1_18[24],stage1_17[32],stage1_16[50]}
   );
   gpc606_5 gpc211 (
      {stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83], stage0_16[84], stage0_16[85]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[15],stage1_18[25],stage1_17[33],stage1_16[51]}
   );
   gpc606_5 gpc212 (
      {stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90], stage0_16[91]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[16],stage1_18[26],stage1_17[34],stage1_16[52]}
   );
   gpc606_5 gpc213 (
      {stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96], stage0_16[97]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[17],stage1_18[27],stage1_17[35],stage1_16[53]}
   );
   gpc606_5 gpc214 (
      {stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102], stage0_16[103]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[18],stage1_18[28],stage1_17[36],stage1_16[54]}
   );
   gpc606_5 gpc215 (
      {stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108], stage0_16[109]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[19],stage1_18[29],stage1_17[37],stage1_16[55]}
   );
   gpc606_5 gpc216 (
      {stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113], stage0_16[114], stage0_16[115]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[20],stage1_18[30],stage1_17[38],stage1_16[56]}
   );
   gpc606_5 gpc217 (
      {stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119], stage0_16[120], stage0_16[121]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[21],stage1_18[31],stage1_17[39],stage1_16[57]}
   );
   gpc606_5 gpc218 (
      {stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126], stage0_16[127]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[22],stage1_18[32],stage1_17[40],stage1_16[58]}
   );
   gpc606_5 gpc219 (
      {stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132], stage0_16[133]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[23],stage1_18[33],stage1_17[41],stage1_16[59]}
   );
   gpc606_5 gpc220 (
      {stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138], stage0_16[139]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[24],stage1_18[34],stage1_17[42],stage1_16[60]}
   );
   gpc606_5 gpc221 (
      {stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144], stage0_16[145]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[25],stage1_18[35],stage1_17[43],stage1_16[61]}
   );
   gpc606_5 gpc222 (
      {stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[26],stage1_18[36],stage1_17[44],stage1_16[62]}
   );
   gpc606_5 gpc223 (
      {stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[27],stage1_18[37],stage1_17[45],stage1_16[63]}
   );
   gpc606_5 gpc224 (
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[14],stage1_19[28],stage1_18[38],stage1_17[46]}
   );
   gpc606_5 gpc225 (
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[15],stage1_19[29],stage1_18[39],stage1_17[47]}
   );
   gpc606_5 gpc226 (
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[2],stage1_20[16],stage1_19[30],stage1_18[40]}
   );
   gpc606_5 gpc227 (
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[3],stage1_20[17],stage1_19[31],stage1_18[41]}
   );
   gpc606_5 gpc228 (
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[4],stage1_20[18],stage1_19[32],stage1_18[42]}
   );
   gpc606_5 gpc229 (
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[5],stage1_20[19],stage1_19[33],stage1_18[43]}
   );
   gpc606_5 gpc230 (
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[6],stage1_20[20],stage1_19[34],stage1_18[44]}
   );
   gpc606_5 gpc231 (
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[7],stage1_20[21],stage1_19[35],stage1_18[45]}
   );
   gpc606_5 gpc232 (
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[8],stage1_20[22],stage1_19[36],stage1_18[46]}
   );
   gpc615_5 gpc233 (
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130]},
      {stage0_19[12]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[9],stage1_20[23],stage1_19[37],stage1_18[47]}
   );
   gpc615_5 gpc234 (
      {stage0_18[131], stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135]},
      {stage0_19[13]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[10],stage1_20[24],stage1_19[38],stage1_18[48]}
   );
   gpc615_5 gpc235 (
      {stage0_18[136], stage0_18[137], stage0_18[138], stage0_18[139], stage0_18[140]},
      {stage0_19[14]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[11],stage1_20[25],stage1_19[39],stage1_18[49]}
   );
   gpc615_5 gpc236 (
      {stage0_18[141], stage0_18[142], stage0_18[143], stage0_18[144], stage0_18[145]},
      {stage0_19[15]},
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65]},
      {stage1_22[10],stage1_21[12],stage1_20[26],stage1_19[40],stage1_18[50]}
   );
   gpc615_5 gpc237 (
      {stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149], stage0_18[150]},
      {stage0_19[16]},
      {stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69], stage0_20[70], stage0_20[71]},
      {stage1_22[11],stage1_21[13],stage1_20[27],stage1_19[41],stage1_18[51]}
   );
   gpc207_4 gpc238 (
      {stage0_19[17], stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage0_21[0], stage0_21[1]},
      {stage1_22[12],stage1_21[14],stage1_20[28],stage1_19[42]}
   );
   gpc207_4 gpc239 (
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29], stage0_19[30]},
      {stage0_21[2], stage0_21[3]},
      {stage1_22[13],stage1_21[15],stage1_20[29],stage1_19[43]}
   );
   gpc207_4 gpc240 (
      {stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35], stage0_19[36], stage0_19[37]},
      {stage0_21[4], stage0_21[5]},
      {stage1_22[14],stage1_21[16],stage1_20[30],stage1_19[44]}
   );
   gpc207_4 gpc241 (
      {stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41], stage0_19[42], stage0_19[43], stage0_19[44]},
      {stage0_21[6], stage0_21[7]},
      {stage1_22[15],stage1_21[17],stage1_20[31],stage1_19[45]}
   );
   gpc606_5 gpc242 (
      {stage0_19[45], stage0_19[46], stage0_19[47], stage0_19[48], stage0_19[49], stage0_19[50]},
      {stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11], stage0_21[12], stage0_21[13]},
      {stage1_23[0],stage1_22[16],stage1_21[18],stage1_20[32],stage1_19[46]}
   );
   gpc606_5 gpc243 (
      {stage0_19[51], stage0_19[52], stage0_19[53], stage0_19[54], stage0_19[55], stage0_19[56]},
      {stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17], stage0_21[18], stage0_21[19]},
      {stage1_23[1],stage1_22[17],stage1_21[19],stage1_20[33],stage1_19[47]}
   );
   gpc606_5 gpc244 (
      {stage0_19[57], stage0_19[58], stage0_19[59], stage0_19[60], stage0_19[61], stage0_19[62]},
      {stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25]},
      {stage1_23[2],stage1_22[18],stage1_21[20],stage1_20[34],stage1_19[48]}
   );
   gpc606_5 gpc245 (
      {stage0_19[63], stage0_19[64], stage0_19[65], stage0_19[66], stage0_19[67], stage0_19[68]},
      {stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30], stage0_21[31]},
      {stage1_23[3],stage1_22[19],stage1_21[21],stage1_20[35],stage1_19[49]}
   );
   gpc606_5 gpc246 (
      {stage0_19[69], stage0_19[70], stage0_19[71], stage0_19[72], stage0_19[73], stage0_19[74]},
      {stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35], stage0_21[36], stage0_21[37]},
      {stage1_23[4],stage1_22[20],stage1_21[22],stage1_20[36],stage1_19[50]}
   );
   gpc606_5 gpc247 (
      {stage0_19[75], stage0_19[76], stage0_19[77], stage0_19[78], stage0_19[79], stage0_19[80]},
      {stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42], stage0_21[43]},
      {stage1_23[5],stage1_22[21],stage1_21[23],stage1_20[37],stage1_19[51]}
   );
   gpc606_5 gpc248 (
      {stage0_19[81], stage0_19[82], stage0_19[83], stage0_19[84], stage0_19[85], stage0_19[86]},
      {stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47], stage0_21[48], stage0_21[49]},
      {stage1_23[6],stage1_22[22],stage1_21[24],stage1_20[38],stage1_19[52]}
   );
   gpc606_5 gpc249 (
      {stage0_19[87], stage0_19[88], stage0_19[89], stage0_19[90], stage0_19[91], stage0_19[92]},
      {stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53], stage0_21[54], stage0_21[55]},
      {stage1_23[7],stage1_22[23],stage1_21[25],stage1_20[39],stage1_19[53]}
   );
   gpc606_5 gpc250 (
      {stage0_19[93], stage0_19[94], stage0_19[95], stage0_19[96], stage0_19[97], stage0_19[98]},
      {stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59], stage0_21[60], stage0_21[61]},
      {stage1_23[8],stage1_22[24],stage1_21[26],stage1_20[40],stage1_19[54]}
   );
   gpc606_5 gpc251 (
      {stage0_19[99], stage0_19[100], stage0_19[101], stage0_19[102], stage0_19[103], stage0_19[104]},
      {stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65], stage0_21[66], stage0_21[67]},
      {stage1_23[9],stage1_22[25],stage1_21[27],stage1_20[41],stage1_19[55]}
   );
   gpc606_5 gpc252 (
      {stage0_19[105], stage0_19[106], stage0_19[107], stage0_19[108], stage0_19[109], stage0_19[110]},
      {stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71], stage0_21[72], stage0_21[73]},
      {stage1_23[10],stage1_22[26],stage1_21[28],stage1_20[42],stage1_19[56]}
   );
   gpc606_5 gpc253 (
      {stage0_19[111], stage0_19[112], stage0_19[113], stage0_19[114], stage0_19[115], stage0_19[116]},
      {stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77], stage0_21[78], stage0_21[79]},
      {stage1_23[11],stage1_22[27],stage1_21[29],stage1_20[43],stage1_19[57]}
   );
   gpc606_5 gpc254 (
      {stage0_19[117], stage0_19[118], stage0_19[119], stage0_19[120], stage0_19[121], stage0_19[122]},
      {stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83], stage0_21[84], stage0_21[85]},
      {stage1_23[12],stage1_22[28],stage1_21[30],stage1_20[44],stage1_19[58]}
   );
   gpc606_5 gpc255 (
      {stage0_19[123], stage0_19[124], stage0_19[125], stage0_19[126], stage0_19[127], stage0_19[128]},
      {stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89], stage0_21[90], stage0_21[91]},
      {stage1_23[13],stage1_22[29],stage1_21[31],stage1_20[45],stage1_19[59]}
   );
   gpc606_5 gpc256 (
      {stage0_19[129], stage0_19[130], stage0_19[131], stage0_19[132], stage0_19[133], stage0_19[134]},
      {stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95], stage0_21[96], stage0_21[97]},
      {stage1_23[14],stage1_22[30],stage1_21[32],stage1_20[46],stage1_19[60]}
   );
   gpc606_5 gpc257 (
      {stage0_19[135], stage0_19[136], stage0_19[137], stage0_19[138], stage0_19[139], stage0_19[140]},
      {stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101], stage0_21[102], stage0_21[103]},
      {stage1_23[15],stage1_22[31],stage1_21[33],stage1_20[47],stage1_19[61]}
   );
   gpc615_5 gpc258 (
      {stage0_19[141], stage0_19[142], stage0_19[143], stage0_19[144], stage0_19[145]},
      {stage0_20[72]},
      {stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107], stage0_21[108], stage0_21[109]},
      {stage1_23[16],stage1_22[32],stage1_21[34],stage1_20[48],stage1_19[62]}
   );
   gpc615_5 gpc259 (
      {stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149], stage0_19[150]},
      {stage0_20[73]},
      {stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113], stage0_21[114], stage0_21[115]},
      {stage1_23[17],stage1_22[33],stage1_21[35],stage1_20[49],stage1_19[63]}
   );
   gpc615_5 gpc260 (
      {stage0_19[151], stage0_19[152], stage0_19[153], stage0_19[154], stage0_19[155]},
      {stage0_20[74]},
      {stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119], stage0_21[120], stage0_21[121]},
      {stage1_23[18],stage1_22[34],stage1_21[36],stage1_20[50],stage1_19[64]}
   );
   gpc606_5 gpc261 (
      {stage0_20[75], stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79], stage0_20[80]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[19],stage1_22[35],stage1_21[37],stage1_20[51]}
   );
   gpc606_5 gpc262 (
      {stage0_20[81], stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85], stage0_20[86]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[20],stage1_22[36],stage1_21[38],stage1_20[52]}
   );
   gpc606_5 gpc263 (
      {stage0_20[87], stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91], stage0_20[92]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[21],stage1_22[37],stage1_21[39],stage1_20[53]}
   );
   gpc606_5 gpc264 (
      {stage0_20[93], stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[22],stage1_22[38],stage1_21[40],stage1_20[54]}
   );
   gpc606_5 gpc265 (
      {stage0_20[99], stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[23],stage1_22[39],stage1_21[41],stage1_20[55]}
   );
   gpc606_5 gpc266 (
      {stage0_20[105], stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109], stage0_20[110]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[24],stage1_22[40],stage1_21[42],stage1_20[56]}
   );
   gpc606_5 gpc267 (
      {stage0_20[111], stage0_20[112], stage0_20[113], stage0_20[114], stage0_20[115], stage0_20[116]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[25],stage1_22[41],stage1_21[43],stage1_20[57]}
   );
   gpc606_5 gpc268 (
      {stage0_20[117], stage0_20[118], stage0_20[119], stage0_20[120], stage0_20[121], stage0_20[122]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[26],stage1_22[42],stage1_21[44],stage1_20[58]}
   );
   gpc606_5 gpc269 (
      {stage0_20[123], stage0_20[124], stage0_20[125], stage0_20[126], stage0_20[127], stage0_20[128]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[27],stage1_22[43],stage1_21[45],stage1_20[59]}
   );
   gpc606_5 gpc270 (
      {stage0_20[129], stage0_20[130], stage0_20[131], stage0_20[132], stage0_20[133], stage0_20[134]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[28],stage1_22[44],stage1_21[46],stage1_20[60]}
   );
   gpc606_5 gpc271 (
      {stage0_20[135], stage0_20[136], stage0_20[137], stage0_20[138], stage0_20[139], stage0_20[140]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[29],stage1_22[45],stage1_21[47],stage1_20[61]}
   );
   gpc606_5 gpc272 (
      {stage0_20[141], stage0_20[142], stage0_20[143], stage0_20[144], stage0_20[145], stage0_20[146]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[30],stage1_22[46],stage1_21[48],stage1_20[62]}
   );
   gpc606_5 gpc273 (
      {stage0_20[147], stage0_20[148], stage0_20[149], stage0_20[150], stage0_20[151], stage0_20[152]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[31],stage1_22[47],stage1_21[49],stage1_20[63]}
   );
   gpc606_5 gpc274 (
      {stage0_20[153], stage0_20[154], stage0_20[155], stage0_20[156], stage0_20[157], stage0_20[158]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[32],stage1_22[48],stage1_21[50],stage1_20[64]}
   );
   gpc615_5 gpc275 (
      {stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125], stage0_21[126]},
      {stage0_22[84]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[14],stage1_23[33],stage1_22[49],stage1_21[51]}
   );
   gpc615_5 gpc276 (
      {stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage0_22[85]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[15],stage1_23[34],stage1_22[50],stage1_21[52]}
   );
   gpc615_5 gpc277 (
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136]},
      {stage0_22[86]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[16],stage1_23[35],stage1_22[51],stage1_21[53]}
   );
   gpc615_5 gpc278 (
      {stage0_21[137], stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141]},
      {stage0_22[87]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[17],stage1_23[36],stage1_22[52],stage1_21[54]}
   );
   gpc615_5 gpc279 (
      {stage0_21[142], stage0_21[143], stage0_21[144], stage0_21[145], stage0_21[146]},
      {stage0_22[88]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[18],stage1_23[37],stage1_22[53],stage1_21[55]}
   );
   gpc606_5 gpc280 (
      {stage0_22[89], stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[5],stage1_24[19],stage1_23[38],stage1_22[54]}
   );
   gpc606_5 gpc281 (
      {stage0_22[95], stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[6],stage1_24[20],stage1_23[39],stage1_22[55]}
   );
   gpc606_5 gpc282 (
      {stage0_22[101], stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[7],stage1_24[21],stage1_23[40],stage1_22[56]}
   );
   gpc606_5 gpc283 (
      {stage0_22[107], stage0_22[108], stage0_22[109], stage0_22[110], stage0_22[111], stage0_22[112]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[8],stage1_24[22],stage1_23[41],stage1_22[57]}
   );
   gpc606_5 gpc284 (
      {stage0_22[113], stage0_22[114], stage0_22[115], stage0_22[116], stage0_22[117], stage0_22[118]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[9],stage1_24[23],stage1_23[42],stage1_22[58]}
   );
   gpc606_5 gpc285 (
      {stage0_22[119], stage0_22[120], stage0_22[121], stage0_22[122], stage0_22[123], stage0_22[124]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[10],stage1_24[24],stage1_23[43],stage1_22[59]}
   );
   gpc606_5 gpc286 (
      {stage0_22[125], stage0_22[126], stage0_22[127], stage0_22[128], stage0_22[129], stage0_22[130]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[11],stage1_24[25],stage1_23[44],stage1_22[60]}
   );
   gpc606_5 gpc287 (
      {stage0_22[131], stage0_22[132], stage0_22[133], stage0_22[134], stage0_22[135], stage0_22[136]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[12],stage1_24[26],stage1_23[45],stage1_22[61]}
   );
   gpc615_5 gpc288 (
      {stage0_22[137], stage0_22[138], stage0_22[139], stage0_22[140], stage0_22[141]},
      {stage0_23[30]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[13],stage1_24[27],stage1_23[46],stage1_22[62]}
   );
   gpc615_5 gpc289 (
      {stage0_22[142], stage0_22[143], stage0_22[144], stage0_22[145], stage0_22[146]},
      {stage0_23[31]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[14],stage1_24[28],stage1_23[47],stage1_22[63]}
   );
   gpc615_5 gpc290 (
      {stage0_22[147], stage0_22[148], stage0_22[149], stage0_22[150], stage0_22[151]},
      {stage0_23[32]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[15],stage1_24[29],stage1_23[48],stage1_22[64]}
   );
   gpc615_5 gpc291 (
      {stage0_22[152], stage0_22[153], stage0_22[154], stage0_22[155], stage0_22[156]},
      {stage0_23[33]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[16],stage1_24[30],stage1_23[49],stage1_22[65]}
   );
   gpc615_5 gpc292 (
      {stage0_22[157], stage0_22[158], stage0_22[159], stage0_22[160], stage0_22[161]},
      {stage0_23[34]},
      {stage0_24[72], stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77]},
      {stage1_26[12],stage1_25[17],stage1_24[31],stage1_23[50],stage1_22[66]}
   );
   gpc606_5 gpc293 (
      {stage0_23[35], stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[13],stage1_25[18],stage1_24[32],stage1_23[51]}
   );
   gpc606_5 gpc294 (
      {stage0_23[41], stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[14],stage1_25[19],stage1_24[33],stage1_23[52]}
   );
   gpc606_5 gpc295 (
      {stage0_23[47], stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[15],stage1_25[20],stage1_24[34],stage1_23[53]}
   );
   gpc606_5 gpc296 (
      {stage0_23[53], stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[16],stage1_25[21],stage1_24[35],stage1_23[54]}
   );
   gpc606_5 gpc297 (
      {stage0_23[59], stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[17],stage1_25[22],stage1_24[36],stage1_23[55]}
   );
   gpc606_5 gpc298 (
      {stage0_23[65], stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[18],stage1_25[23],stage1_24[37],stage1_23[56]}
   );
   gpc606_5 gpc299 (
      {stage0_23[71], stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[19],stage1_25[24],stage1_24[38],stage1_23[57]}
   );
   gpc606_5 gpc300 (
      {stage0_24[78], stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[7],stage1_26[20],stage1_25[25],stage1_24[39]}
   );
   gpc606_5 gpc301 (
      {stage0_24[84], stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[8],stage1_26[21],stage1_25[26],stage1_24[40]}
   );
   gpc606_5 gpc302 (
      {stage0_24[90], stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[9],stage1_26[22],stage1_25[27],stage1_24[41]}
   );
   gpc606_5 gpc303 (
      {stage0_24[96], stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[10],stage1_26[23],stage1_25[28],stage1_24[42]}
   );
   gpc606_5 gpc304 (
      {stage0_24[102], stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[11],stage1_26[24],stage1_25[29],stage1_24[43]}
   );
   gpc606_5 gpc305 (
      {stage0_24[108], stage0_24[109], stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[12],stage1_26[25],stage1_25[30],stage1_24[44]}
   );
   gpc606_5 gpc306 (
      {stage0_24[114], stage0_24[115], stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[13],stage1_26[26],stage1_25[31],stage1_24[45]}
   );
   gpc606_5 gpc307 (
      {stage0_24[120], stage0_24[121], stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[14],stage1_26[27],stage1_25[32],stage1_24[46]}
   );
   gpc615_5 gpc308 (
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46]},
      {stage0_26[48]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[8],stage1_27[15],stage1_26[28],stage1_25[33]}
   );
   gpc615_5 gpc309 (
      {stage0_25[47], stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51]},
      {stage0_26[49]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[9],stage1_27[16],stage1_26[29],stage1_25[34]}
   );
   gpc615_5 gpc310 (
      {stage0_25[52], stage0_25[53], stage0_25[54], stage0_25[55], stage0_25[56]},
      {stage0_26[50]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[10],stage1_27[17],stage1_26[30],stage1_25[35]}
   );
   gpc615_5 gpc311 (
      {stage0_25[57], stage0_25[58], stage0_25[59], stage0_25[60], stage0_25[61]},
      {stage0_26[51]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[11],stage1_27[18],stage1_26[31],stage1_25[36]}
   );
   gpc615_5 gpc312 (
      {stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65], stage0_25[66]},
      {stage0_26[52]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[12],stage1_27[19],stage1_26[32],stage1_25[37]}
   );
   gpc615_5 gpc313 (
      {stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_26[53]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[13],stage1_27[20],stage1_26[33],stage1_25[38]}
   );
   gpc615_5 gpc314 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76]},
      {stage0_26[54]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[14],stage1_27[21],stage1_26[34],stage1_25[39]}
   );
   gpc615_5 gpc315 (
      {stage0_25[77], stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81]},
      {stage0_26[55]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[15],stage1_27[22],stage1_26[35],stage1_25[40]}
   );
   gpc615_5 gpc316 (
      {stage0_25[82], stage0_25[83], stage0_25[84], stage0_25[85], stage0_25[86]},
      {stage0_26[56]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[16],stage1_27[23],stage1_26[36],stage1_25[41]}
   );
   gpc615_5 gpc317 (
      {stage0_25[87], stage0_25[88], stage0_25[89], stage0_25[90], stage0_25[91]},
      {stage0_26[57]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[17],stage1_27[24],stage1_26[37],stage1_25[42]}
   );
   gpc615_5 gpc318 (
      {stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95], stage0_25[96]},
      {stage0_26[58]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[18],stage1_27[25],stage1_26[38],stage1_25[43]}
   );
   gpc615_5 gpc319 (
      {stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_26[59]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[19],stage1_27[26],stage1_26[39],stage1_25[44]}
   );
   gpc615_5 gpc320 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106]},
      {stage0_26[60]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[20],stage1_27[27],stage1_26[40],stage1_25[45]}
   );
   gpc615_5 gpc321 (
      {stage0_25[107], stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111]},
      {stage0_26[61]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[21],stage1_27[28],stage1_26[41],stage1_25[46]}
   );
   gpc615_5 gpc322 (
      {stage0_25[112], stage0_25[113], stage0_25[114], stage0_25[115], stage0_25[116]},
      {stage0_26[62]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[22],stage1_27[29],stage1_26[42],stage1_25[47]}
   );
   gpc615_5 gpc323 (
      {stage0_25[117], stage0_25[118], stage0_25[119], stage0_25[120], stage0_25[121]},
      {stage0_26[63]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[23],stage1_27[30],stage1_26[43],stage1_25[48]}
   );
   gpc615_5 gpc324 (
      {stage0_25[122], stage0_25[123], stage0_25[124], stage0_25[125], stage0_25[126]},
      {stage0_26[64]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[24],stage1_27[31],stage1_26[44],stage1_25[49]}
   );
   gpc606_5 gpc325 (
      {stage0_26[65], stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[17],stage1_28[25],stage1_27[32],stage1_26[45]}
   );
   gpc606_5 gpc326 (
      {stage0_26[71], stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[18],stage1_28[26],stage1_27[33],stage1_26[46]}
   );
   gpc606_5 gpc327 (
      {stage0_26[77], stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[19],stage1_28[27],stage1_27[34],stage1_26[47]}
   );
   gpc606_5 gpc328 (
      {stage0_26[83], stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88]},
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage1_30[3],stage1_29[20],stage1_28[28],stage1_27[35],stage1_26[48]}
   );
   gpc606_5 gpc329 (
      {stage0_26[89], stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94]},
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage1_30[4],stage1_29[21],stage1_28[29],stage1_27[36],stage1_26[49]}
   );
   gpc606_5 gpc330 (
      {stage0_26[95], stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100]},
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage1_30[5],stage1_29[22],stage1_28[30],stage1_27[37],stage1_26[50]}
   );
   gpc606_5 gpc331 (
      {stage0_26[101], stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106]},
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage1_30[6],stage1_29[23],stage1_28[31],stage1_27[38],stage1_26[51]}
   );
   gpc606_5 gpc332 (
      {stage0_26[107], stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112]},
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage1_30[7],stage1_29[24],stage1_28[32],stage1_27[39],stage1_26[52]}
   );
   gpc606_5 gpc333 (
      {stage0_26[113], stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118]},
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage1_30[8],stage1_29[25],stage1_28[33],stage1_27[40],stage1_26[53]}
   );
   gpc606_5 gpc334 (
      {stage0_26[119], stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124]},
      {stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59]},
      {stage1_30[9],stage1_29[26],stage1_28[34],stage1_27[41],stage1_26[54]}
   );
   gpc606_5 gpc335 (
      {stage0_26[125], stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130]},
      {stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65]},
      {stage1_30[10],stage1_29[27],stage1_28[35],stage1_27[42],stage1_26[55]}
   );
   gpc606_5 gpc336 (
      {stage0_26[131], stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136]},
      {stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71]},
      {stage1_30[11],stage1_29[28],stage1_28[36],stage1_27[43],stage1_26[56]}
   );
   gpc606_5 gpc337 (
      {stage0_26[137], stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142]},
      {stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77]},
      {stage1_30[12],stage1_29[29],stage1_28[37],stage1_27[44],stage1_26[57]}
   );
   gpc606_5 gpc338 (
      {stage0_26[143], stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148]},
      {stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83]},
      {stage1_30[13],stage1_29[30],stage1_28[38],stage1_27[45],stage1_26[58]}
   );
   gpc615_5 gpc339 (
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106]},
      {stage0_28[84]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[14],stage1_29[31],stage1_28[39],stage1_27[46]}
   );
   gpc615_5 gpc340 (
      {stage0_27[107], stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111]},
      {stage0_28[85]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[15],stage1_29[32],stage1_28[40],stage1_27[47]}
   );
   gpc615_5 gpc341 (
      {stage0_27[112], stage0_27[113], stage0_27[114], stage0_27[115], stage0_27[116]},
      {stage0_28[86]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[16],stage1_29[33],stage1_28[41],stage1_27[48]}
   );
   gpc615_5 gpc342 (
      {stage0_27[117], stage0_27[118], stage0_27[119], stage0_27[120], stage0_27[121]},
      {stage0_28[87]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[17],stage1_29[34],stage1_28[42],stage1_27[49]}
   );
   gpc615_5 gpc343 (
      {stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125], stage0_27[126]},
      {stage0_28[88]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[18],stage1_29[35],stage1_28[43],stage1_27[50]}
   );
   gpc615_5 gpc344 (
      {stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage0_28[89]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[19],stage1_29[36],stage1_28[44],stage1_27[51]}
   );
   gpc615_5 gpc345 (
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136]},
      {stage0_28[90]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[20],stage1_29[37],stage1_28[45],stage1_27[52]}
   );
   gpc615_5 gpc346 (
      {stage0_27[137], stage0_27[138], stage0_27[139], stage0_27[140], stage0_27[141]},
      {stage0_28[91]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[21],stage1_29[38],stage1_28[46],stage1_27[53]}
   );
   gpc606_5 gpc347 (
      {stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95], stage0_28[96], stage0_28[97]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[8],stage1_30[22],stage1_29[39],stage1_28[47]}
   );
   gpc606_5 gpc348 (
      {stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101], stage0_28[102], stage0_28[103]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[9],stage1_30[23],stage1_29[40],stage1_28[48]}
   );
   gpc606_5 gpc349 (
      {stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107], stage0_28[108], stage0_28[109]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[10],stage1_30[24],stage1_29[41],stage1_28[49]}
   );
   gpc606_5 gpc350 (
      {stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114], stage0_28[115]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[11],stage1_30[25],stage1_29[42],stage1_28[50]}
   );
   gpc606_5 gpc351 (
      {stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120], stage0_28[121]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[12],stage1_30[26],stage1_29[43],stage1_28[51]}
   );
   gpc606_5 gpc352 (
      {stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126], stage0_28[127]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[13],stage1_30[27],stage1_29[44],stage1_28[52]}
   );
   gpc606_5 gpc353 (
      {stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132], stage0_28[133]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[14],stage1_30[28],stage1_29[45],stage1_28[53]}
   );
   gpc606_5 gpc354 (
      {stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138], stage0_28[139]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[15],stage1_30[29],stage1_29[46],stage1_28[54]}
   );
   gpc606_5 gpc355 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[8],stage1_31[16],stage1_30[30],stage1_29[47]}
   );
   gpc606_5 gpc356 (
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[9],stage1_31[17],stage1_30[31],stage1_29[48]}
   );
   gpc606_5 gpc357 (
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[10],stage1_31[18],stage1_30[32],stage1_29[49]}
   );
   gpc606_5 gpc358 (
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[11],stage1_31[19],stage1_30[33],stage1_29[50]}
   );
   gpc606_5 gpc359 (
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[12],stage1_31[20],stage1_30[34],stage1_29[51]}
   );
   gpc606_5 gpc360 (
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[13],stage1_31[21],stage1_30[35],stage1_29[52]}
   );
   gpc606_5 gpc361 (
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[14],stage1_31[22],stage1_30[36],stage1_29[53]}
   );
   gpc606_5 gpc362 (
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[15],stage1_31[23],stage1_30[37],stage1_29[54]}
   );
   gpc606_5 gpc363 (
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[16],stage1_31[24],stage1_30[38],stage1_29[55]}
   );
   gpc606_5 gpc364 (
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[17],stage1_31[25],stage1_30[39],stage1_29[56]}
   );
   gpc606_5 gpc365 (
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[18],stage1_31[26],stage1_30[40],stage1_29[57]}
   );
   gpc606_5 gpc366 (
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[19],stage1_31[27],stage1_30[41],stage1_29[58]}
   );
   gpc606_5 gpc367 (
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[20],stage1_31[28],stage1_30[42],stage1_29[59]}
   );
   gpc606_5 gpc368 (
      {stage0_29[126], stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[21],stage1_31[29],stage1_30[43],stage1_29[60]}
   );
   gpc606_5 gpc369 (
      {stage0_29[132], stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[22],stage1_31[30],stage1_30[44],stage1_29[61]}
   );
   gpc606_5 gpc370 (
      {stage0_29[138], stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[23],stage1_31[31],stage1_30[45],stage1_29[62]}
   );
   gpc1406_5 gpc371 (
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3]},
      {stage0_33[0]},
      {stage1_34[0],stage1_33[16],stage1_32[24],stage1_31[32],stage1_30[46]}
   );
   gpc207_4 gpc372 (
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59], stage0_30[60]},
      {stage0_32[4], stage0_32[5]},
      {stage1_33[17],stage1_32[25],stage1_31[33],stage1_30[47]}
   );
   gpc207_4 gpc373 (
      {stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65], stage0_30[66], stage0_30[67]},
      {stage0_32[6], stage0_32[7]},
      {stage1_33[18],stage1_32[26],stage1_31[34],stage1_30[48]}
   );
   gpc207_4 gpc374 (
      {stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71], stage0_30[72], stage0_30[73], stage0_30[74]},
      {stage0_32[8], stage0_32[9]},
      {stage1_33[19],stage1_32[27],stage1_31[35],stage1_30[49]}
   );
   gpc207_4 gpc375 (
      {stage0_30[75], stage0_30[76], stage0_30[77], stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81]},
      {stage0_32[10], stage0_32[11]},
      {stage1_33[20],stage1_32[28],stage1_31[36],stage1_30[50]}
   );
   gpc207_4 gpc376 (
      {stage0_30[82], stage0_30[83], stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88]},
      {stage0_32[12], stage0_32[13]},
      {stage1_33[21],stage1_32[29],stage1_31[37],stage1_30[51]}
   );
   gpc207_4 gpc377 (
      {stage0_30[89], stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage0_32[14], stage0_32[15]},
      {stage1_33[22],stage1_32[30],stage1_31[38],stage1_30[52]}
   );
   gpc615_5 gpc378 (
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100]},
      {stage0_31[96]},
      {stage0_32[16], stage0_32[17], stage0_32[18], stage0_32[19], stage0_32[20], stage0_32[21]},
      {stage1_34[1],stage1_33[23],stage1_32[31],stage1_31[39],stage1_30[53]}
   );
   gpc615_5 gpc379 (
      {stage0_30[101], stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105]},
      {stage0_31[97]},
      {stage0_32[22], stage0_32[23], stage0_32[24], stage0_32[25], stage0_32[26], stage0_32[27]},
      {stage1_34[2],stage1_33[24],stage1_32[32],stage1_31[40],stage1_30[54]}
   );
   gpc615_5 gpc380 (
      {stage0_30[106], stage0_30[107], stage0_30[108], stage0_30[109], stage0_30[110]},
      {stage0_31[98]},
      {stage0_32[28], stage0_32[29], stage0_32[30], stage0_32[31], stage0_32[32], stage0_32[33]},
      {stage1_34[3],stage1_33[25],stage1_32[33],stage1_31[41],stage1_30[55]}
   );
   gpc615_5 gpc381 (
      {stage0_31[99], stage0_31[100], stage0_31[101], stage0_31[102], stage0_31[103]},
      {stage0_32[34]},
      {stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5], stage0_33[6]},
      {stage1_35[0],stage1_34[4],stage1_33[26],stage1_32[34],stage1_31[42]}
   );
   gpc615_5 gpc382 (
      {stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107], stage0_31[108]},
      {stage0_32[35]},
      {stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11], stage0_33[12]},
      {stage1_35[1],stage1_34[5],stage1_33[27],stage1_32[35],stage1_31[43]}
   );
   gpc606_5 gpc383 (
      {stage0_32[36], stage0_32[37], stage0_32[38], stage0_32[39], stage0_32[40], stage0_32[41]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[2],stage1_34[6],stage1_33[28],stage1_32[36]}
   );
   gpc606_5 gpc384 (
      {stage0_32[42], stage0_32[43], stage0_32[44], stage0_32[45], stage0_32[46], stage0_32[47]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[3],stage1_34[7],stage1_33[29],stage1_32[37]}
   );
   gpc606_5 gpc385 (
      {stage0_32[48], stage0_32[49], stage0_32[50], stage0_32[51], stage0_32[52], stage0_32[53]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[4],stage1_34[8],stage1_33[30],stage1_32[38]}
   );
   gpc615_5 gpc386 (
      {stage0_32[54], stage0_32[55], stage0_32[56], stage0_32[57], stage0_32[58]},
      {stage0_33[13]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[5],stage1_34[9],stage1_33[31],stage1_32[39]}
   );
   gpc615_5 gpc387 (
      {stage0_32[59], stage0_32[60], stage0_32[61], stage0_32[62], stage0_32[63]},
      {stage0_33[14]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[6],stage1_34[10],stage1_33[32],stage1_32[40]}
   );
   gpc615_5 gpc388 (
      {stage0_32[64], stage0_32[65], stage0_32[66], stage0_32[67], stage0_32[68]},
      {stage0_33[15]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[7],stage1_34[11],stage1_33[33],stage1_32[41]}
   );
   gpc615_5 gpc389 (
      {stage0_32[69], stage0_32[70], stage0_32[71], stage0_32[72], stage0_32[73]},
      {stage0_33[16]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[8],stage1_34[12],stage1_33[34],stage1_32[42]}
   );
   gpc615_5 gpc390 (
      {stage0_32[74], stage0_32[75], stage0_32[76], stage0_32[77], stage0_32[78]},
      {stage0_33[17]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[9],stage1_34[13],stage1_33[35],stage1_32[43]}
   );
   gpc615_5 gpc391 (
      {stage0_32[79], stage0_32[80], stage0_32[81], stage0_32[82], stage0_32[83]},
      {stage0_33[18]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[10],stage1_34[14],stage1_33[36],stage1_32[44]}
   );
   gpc615_5 gpc392 (
      {stage0_32[84], stage0_32[85], stage0_32[86], stage0_32[87], stage0_32[88]},
      {stage0_33[19]},
      {stage0_34[54], stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage1_36[9],stage1_35[11],stage1_34[15],stage1_33[37],stage1_32[45]}
   );
   gpc615_5 gpc393 (
      {stage0_32[89], stage0_32[90], stage0_32[91], stage0_32[92], stage0_32[93]},
      {stage0_33[20]},
      {stage0_34[60], stage0_34[61], stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65]},
      {stage1_36[10],stage1_35[12],stage1_34[16],stage1_33[38],stage1_32[46]}
   );
   gpc615_5 gpc394 (
      {stage0_32[94], stage0_32[95], stage0_32[96], stage0_32[97], stage0_32[98]},
      {stage0_33[21]},
      {stage0_34[66], stage0_34[67], stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71]},
      {stage1_36[11],stage1_35[13],stage1_34[17],stage1_33[39],stage1_32[47]}
   );
   gpc615_5 gpc395 (
      {stage0_32[99], stage0_32[100], stage0_32[101], stage0_32[102], stage0_32[103]},
      {stage0_33[22]},
      {stage0_34[72], stage0_34[73], stage0_34[74], stage0_34[75], stage0_34[76], stage0_34[77]},
      {stage1_36[12],stage1_35[14],stage1_34[18],stage1_33[40],stage1_32[48]}
   );
   gpc615_5 gpc396 (
      {stage0_32[104], stage0_32[105], stage0_32[106], stage0_32[107], stage0_32[108]},
      {stage0_33[23]},
      {stage0_34[78], stage0_34[79], stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83]},
      {stage1_36[13],stage1_35[15],stage1_34[19],stage1_33[41],stage1_32[49]}
   );
   gpc615_5 gpc397 (
      {stage0_32[109], stage0_32[110], stage0_32[111], stage0_32[112], stage0_32[113]},
      {stage0_33[24]},
      {stage0_34[84], stage0_34[85], stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89]},
      {stage1_36[14],stage1_35[16],stage1_34[20],stage1_33[42],stage1_32[50]}
   );
   gpc615_5 gpc398 (
      {stage0_32[114], stage0_32[115], stage0_32[116], stage0_32[117], stage0_32[118]},
      {stage0_33[25]},
      {stage0_34[90], stage0_34[91], stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95]},
      {stage1_36[15],stage1_35[17],stage1_34[21],stage1_33[43],stage1_32[51]}
   );
   gpc615_5 gpc399 (
      {stage0_32[119], stage0_32[120], stage0_32[121], stage0_32[122], stage0_32[123]},
      {stage0_33[26]},
      {stage0_34[96], stage0_34[97], stage0_34[98], stage0_34[99], stage0_34[100], stage0_34[101]},
      {stage1_36[16],stage1_35[18],stage1_34[22],stage1_33[44],stage1_32[52]}
   );
   gpc615_5 gpc400 (
      {stage0_32[124], stage0_32[125], stage0_32[126], stage0_32[127], stage0_32[128]},
      {stage0_33[27]},
      {stage0_34[102], stage0_34[103], stage0_34[104], stage0_34[105], stage0_34[106], stage0_34[107]},
      {stage1_36[17],stage1_35[19],stage1_34[23],stage1_33[45],stage1_32[53]}
   );
   gpc606_5 gpc401 (
      {stage0_33[28], stage0_33[29], stage0_33[30], stage0_33[31], stage0_33[32], stage0_33[33]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[18],stage1_35[20],stage1_34[24],stage1_33[46]}
   );
   gpc606_5 gpc402 (
      {stage0_33[34], stage0_33[35], stage0_33[36], stage0_33[37], stage0_33[38], stage0_33[39]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[19],stage1_35[21],stage1_34[25],stage1_33[47]}
   );
   gpc606_5 gpc403 (
      {stage0_33[40], stage0_33[41], stage0_33[42], stage0_33[43], stage0_33[44], stage0_33[45]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[20],stage1_35[22],stage1_34[26],stage1_33[48]}
   );
   gpc606_5 gpc404 (
      {stage0_33[46], stage0_33[47], stage0_33[48], stage0_33[49], stage0_33[50], stage0_33[51]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[21],stage1_35[23],stage1_34[27],stage1_33[49]}
   );
   gpc606_5 gpc405 (
      {stage0_33[52], stage0_33[53], stage0_33[54], stage0_33[55], stage0_33[56], stage0_33[57]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[22],stage1_35[24],stage1_34[28],stage1_33[50]}
   );
   gpc606_5 gpc406 (
      {stage0_33[58], stage0_33[59], stage0_33[60], stage0_33[61], stage0_33[62], stage0_33[63]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[23],stage1_35[25],stage1_34[29],stage1_33[51]}
   );
   gpc606_5 gpc407 (
      {stage0_33[64], stage0_33[65], stage0_33[66], stage0_33[67], stage0_33[68], stage0_33[69]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[24],stage1_35[26],stage1_34[30],stage1_33[52]}
   );
   gpc606_5 gpc408 (
      {stage0_33[70], stage0_33[71], stage0_33[72], stage0_33[73], stage0_33[74], stage0_33[75]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[25],stage1_35[27],stage1_34[31],stage1_33[53]}
   );
   gpc606_5 gpc409 (
      {stage0_33[76], stage0_33[77], stage0_33[78], stage0_33[79], stage0_33[80], stage0_33[81]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[26],stage1_35[28],stage1_34[32],stage1_33[54]}
   );
   gpc606_5 gpc410 (
      {stage0_33[82], stage0_33[83], stage0_33[84], stage0_33[85], stage0_33[86], stage0_33[87]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[27],stage1_35[29],stage1_34[33],stage1_33[55]}
   );
   gpc606_5 gpc411 (
      {stage0_33[88], stage0_33[89], stage0_33[90], stage0_33[91], stage0_33[92], stage0_33[93]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[28],stage1_35[30],stage1_34[34],stage1_33[56]}
   );
   gpc606_5 gpc412 (
      {stage0_33[94], stage0_33[95], stage0_33[96], stage0_33[97], stage0_33[98], stage0_33[99]},
      {stage0_35[66], stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage1_37[11],stage1_36[29],stage1_35[31],stage1_34[35],stage1_33[57]}
   );
   gpc606_5 gpc413 (
      {stage0_33[100], stage0_33[101], stage0_33[102], stage0_33[103], stage0_33[104], stage0_33[105]},
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76], stage0_35[77]},
      {stage1_37[12],stage1_36[30],stage1_35[32],stage1_34[36],stage1_33[58]}
   );
   gpc606_5 gpc414 (
      {stage0_33[106], stage0_33[107], stage0_33[108], stage0_33[109], stage0_33[110], stage0_33[111]},
      {stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81], stage0_35[82], stage0_35[83]},
      {stage1_37[13],stage1_36[31],stage1_35[33],stage1_34[37],stage1_33[59]}
   );
   gpc606_5 gpc415 (
      {stage0_33[112], stage0_33[113], stage0_33[114], stage0_33[115], stage0_33[116], stage0_33[117]},
      {stage0_35[84], stage0_35[85], stage0_35[86], stage0_35[87], stage0_35[88], stage0_35[89]},
      {stage1_37[14],stage1_36[32],stage1_35[34],stage1_34[38],stage1_33[60]}
   );
   gpc606_5 gpc416 (
      {stage0_33[118], stage0_33[119], stage0_33[120], stage0_33[121], stage0_33[122], stage0_33[123]},
      {stage0_35[90], stage0_35[91], stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95]},
      {stage1_37[15],stage1_36[33],stage1_35[35],stage1_34[39],stage1_33[61]}
   );
   gpc606_5 gpc417 (
      {stage0_33[124], stage0_33[125], stage0_33[126], stage0_33[127], stage0_33[128], stage0_33[129]},
      {stage0_35[96], stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage1_37[16],stage1_36[34],stage1_35[36],stage1_34[40],stage1_33[62]}
   );
   gpc606_5 gpc418 (
      {stage0_33[130], stage0_33[131], stage0_33[132], stage0_33[133], stage0_33[134], stage0_33[135]},
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106], stage0_35[107]},
      {stage1_37[17],stage1_36[35],stage1_35[37],stage1_34[41],stage1_33[63]}
   );
   gpc615_5 gpc419 (
      {stage0_34[108], stage0_34[109], stage0_34[110], stage0_34[111], stage0_34[112]},
      {stage0_35[108]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[18],stage1_36[36],stage1_35[38],stage1_34[42]}
   );
   gpc615_5 gpc420 (
      {stage0_34[113], stage0_34[114], stage0_34[115], stage0_34[116], stage0_34[117]},
      {stage0_35[109]},
      {stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11]},
      {stage1_38[1],stage1_37[19],stage1_36[37],stage1_35[39],stage1_34[43]}
   );
   gpc615_5 gpc421 (
      {stage0_34[118], stage0_34[119], stage0_34[120], stage0_34[121], stage0_34[122]},
      {stage0_35[110]},
      {stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16], stage0_36[17]},
      {stage1_38[2],stage1_37[20],stage1_36[38],stage1_35[40],stage1_34[44]}
   );
   gpc615_5 gpc422 (
      {stage0_34[123], stage0_34[124], stage0_34[125], stage0_34[126], stage0_34[127]},
      {stage0_35[111]},
      {stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21], stage0_36[22], stage0_36[23]},
      {stage1_38[3],stage1_37[21],stage1_36[39],stage1_35[41],stage1_34[45]}
   );
   gpc615_5 gpc423 (
      {stage0_34[128], stage0_34[129], stage0_34[130], stage0_34[131], stage0_34[132]},
      {stage0_35[112]},
      {stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27], stage0_36[28], stage0_36[29]},
      {stage1_38[4],stage1_37[22],stage1_36[40],stage1_35[42],stage1_34[46]}
   );
   gpc615_5 gpc424 (
      {stage0_34[133], stage0_34[134], stage0_34[135], stage0_34[136], stage0_34[137]},
      {stage0_35[113]},
      {stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33], stage0_36[34], stage0_36[35]},
      {stage1_38[5],stage1_37[23],stage1_36[41],stage1_35[43],stage1_34[47]}
   );
   gpc615_5 gpc425 (
      {stage0_34[138], stage0_34[139], stage0_34[140], stage0_34[141], stage0_34[142]},
      {stage0_35[114]},
      {stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39], stage0_36[40], stage0_36[41]},
      {stage1_38[6],stage1_37[24],stage1_36[42],stage1_35[44],stage1_34[48]}
   );
   gpc615_5 gpc426 (
      {stage0_34[143], stage0_34[144], stage0_34[145], stage0_34[146], stage0_34[147]},
      {stage0_35[115]},
      {stage0_36[42], stage0_36[43], stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47]},
      {stage1_38[7],stage1_37[25],stage1_36[43],stage1_35[45],stage1_34[49]}
   );
   gpc615_5 gpc427 (
      {stage0_34[148], stage0_34[149], stage0_34[150], stage0_34[151], stage0_34[152]},
      {stage0_35[116]},
      {stage0_36[48], stage0_36[49], stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53]},
      {stage1_38[8],stage1_37[26],stage1_36[44],stage1_35[46],stage1_34[50]}
   );
   gpc615_5 gpc428 (
      {stage0_34[153], stage0_34[154], stage0_34[155], stage0_34[156], stage0_34[157]},
      {stage0_35[117]},
      {stage0_36[54], stage0_36[55], stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59]},
      {stage1_38[9],stage1_37[27],stage1_36[45],stage1_35[47],stage1_34[51]}
   );
   gpc615_5 gpc429 (
      {stage0_35[118], stage0_35[119], stage0_35[120], stage0_35[121], stage0_35[122]},
      {stage0_36[60]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[10],stage1_37[28],stage1_36[46],stage1_35[48]}
   );
   gpc615_5 gpc430 (
      {stage0_35[123], stage0_35[124], stage0_35[125], stage0_35[126], stage0_35[127]},
      {stage0_36[61]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[11],stage1_37[29],stage1_36[47],stage1_35[49]}
   );
   gpc615_5 gpc431 (
      {stage0_35[128], stage0_35[129], stage0_35[130], stage0_35[131], stage0_35[132]},
      {stage0_36[62]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[12],stage1_37[30],stage1_36[48],stage1_35[50]}
   );
   gpc615_5 gpc432 (
      {stage0_35[133], stage0_35[134], stage0_35[135], stage0_35[136], stage0_35[137]},
      {stage0_36[63]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[13],stage1_37[31],stage1_36[49],stage1_35[51]}
   );
   gpc615_5 gpc433 (
      {stage0_35[138], stage0_35[139], stage0_35[140], stage0_35[141], stage0_35[142]},
      {stage0_36[64]},
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage1_39[4],stage1_38[14],stage1_37[32],stage1_36[50],stage1_35[52]}
   );
   gpc615_5 gpc434 (
      {stage0_35[143], stage0_35[144], stage0_35[145], stage0_35[146], stage0_35[147]},
      {stage0_36[65]},
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage1_39[5],stage1_38[15],stage1_37[33],stage1_36[51],stage1_35[53]}
   );
   gpc615_5 gpc435 (
      {stage0_35[148], stage0_35[149], stage0_35[150], stage0_35[151], stage0_35[152]},
      {stage0_36[66]},
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage1_39[6],stage1_38[16],stage1_37[34],stage1_36[52],stage1_35[54]}
   );
   gpc615_5 gpc436 (
      {stage0_35[153], stage0_35[154], stage0_35[155], stage0_35[156], stage0_35[157]},
      {stage0_36[67]},
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage1_39[7],stage1_38[17],stage1_37[35],stage1_36[53],stage1_35[55]}
   );
   gpc606_5 gpc437 (
      {stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71], stage0_36[72], stage0_36[73]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[8],stage1_38[18],stage1_37[36],stage1_36[54]}
   );
   gpc606_5 gpc438 (
      {stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77], stage0_36[78], stage0_36[79]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[9],stage1_38[19],stage1_37[37],stage1_36[55]}
   );
   gpc606_5 gpc439 (
      {stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83], stage0_36[84], stage0_36[85]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[10],stage1_38[20],stage1_37[38],stage1_36[56]}
   );
   gpc606_5 gpc440 (
      {stage0_36[86], stage0_36[87], stage0_36[88], stage0_36[89], stage0_36[90], stage0_36[91]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[11],stage1_38[21],stage1_37[39],stage1_36[57]}
   );
   gpc606_5 gpc441 (
      {stage0_36[92], stage0_36[93], stage0_36[94], stage0_36[95], stage0_36[96], stage0_36[97]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[12],stage1_38[22],stage1_37[40],stage1_36[58]}
   );
   gpc606_5 gpc442 (
      {stage0_36[98], stage0_36[99], stage0_36[100], stage0_36[101], stage0_36[102], stage0_36[103]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[13],stage1_38[23],stage1_37[41],stage1_36[59]}
   );
   gpc606_5 gpc443 (
      {stage0_36[104], stage0_36[105], stage0_36[106], stage0_36[107], stage0_36[108], stage0_36[109]},
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41]},
      {stage1_40[6],stage1_39[14],stage1_38[24],stage1_37[42],stage1_36[60]}
   );
   gpc606_5 gpc444 (
      {stage0_36[110], stage0_36[111], stage0_36[112], stage0_36[113], stage0_36[114], stage0_36[115]},
      {stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47]},
      {stage1_40[7],stage1_39[15],stage1_38[25],stage1_37[43],stage1_36[61]}
   );
   gpc606_5 gpc445 (
      {stage0_36[116], stage0_36[117], stage0_36[118], stage0_36[119], stage0_36[120], stage0_36[121]},
      {stage0_38[48], stage0_38[49], stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53]},
      {stage1_40[8],stage1_39[16],stage1_38[26],stage1_37[44],stage1_36[62]}
   );
   gpc606_5 gpc446 (
      {stage0_36[122], stage0_36[123], stage0_36[124], stage0_36[125], stage0_36[126], stage0_36[127]},
      {stage0_38[54], stage0_38[55], stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59]},
      {stage1_40[9],stage1_39[17],stage1_38[27],stage1_37[45],stage1_36[63]}
   );
   gpc606_5 gpc447 (
      {stage0_36[128], stage0_36[129], stage0_36[130], stage0_36[131], stage0_36[132], stage0_36[133]},
      {stage0_38[60], stage0_38[61], stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65]},
      {stage1_40[10],stage1_39[18],stage1_38[28],stage1_37[46],stage1_36[64]}
   );
   gpc606_5 gpc448 (
      {stage0_36[134], stage0_36[135], stage0_36[136], stage0_36[137], stage0_36[138], stage0_36[139]},
      {stage0_38[66], stage0_38[67], stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71]},
      {stage1_40[11],stage1_39[19],stage1_38[29],stage1_37[47],stage1_36[65]}
   );
   gpc606_5 gpc449 (
      {stage0_36[140], stage0_36[141], stage0_36[142], stage0_36[143], stage0_36[144], stage0_36[145]},
      {stage0_38[72], stage0_38[73], stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77]},
      {stage1_40[12],stage1_39[20],stage1_38[30],stage1_37[48],stage1_36[66]}
   );
   gpc606_5 gpc450 (
      {stage0_37[48], stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[13],stage1_39[21],stage1_38[31],stage1_37[49]}
   );
   gpc606_5 gpc451 (
      {stage0_37[54], stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[14],stage1_39[22],stage1_38[32],stage1_37[50]}
   );
   gpc606_5 gpc452 (
      {stage0_37[60], stage0_37[61], stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[15],stage1_39[23],stage1_38[33],stage1_37[51]}
   );
   gpc606_5 gpc453 (
      {stage0_37[66], stage0_37[67], stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[16],stage1_39[24],stage1_38[34],stage1_37[52]}
   );
   gpc606_5 gpc454 (
      {stage0_37[72], stage0_37[73], stage0_37[74], stage0_37[75], stage0_37[76], stage0_37[77]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[17],stage1_39[25],stage1_38[35],stage1_37[53]}
   );
   gpc606_5 gpc455 (
      {stage0_37[78], stage0_37[79], stage0_37[80], stage0_37[81], stage0_37[82], stage0_37[83]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[18],stage1_39[26],stage1_38[36],stage1_37[54]}
   );
   gpc606_5 gpc456 (
      {stage0_37[84], stage0_37[85], stage0_37[86], stage0_37[87], stage0_37[88], stage0_37[89]},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[19],stage1_39[27],stage1_38[37],stage1_37[55]}
   );
   gpc615_5 gpc457 (
      {stage0_38[78], stage0_38[79], stage0_38[80], stage0_38[81], stage0_38[82]},
      {stage0_39[42]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[7],stage1_40[20],stage1_39[28],stage1_38[38]}
   );
   gpc615_5 gpc458 (
      {stage0_38[83], stage0_38[84], stage0_38[85], stage0_38[86], stage0_38[87]},
      {stage0_39[43]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[8],stage1_40[21],stage1_39[29],stage1_38[39]}
   );
   gpc615_5 gpc459 (
      {stage0_38[88], stage0_38[89], stage0_38[90], stage0_38[91], stage0_38[92]},
      {stage0_39[44]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[9],stage1_40[22],stage1_39[30],stage1_38[40]}
   );
   gpc615_5 gpc460 (
      {stage0_38[93], stage0_38[94], stage0_38[95], stage0_38[96], stage0_38[97]},
      {stage0_39[45]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[10],stage1_40[23],stage1_39[31],stage1_38[41]}
   );
   gpc615_5 gpc461 (
      {stage0_38[98], stage0_38[99], stage0_38[100], stage0_38[101], stage0_38[102]},
      {stage0_39[46]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[11],stage1_40[24],stage1_39[32],stage1_38[42]}
   );
   gpc615_5 gpc462 (
      {stage0_38[103], stage0_38[104], stage0_38[105], stage0_38[106], stage0_38[107]},
      {stage0_39[47]},
      {stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33], stage0_40[34], stage0_40[35]},
      {stage1_42[5],stage1_41[12],stage1_40[25],stage1_39[33],stage1_38[43]}
   );
   gpc615_5 gpc463 (
      {stage0_38[108], stage0_38[109], stage0_38[110], stage0_38[111], stage0_38[112]},
      {stage0_39[48]},
      {stage0_40[36], stage0_40[37], stage0_40[38], stage0_40[39], stage0_40[40], stage0_40[41]},
      {stage1_42[6],stage1_41[13],stage1_40[26],stage1_39[34],stage1_38[44]}
   );
   gpc615_5 gpc464 (
      {stage0_38[113], stage0_38[114], stage0_38[115], stage0_38[116], stage0_38[117]},
      {stage0_39[49]},
      {stage0_40[42], stage0_40[43], stage0_40[44], stage0_40[45], stage0_40[46], stage0_40[47]},
      {stage1_42[7],stage1_41[14],stage1_40[27],stage1_39[35],stage1_38[45]}
   );
   gpc615_5 gpc465 (
      {stage0_38[118], stage0_38[119], stage0_38[120], stage0_38[121], stage0_38[122]},
      {stage0_39[50]},
      {stage0_40[48], stage0_40[49], stage0_40[50], stage0_40[51], stage0_40[52], stage0_40[53]},
      {stage1_42[8],stage1_41[15],stage1_40[28],stage1_39[36],stage1_38[46]}
   );
   gpc615_5 gpc466 (
      {stage0_38[123], stage0_38[124], stage0_38[125], stage0_38[126], stage0_38[127]},
      {stage0_39[51]},
      {stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57], stage0_40[58], stage0_40[59]},
      {stage1_42[9],stage1_41[16],stage1_40[29],stage1_39[37],stage1_38[47]}
   );
   gpc615_5 gpc467 (
      {stage0_38[128], stage0_38[129], stage0_38[130], stage0_38[131], stage0_38[132]},
      {stage0_39[52]},
      {stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63], stage0_40[64], stage0_40[65]},
      {stage1_42[10],stage1_41[17],stage1_40[30],stage1_39[38],stage1_38[48]}
   );
   gpc615_5 gpc468 (
      {stage0_38[133], stage0_38[134], stage0_38[135], stage0_38[136], stage0_38[137]},
      {stage0_39[53]},
      {stage0_40[66], stage0_40[67], stage0_40[68], stage0_40[69], stage0_40[70], stage0_40[71]},
      {stage1_42[11],stage1_41[18],stage1_40[31],stage1_39[39],stage1_38[49]}
   );
   gpc615_5 gpc469 (
      {stage0_38[138], stage0_38[139], stage0_38[140], stage0_38[141], stage0_38[142]},
      {stage0_39[54]},
      {stage0_40[72], stage0_40[73], stage0_40[74], stage0_40[75], stage0_40[76], stage0_40[77]},
      {stage1_42[12],stage1_41[19],stage1_40[32],stage1_39[40],stage1_38[50]}
   );
   gpc615_5 gpc470 (
      {stage0_38[143], stage0_38[144], stage0_38[145], stage0_38[146], stage0_38[147]},
      {stage0_39[55]},
      {stage0_40[78], stage0_40[79], stage0_40[80], stage0_40[81], stage0_40[82], stage0_40[83]},
      {stage1_42[13],stage1_41[20],stage1_40[33],stage1_39[41],stage1_38[51]}
   );
   gpc615_5 gpc471 (
      {stage0_39[56], stage0_39[57], stage0_39[58], stage0_39[59], stage0_39[60]},
      {stage0_40[84]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[14],stage1_41[21],stage1_40[34],stage1_39[42]}
   );
   gpc615_5 gpc472 (
      {stage0_39[61], stage0_39[62], stage0_39[63], stage0_39[64], stage0_39[65]},
      {stage0_40[85]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[15],stage1_41[22],stage1_40[35],stage1_39[43]}
   );
   gpc615_5 gpc473 (
      {stage0_39[66], stage0_39[67], stage0_39[68], stage0_39[69], stage0_39[70]},
      {stage0_40[86]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[16],stage1_41[23],stage1_40[36],stage1_39[44]}
   );
   gpc615_5 gpc474 (
      {stage0_39[71], stage0_39[72], stage0_39[73], stage0_39[74], stage0_39[75]},
      {stage0_40[87]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[17],stage1_41[24],stage1_40[37],stage1_39[45]}
   );
   gpc615_5 gpc475 (
      {stage0_39[76], stage0_39[77], stage0_39[78], stage0_39[79], stage0_39[80]},
      {stage0_40[88]},
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage1_43[4],stage1_42[18],stage1_41[25],stage1_40[38],stage1_39[46]}
   );
   gpc615_5 gpc476 (
      {stage0_39[81], stage0_39[82], stage0_39[83], stage0_39[84], stage0_39[85]},
      {stage0_40[89]},
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage1_43[5],stage1_42[19],stage1_41[26],stage1_40[39],stage1_39[47]}
   );
   gpc615_5 gpc477 (
      {stage0_39[86], stage0_39[87], stage0_39[88], stage0_39[89], stage0_39[90]},
      {stage0_40[90]},
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage1_43[6],stage1_42[20],stage1_41[27],stage1_40[40],stage1_39[48]}
   );
   gpc615_5 gpc478 (
      {stage0_39[91], stage0_39[92], stage0_39[93], stage0_39[94], stage0_39[95]},
      {stage0_40[91]},
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage1_43[7],stage1_42[21],stage1_41[28],stage1_40[41],stage1_39[49]}
   );
   gpc615_5 gpc479 (
      {stage0_39[96], stage0_39[97], stage0_39[98], stage0_39[99], stage0_39[100]},
      {stage0_40[92]},
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage1_43[8],stage1_42[22],stage1_41[29],stage1_40[42],stage1_39[50]}
   );
   gpc615_5 gpc480 (
      {stage0_39[101], stage0_39[102], stage0_39[103], stage0_39[104], stage0_39[105]},
      {stage0_40[93]},
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage1_43[9],stage1_42[23],stage1_41[30],stage1_40[43],stage1_39[51]}
   );
   gpc615_5 gpc481 (
      {stage0_39[106], stage0_39[107], stage0_39[108], stage0_39[109], stage0_39[110]},
      {stage0_40[94]},
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage1_43[10],stage1_42[24],stage1_41[31],stage1_40[44],stage1_39[52]}
   );
   gpc615_5 gpc482 (
      {stage0_39[111], stage0_39[112], stage0_39[113], stage0_39[114], stage0_39[115]},
      {stage0_40[95]},
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage1_43[11],stage1_42[25],stage1_41[32],stage1_40[45],stage1_39[53]}
   );
   gpc615_5 gpc483 (
      {stage0_39[116], stage0_39[117], stage0_39[118], stage0_39[119], stage0_39[120]},
      {stage0_40[96]},
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage1_43[12],stage1_42[26],stage1_41[33],stage1_40[46],stage1_39[54]}
   );
   gpc615_5 gpc484 (
      {stage0_39[121], stage0_39[122], stage0_39[123], stage0_39[124], stage0_39[125]},
      {stage0_40[97]},
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage1_43[13],stage1_42[27],stage1_41[34],stage1_40[47],stage1_39[55]}
   );
   gpc615_5 gpc485 (
      {stage0_39[126], stage0_39[127], stage0_39[128], stage0_39[129], stage0_39[130]},
      {stage0_40[98]},
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage1_43[14],stage1_42[28],stage1_41[35],stage1_40[48],stage1_39[56]}
   );
   gpc615_5 gpc486 (
      {stage0_39[131], stage0_39[132], stage0_39[133], stage0_39[134], stage0_39[135]},
      {stage0_40[99]},
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage1_43[15],stage1_42[29],stage1_41[36],stage1_40[49],stage1_39[57]}
   );
   gpc615_5 gpc487 (
      {stage0_39[136], stage0_39[137], stage0_39[138], stage0_39[139], stage0_39[140]},
      {stage0_40[100]},
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100], stage0_41[101]},
      {stage1_43[16],stage1_42[30],stage1_41[37],stage1_40[50],stage1_39[58]}
   );
   gpc615_5 gpc488 (
      {stage0_39[141], stage0_39[142], stage0_39[143], stage0_39[144], stage0_39[145]},
      {stage0_40[101]},
      {stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105], stage0_41[106], stage0_41[107]},
      {stage1_43[17],stage1_42[31],stage1_41[38],stage1_40[51],stage1_39[59]}
   );
   gpc615_5 gpc489 (
      {stage0_39[146], stage0_39[147], stage0_39[148], stage0_39[149], stage0_39[150]},
      {stage0_40[102]},
      {stage0_41[108], stage0_41[109], stage0_41[110], stage0_41[111], stage0_41[112], stage0_41[113]},
      {stage1_43[18],stage1_42[32],stage1_41[39],stage1_40[52],stage1_39[60]}
   );
   gpc615_5 gpc490 (
      {stage0_39[151], stage0_39[152], stage0_39[153], stage0_39[154], stage0_39[155]},
      {stage0_40[103]},
      {stage0_41[114], stage0_41[115], stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119]},
      {stage1_43[19],stage1_42[33],stage1_41[40],stage1_40[53],stage1_39[61]}
   );
   gpc606_5 gpc491 (
      {stage0_40[104], stage0_40[105], stage0_40[106], stage0_40[107], stage0_40[108], stage0_40[109]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[20],stage1_42[34],stage1_41[41],stage1_40[54]}
   );
   gpc606_5 gpc492 (
      {stage0_40[110], stage0_40[111], stage0_40[112], stage0_40[113], stage0_40[114], stage0_40[115]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[21],stage1_42[35],stage1_41[42],stage1_40[55]}
   );
   gpc606_5 gpc493 (
      {stage0_40[116], stage0_40[117], stage0_40[118], stage0_40[119], stage0_40[120], stage0_40[121]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[22],stage1_42[36],stage1_41[43],stage1_40[56]}
   );
   gpc606_5 gpc494 (
      {stage0_40[122], stage0_40[123], stage0_40[124], stage0_40[125], stage0_40[126], stage0_40[127]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[23],stage1_42[37],stage1_41[44],stage1_40[57]}
   );
   gpc606_5 gpc495 (
      {stage0_40[128], stage0_40[129], stage0_40[130], stage0_40[131], stage0_40[132], stage0_40[133]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[24],stage1_42[38],stage1_41[45],stage1_40[58]}
   );
   gpc606_5 gpc496 (
      {stage0_40[134], stage0_40[135], stage0_40[136], stage0_40[137], stage0_40[138], stage0_40[139]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[25],stage1_42[39],stage1_41[46],stage1_40[59]}
   );
   gpc606_5 gpc497 (
      {stage0_41[120], stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[6],stage1_43[26],stage1_42[40],stage1_41[47]}
   );
   gpc606_5 gpc498 (
      {stage0_41[126], stage0_41[127], stage0_41[128], stage0_41[129], stage0_41[130], stage0_41[131]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[7],stage1_43[27],stage1_42[41],stage1_41[48]}
   );
   gpc606_5 gpc499 (
      {stage0_41[132], stage0_41[133], stage0_41[134], stage0_41[135], stage0_41[136], stage0_41[137]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[8],stage1_43[28],stage1_42[42],stage1_41[49]}
   );
   gpc606_5 gpc500 (
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[3],stage1_44[9],stage1_43[29],stage1_42[43]}
   );
   gpc606_5 gpc501 (
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[4],stage1_44[10],stage1_43[30],stage1_42[44]}
   );
   gpc606_5 gpc502 (
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[5],stage1_44[11],stage1_43[31],stage1_42[45]}
   );
   gpc606_5 gpc503 (
      {stage0_42[54], stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[6],stage1_44[12],stage1_43[32],stage1_42[46]}
   );
   gpc606_5 gpc504 (
      {stage0_42[60], stage0_42[61], stage0_42[62], stage0_42[63], stage0_42[64], stage0_42[65]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[7],stage1_44[13],stage1_43[33],stage1_42[47]}
   );
   gpc615_5 gpc505 (
      {stage0_42[66], stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70]},
      {stage0_43[18]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[8],stage1_44[14],stage1_43[34],stage1_42[48]}
   );
   gpc615_5 gpc506 (
      {stage0_42[71], stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75]},
      {stage0_43[19]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[9],stage1_44[15],stage1_43[35],stage1_42[49]}
   );
   gpc615_5 gpc507 (
      {stage0_42[76], stage0_42[77], stage0_42[78], stage0_42[79], stage0_42[80]},
      {stage0_43[20]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[10],stage1_44[16],stage1_43[36],stage1_42[50]}
   );
   gpc615_5 gpc508 (
      {stage0_42[81], stage0_42[82], stage0_42[83], stage0_42[84], stage0_42[85]},
      {stage0_43[21]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[11],stage1_44[17],stage1_43[37],stage1_42[51]}
   );
   gpc615_5 gpc509 (
      {stage0_42[86], stage0_42[87], stage0_42[88], stage0_42[89], stage0_42[90]},
      {stage0_43[22]},
      {stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57], stage0_44[58], stage0_44[59]},
      {stage1_46[9],stage1_45[12],stage1_44[18],stage1_43[38],stage1_42[52]}
   );
   gpc615_5 gpc510 (
      {stage0_42[91], stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95]},
      {stage0_43[23]},
      {stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64], stage0_44[65]},
      {stage1_46[10],stage1_45[13],stage1_44[19],stage1_43[39],stage1_42[53]}
   );
   gpc615_5 gpc511 (
      {stage0_42[96], stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100]},
      {stage0_43[24]},
      {stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70], stage0_44[71]},
      {stage1_46[11],stage1_45[14],stage1_44[20],stage1_43[40],stage1_42[54]}
   );
   gpc615_5 gpc512 (
      {stage0_42[101], stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105]},
      {stage0_43[25]},
      {stage0_44[72], stage0_44[73], stage0_44[74], stage0_44[75], stage0_44[76], stage0_44[77]},
      {stage1_46[12],stage1_45[15],stage1_44[21],stage1_43[41],stage1_42[55]}
   );
   gpc615_5 gpc513 (
      {stage0_42[106], stage0_42[107], stage0_42[108], stage0_42[109], stage0_42[110]},
      {stage0_43[26]},
      {stage0_44[78], stage0_44[79], stage0_44[80], stage0_44[81], stage0_44[82], stage0_44[83]},
      {stage1_46[13],stage1_45[16],stage1_44[22],stage1_43[42],stage1_42[56]}
   );
   gpc615_5 gpc514 (
      {stage0_42[111], stage0_42[112], stage0_42[113], stage0_42[114], stage0_42[115]},
      {stage0_43[27]},
      {stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88], stage0_44[89]},
      {stage1_46[14],stage1_45[17],stage1_44[23],stage1_43[43],stage1_42[57]}
   );
   gpc615_5 gpc515 (
      {stage0_42[116], stage0_42[117], stage0_42[118], stage0_42[119], stage0_42[120]},
      {stage0_43[28]},
      {stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94], stage0_44[95]},
      {stage1_46[15],stage1_45[18],stage1_44[24],stage1_43[44],stage1_42[58]}
   );
   gpc615_5 gpc516 (
      {stage0_42[121], stage0_42[122], stage0_42[123], stage0_42[124], stage0_42[125]},
      {stage0_43[29]},
      {stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100], stage0_44[101]},
      {stage1_46[16],stage1_45[19],stage1_44[25],stage1_43[45],stage1_42[59]}
   );
   gpc606_5 gpc517 (
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[17],stage1_45[20],stage1_44[26],stage1_43[46]}
   );
   gpc606_5 gpc518 (
      {stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39], stage0_43[40], stage0_43[41]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[18],stage1_45[21],stage1_44[27],stage1_43[47]}
   );
   gpc606_5 gpc519 (
      {stage0_43[42], stage0_43[43], stage0_43[44], stage0_43[45], stage0_43[46], stage0_43[47]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[19],stage1_45[22],stage1_44[28],stage1_43[48]}
   );
   gpc606_5 gpc520 (
      {stage0_43[48], stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[20],stage1_45[23],stage1_44[29],stage1_43[49]}
   );
   gpc606_5 gpc521 (
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58], stage0_43[59]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[21],stage1_45[24],stage1_44[30],stage1_43[50]}
   );
   gpc606_5 gpc522 (
      {stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63], stage0_43[64], stage0_43[65]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[22],stage1_45[25],stage1_44[31],stage1_43[51]}
   );
   gpc606_5 gpc523 (
      {stage0_43[66], stage0_43[67], stage0_43[68], stage0_43[69], stage0_43[70], stage0_43[71]},
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage1_47[6],stage1_46[23],stage1_45[26],stage1_44[32],stage1_43[52]}
   );
   gpc606_5 gpc524 (
      {stage0_43[72], stage0_43[73], stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77]},
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage1_47[7],stage1_46[24],stage1_45[27],stage1_44[33],stage1_43[53]}
   );
   gpc606_5 gpc525 (
      {stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106], stage0_44[107]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[8],stage1_46[25],stage1_45[28],stage1_44[34]}
   );
   gpc606_5 gpc526 (
      {stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112], stage0_44[113]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[9],stage1_46[26],stage1_45[29],stage1_44[35]}
   );
   gpc606_5 gpc527 (
      {stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118], stage0_44[119]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[10],stage1_46[27],stage1_45[30],stage1_44[36]}
   );
   gpc606_5 gpc528 (
      {stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124], stage0_44[125]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[11],stage1_46[28],stage1_45[31],stage1_44[37]}
   );
   gpc606_5 gpc529 (
      {stage0_44[126], stage0_44[127], stage0_44[128], stage0_44[129], stage0_44[130], stage0_44[131]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[12],stage1_46[29],stage1_45[32],stage1_44[38]}
   );
   gpc606_5 gpc530 (
      {stage0_44[132], stage0_44[133], stage0_44[134], stage0_44[135], stage0_44[136], stage0_44[137]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[13],stage1_46[30],stage1_45[33],stage1_44[39]}
   );
   gpc606_5 gpc531 (
      {stage0_44[138], stage0_44[139], stage0_44[140], stage0_44[141], stage0_44[142], stage0_44[143]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[14],stage1_46[31],stage1_45[34],stage1_44[40]}
   );
   gpc606_5 gpc532 (
      {stage0_44[144], stage0_44[145], stage0_44[146], stage0_44[147], stage0_44[148], stage0_44[149]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[15],stage1_46[32],stage1_45[35],stage1_44[41]}
   );
   gpc615_5 gpc533 (
      {stage0_44[150], stage0_44[151], stage0_44[152], stage0_44[153], stage0_44[154]},
      {stage0_45[48]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[16],stage1_46[33],stage1_45[36],stage1_44[42]}
   );
   gpc615_5 gpc534 (
      {stage0_44[155], stage0_44[156], stage0_44[157], stage0_44[158], stage0_44[159]},
      {stage0_45[49]},
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage1_48[9],stage1_47[17],stage1_46[34],stage1_45[37],stage1_44[43]}
   );
   gpc606_5 gpc535 (
      {stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53], stage0_45[54], stage0_45[55]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[10],stage1_47[18],stage1_46[35],stage1_45[38]}
   );
   gpc615_5 gpc536 (
      {stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59], stage0_45[60]},
      {stage0_46[60]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[11],stage1_47[19],stage1_46[36],stage1_45[39]}
   );
   gpc615_5 gpc537 (
      {stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage0_46[61]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[12],stage1_47[20],stage1_46[37],stage1_45[40]}
   );
   gpc615_5 gpc538 (
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70]},
      {stage0_46[62]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[13],stage1_47[21],stage1_46[38],stage1_45[41]}
   );
   gpc615_5 gpc539 (
      {stage0_45[71], stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75]},
      {stage0_46[63]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[14],stage1_47[22],stage1_46[39],stage1_45[42]}
   );
   gpc615_5 gpc540 (
      {stage0_45[76], stage0_45[77], stage0_45[78], stage0_45[79], stage0_45[80]},
      {stage0_46[64]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[15],stage1_47[23],stage1_46[40],stage1_45[43]}
   );
   gpc615_5 gpc541 (
      {stage0_45[81], stage0_45[82], stage0_45[83], stage0_45[84], stage0_45[85]},
      {stage0_46[65]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[16],stage1_47[24],stage1_46[41],stage1_45[44]}
   );
   gpc615_5 gpc542 (
      {stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89], stage0_45[90]},
      {stage0_46[66]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[17],stage1_47[25],stage1_46[42],stage1_45[45]}
   );
   gpc615_5 gpc543 (
      {stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage0_46[67]},
      {stage0_47[48], stage0_47[49], stage0_47[50], stage0_47[51], stage0_47[52], stage0_47[53]},
      {stage1_49[8],stage1_48[18],stage1_47[26],stage1_46[43],stage1_45[46]}
   );
   gpc615_5 gpc544 (
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100]},
      {stage0_46[68]},
      {stage0_47[54], stage0_47[55], stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59]},
      {stage1_49[9],stage1_48[19],stage1_47[27],stage1_46[44],stage1_45[47]}
   );
   gpc615_5 gpc545 (
      {stage0_45[101], stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105]},
      {stage0_46[69]},
      {stage0_47[60], stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65]},
      {stage1_49[10],stage1_48[20],stage1_47[28],stage1_46[45],stage1_45[48]}
   );
   gpc615_5 gpc546 (
      {stage0_45[106], stage0_45[107], stage0_45[108], stage0_45[109], stage0_45[110]},
      {stage0_46[70]},
      {stage0_47[66], stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71]},
      {stage1_49[11],stage1_48[21],stage1_47[29],stage1_46[46],stage1_45[49]}
   );
   gpc615_5 gpc547 (
      {stage0_45[111], stage0_45[112], stage0_45[113], stage0_45[114], stage0_45[115]},
      {stage0_46[71]},
      {stage0_47[72], stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage1_49[12],stage1_48[22],stage1_47[30],stage1_46[47],stage1_45[50]}
   );
   gpc615_5 gpc548 (
      {stage0_45[116], stage0_45[117], stage0_45[118], stage0_45[119], stage0_45[120]},
      {stage0_46[72]},
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82], stage0_47[83]},
      {stage1_49[13],stage1_48[23],stage1_47[31],stage1_46[48],stage1_45[51]}
   );
   gpc117_4 gpc549 (
      {stage0_46[73], stage0_46[74], stage0_46[75], stage0_46[76], stage0_46[77], stage0_46[78], stage0_46[79]},
      {stage0_47[84]},
      {stage0_48[0]},
      {stage1_49[14],stage1_48[24],stage1_47[32],stage1_46[49]}
   );
   gpc117_4 gpc550 (
      {stage0_46[80], stage0_46[81], stage0_46[82], stage0_46[83], stage0_46[84], stage0_46[85], stage0_46[86]},
      {stage0_47[85]},
      {stage0_48[1]},
      {stage1_49[15],stage1_48[25],stage1_47[33],stage1_46[50]}
   );
   gpc117_4 gpc551 (
      {stage0_46[87], stage0_46[88], stage0_46[89], stage0_46[90], stage0_46[91], stage0_46[92], stage0_46[93]},
      {stage0_47[86]},
      {stage0_48[2]},
      {stage1_49[16],stage1_48[26],stage1_47[34],stage1_46[51]}
   );
   gpc117_4 gpc552 (
      {stage0_46[94], stage0_46[95], stage0_46[96], stage0_46[97], stage0_46[98], stage0_46[99], stage0_46[100]},
      {stage0_47[87]},
      {stage0_48[3]},
      {stage1_49[17],stage1_48[27],stage1_47[35],stage1_46[52]}
   );
   gpc117_4 gpc553 (
      {stage0_46[101], stage0_46[102], stage0_46[103], stage0_46[104], stage0_46[105], stage0_46[106], stage0_46[107]},
      {stage0_47[88]},
      {stage0_48[4]},
      {stage1_49[18],stage1_48[28],stage1_47[36],stage1_46[53]}
   );
   gpc117_4 gpc554 (
      {stage0_46[108], stage0_46[109], stage0_46[110], stage0_46[111], stage0_46[112], stage0_46[113], stage0_46[114]},
      {stage0_47[89]},
      {stage0_48[5]},
      {stage1_49[19],stage1_48[29],stage1_47[37],stage1_46[54]}
   );
   gpc117_4 gpc555 (
      {stage0_46[115], stage0_46[116], stage0_46[117], stage0_46[118], stage0_46[119], stage0_46[120], stage0_46[121]},
      {stage0_47[90]},
      {stage0_48[6]},
      {stage1_49[20],stage1_48[30],stage1_47[38],stage1_46[55]}
   );
   gpc606_5 gpc556 (
      {stage0_46[122], stage0_46[123], stage0_46[124], stage0_46[125], stage0_46[126], stage0_46[127]},
      {stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11], stage0_48[12]},
      {stage1_50[0],stage1_49[21],stage1_48[31],stage1_47[39],stage1_46[56]}
   );
   gpc606_5 gpc557 (
      {stage0_46[128], stage0_46[129], stage0_46[130], stage0_46[131], stage0_46[132], stage0_46[133]},
      {stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17], stage0_48[18]},
      {stage1_50[1],stage1_49[22],stage1_48[32],stage1_47[40],stage1_46[57]}
   );
   gpc606_5 gpc558 (
      {stage0_46[134], stage0_46[135], stage0_46[136], stage0_46[137], stage0_46[138], stage0_46[139]},
      {stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23], stage0_48[24]},
      {stage1_50[2],stage1_49[23],stage1_48[33],stage1_47[41],stage1_46[58]}
   );
   gpc606_5 gpc559 (
      {stage0_46[140], stage0_46[141], stage0_46[142], stage0_46[143], stage0_46[144], stage0_46[145]},
      {stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29], stage0_48[30]},
      {stage1_50[3],stage1_49[24],stage1_48[34],stage1_47[42],stage1_46[59]}
   );
   gpc615_5 gpc560 (
      {stage0_46[146], stage0_46[147], stage0_46[148], stage0_46[149], stage0_46[150]},
      {stage0_47[91]},
      {stage0_48[31], stage0_48[32], stage0_48[33], stage0_48[34], stage0_48[35], stage0_48[36]},
      {stage1_50[4],stage1_49[25],stage1_48[35],stage1_47[43],stage1_46[60]}
   );
   gpc615_5 gpc561 (
      {stage0_46[151], stage0_46[152], stage0_46[153], stage0_46[154], stage0_46[155]},
      {stage0_47[92]},
      {stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41], stage0_48[42]},
      {stage1_50[5],stage1_49[26],stage1_48[36],stage1_47[44],stage1_46[61]}
   );
   gpc615_5 gpc562 (
      {stage0_46[156], stage0_46[157], stage0_46[158], stage0_46[159], stage0_46[160]},
      {stage0_47[93]},
      {stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47], stage0_48[48]},
      {stage1_50[6],stage1_49[27],stage1_48[37],stage1_47[45],stage1_46[62]}
   );
   gpc606_5 gpc563 (
      {stage0_47[94], stage0_47[95], stage0_47[96], stage0_47[97], stage0_47[98], stage0_47[99]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[7],stage1_49[28],stage1_48[38],stage1_47[46]}
   );
   gpc606_5 gpc564 (
      {stage0_47[100], stage0_47[101], stage0_47[102], stage0_47[103], stage0_47[104], stage0_47[105]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[8],stage1_49[29],stage1_48[39],stage1_47[47]}
   );
   gpc606_5 gpc565 (
      {stage0_47[106], stage0_47[107], stage0_47[108], stage0_47[109], stage0_47[110], stage0_47[111]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[9],stage1_49[30],stage1_48[40],stage1_47[48]}
   );
   gpc606_5 gpc566 (
      {stage0_47[112], stage0_47[113], stage0_47[114], stage0_47[115], stage0_47[116], stage0_47[117]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[10],stage1_49[31],stage1_48[41],stage1_47[49]}
   );
   gpc606_5 gpc567 (
      {stage0_47[118], stage0_47[119], stage0_47[120], stage0_47[121], stage0_47[122], stage0_47[123]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[11],stage1_49[32],stage1_48[42],stage1_47[50]}
   );
   gpc606_5 gpc568 (
      {stage0_47[124], stage0_47[125], stage0_47[126], stage0_47[127], stage0_47[128], stage0_47[129]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[12],stage1_49[33],stage1_48[43],stage1_47[51]}
   );
   gpc606_5 gpc569 (
      {stage0_47[130], stage0_47[131], stage0_47[132], stage0_47[133], stage0_47[134], stage0_47[135]},
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage1_51[6],stage1_50[13],stage1_49[34],stage1_48[44],stage1_47[52]}
   );
   gpc606_5 gpc570 (
      {stage0_47[136], stage0_47[137], stage0_47[138], stage0_47[139], stage0_47[140], stage0_47[141]},
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46], stage0_49[47]},
      {stage1_51[7],stage1_50[14],stage1_49[35],stage1_48[45],stage1_47[53]}
   );
   gpc615_5 gpc571 (
      {stage0_47[142], stage0_47[143], stage0_47[144], stage0_47[145], stage0_47[146]},
      {stage0_48[49]},
      {stage0_49[48], stage0_49[49], stage0_49[50], stage0_49[51], stage0_49[52], stage0_49[53]},
      {stage1_51[8],stage1_50[15],stage1_49[36],stage1_48[46],stage1_47[54]}
   );
   gpc615_5 gpc572 (
      {stage0_47[147], stage0_47[148], stage0_47[149], stage0_47[150], stage0_47[151]},
      {stage0_48[50]},
      {stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58], stage0_49[59]},
      {stage1_51[9],stage1_50[16],stage1_49[37],stage1_48[47],stage1_47[55]}
   );
   gpc615_5 gpc573 (
      {stage0_47[152], stage0_47[153], stage0_47[154], stage0_47[155], stage0_47[156]},
      {stage0_48[51]},
      {stage0_49[60], stage0_49[61], stage0_49[62], stage0_49[63], stage0_49[64], stage0_49[65]},
      {stage1_51[10],stage1_50[17],stage1_49[38],stage1_48[48],stage1_47[56]}
   );
   gpc615_5 gpc574 (
      {stage0_47[157], stage0_47[158], stage0_47[159], stage0_47[160], stage0_47[161]},
      {stage0_48[52]},
      {stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70], stage0_49[71]},
      {stage1_51[11],stage1_50[18],stage1_49[39],stage1_48[49],stage1_47[57]}
   );
   gpc606_5 gpc575 (
      {stage0_48[53], stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57], stage0_48[58]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[12],stage1_50[19],stage1_49[40],stage1_48[50]}
   );
   gpc606_5 gpc576 (
      {stage0_48[59], stage0_48[60], stage0_48[61], stage0_48[62], stage0_48[63], stage0_48[64]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[13],stage1_50[20],stage1_49[41],stage1_48[51]}
   );
   gpc606_5 gpc577 (
      {stage0_48[65], stage0_48[66], stage0_48[67], stage0_48[68], stage0_48[69], stage0_48[70]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[14],stage1_50[21],stage1_49[42],stage1_48[52]}
   );
   gpc615_5 gpc578 (
      {stage0_48[71], stage0_48[72], stage0_48[73], stage0_48[74], stage0_48[75]},
      {stage0_49[72]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[15],stage1_50[22],stage1_49[43],stage1_48[53]}
   );
   gpc615_5 gpc579 (
      {stage0_48[76], stage0_48[77], stage0_48[78], stage0_48[79], stage0_48[80]},
      {stage0_49[73]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[16],stage1_50[23],stage1_49[44],stage1_48[54]}
   );
   gpc615_5 gpc580 (
      {stage0_48[81], stage0_48[82], stage0_48[83], stage0_48[84], stage0_48[85]},
      {stage0_49[74]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[17],stage1_50[24],stage1_49[45],stage1_48[55]}
   );
   gpc615_5 gpc581 (
      {stage0_48[86], stage0_48[87], stage0_48[88], stage0_48[89], stage0_48[90]},
      {stage0_49[75]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[18],stage1_50[25],stage1_49[46],stage1_48[56]}
   );
   gpc615_5 gpc582 (
      {stage0_48[91], stage0_48[92], stage0_48[93], stage0_48[94], stage0_48[95]},
      {stage0_49[76]},
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47]},
      {stage1_52[7],stage1_51[19],stage1_50[26],stage1_49[47],stage1_48[57]}
   );
   gpc615_5 gpc583 (
      {stage0_48[96], stage0_48[97], stage0_48[98], stage0_48[99], stage0_48[100]},
      {stage0_49[77]},
      {stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53]},
      {stage1_52[8],stage1_51[20],stage1_50[27],stage1_49[48],stage1_48[58]}
   );
   gpc615_5 gpc584 (
      {stage0_48[101], stage0_48[102], stage0_48[103], stage0_48[104], stage0_48[105]},
      {stage0_49[78]},
      {stage0_50[54], stage0_50[55], stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59]},
      {stage1_52[9],stage1_51[21],stage1_50[28],stage1_49[49],stage1_48[59]}
   );
   gpc615_5 gpc585 (
      {stage0_48[106], stage0_48[107], stage0_48[108], stage0_48[109], stage0_48[110]},
      {stage0_49[79]},
      {stage0_50[60], stage0_50[61], stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65]},
      {stage1_52[10],stage1_51[22],stage1_50[29],stage1_49[50],stage1_48[60]}
   );
   gpc615_5 gpc586 (
      {stage0_48[111], stage0_48[112], stage0_48[113], stage0_48[114], stage0_48[115]},
      {stage0_49[80]},
      {stage0_50[66], stage0_50[67], stage0_50[68], stage0_50[69], stage0_50[70], stage0_50[71]},
      {stage1_52[11],stage1_51[23],stage1_50[30],stage1_49[51],stage1_48[61]}
   );
   gpc615_5 gpc587 (
      {stage0_48[116], stage0_48[117], stage0_48[118], stage0_48[119], stage0_48[120]},
      {stage0_49[81]},
      {stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75], stage0_50[76], stage0_50[77]},
      {stage1_52[12],stage1_51[24],stage1_50[31],stage1_49[52],stage1_48[62]}
   );
   gpc615_5 gpc588 (
      {stage0_48[121], stage0_48[122], stage0_48[123], stage0_48[124], stage0_48[125]},
      {stage0_49[82]},
      {stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81], stage0_50[82], stage0_50[83]},
      {stage1_52[13],stage1_51[25],stage1_50[32],stage1_49[53],stage1_48[63]}
   );
   gpc615_5 gpc589 (
      {stage0_48[126], stage0_48[127], stage0_48[128], stage0_48[129], stage0_48[130]},
      {stage0_49[83]},
      {stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87], stage0_50[88], stage0_50[89]},
      {stage1_52[14],stage1_51[26],stage1_50[33],stage1_49[54],stage1_48[64]}
   );
   gpc615_5 gpc590 (
      {stage0_48[131], stage0_48[132], stage0_48[133], stage0_48[134], stage0_48[135]},
      {stage0_49[84]},
      {stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93], stage0_50[94], stage0_50[95]},
      {stage1_52[15],stage1_51[27],stage1_50[34],stage1_49[55],stage1_48[65]}
   );
   gpc615_5 gpc591 (
      {stage0_48[136], stage0_48[137], stage0_48[138], stage0_48[139], stage0_48[140]},
      {stage0_49[85]},
      {stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99], stage0_50[100], stage0_50[101]},
      {stage1_52[16],stage1_51[28],stage1_50[35],stage1_49[56],stage1_48[66]}
   );
   gpc615_5 gpc592 (
      {stage0_48[141], stage0_48[142], stage0_48[143], stage0_48[144], stage0_48[145]},
      {stage0_49[86]},
      {stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105], stage0_50[106], stage0_50[107]},
      {stage1_52[17],stage1_51[29],stage1_50[36],stage1_49[57],stage1_48[67]}
   );
   gpc615_5 gpc593 (
      {stage0_48[146], stage0_48[147], stage0_48[148], stage0_48[149], stage0_48[150]},
      {stage0_49[87]},
      {stage0_50[108], stage0_50[109], stage0_50[110], stage0_50[111], stage0_50[112], stage0_50[113]},
      {stage1_52[18],stage1_51[30],stage1_50[37],stage1_49[58],stage1_48[68]}
   );
   gpc615_5 gpc594 (
      {stage0_48[151], stage0_48[152], stage0_48[153], stage0_48[154], stage0_48[155]},
      {stage0_49[88]},
      {stage0_50[114], stage0_50[115], stage0_50[116], stage0_50[117], stage0_50[118], stage0_50[119]},
      {stage1_52[19],stage1_51[31],stage1_50[38],stage1_49[59],stage1_48[69]}
   );
   gpc615_5 gpc595 (
      {stage0_48[156], stage0_48[157], stage0_48[158], stage0_48[159], stage0_48[160]},
      {stage0_49[89]},
      {stage0_50[120], stage0_50[121], stage0_50[122], stage0_50[123], stage0_50[124], stage0_50[125]},
      {stage1_52[20],stage1_51[32],stage1_50[39],stage1_49[60],stage1_48[70]}
   );
   gpc606_5 gpc596 (
      {stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94], stage0_49[95]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[21],stage1_51[33],stage1_50[40],stage1_49[61]}
   );
   gpc606_5 gpc597 (
      {stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100], stage0_49[101]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[22],stage1_51[34],stage1_50[41],stage1_49[62]}
   );
   gpc615_5 gpc598 (
      {stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106]},
      {stage0_50[126]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[23],stage1_51[35],stage1_50[42],stage1_49[63]}
   );
   gpc615_5 gpc599 (
      {stage0_49[107], stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111]},
      {stage0_50[127]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[24],stage1_51[36],stage1_50[43],stage1_49[64]}
   );
   gpc615_5 gpc600 (
      {stage0_49[112], stage0_49[113], stage0_49[114], stage0_49[115], stage0_49[116]},
      {stage0_50[128]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[25],stage1_51[37],stage1_50[44],stage1_49[65]}
   );
   gpc615_5 gpc601 (
      {stage0_49[117], stage0_49[118], stage0_49[119], stage0_49[120], stage0_49[121]},
      {stage0_50[129]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[26],stage1_51[38],stage1_50[45],stage1_49[66]}
   );
   gpc615_5 gpc602 (
      {stage0_49[122], stage0_49[123], stage0_49[124], stage0_49[125], stage0_49[126]},
      {stage0_50[130]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[27],stage1_51[39],stage1_50[46],stage1_49[67]}
   );
   gpc615_5 gpc603 (
      {stage0_49[127], stage0_49[128], stage0_49[129], stage0_49[130], stage0_49[131]},
      {stage0_50[131]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[28],stage1_51[40],stage1_50[47],stage1_49[68]}
   );
   gpc615_5 gpc604 (
      {stage0_49[132], stage0_49[133], stage0_49[134], stage0_49[135], stage0_49[136]},
      {stage0_50[132]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[29],stage1_51[41],stage1_50[48],stage1_49[69]}
   );
   gpc615_5 gpc605 (
      {stage0_49[137], stage0_49[138], stage0_49[139], stage0_49[140], stage0_49[141]},
      {stage0_50[133]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[30],stage1_51[42],stage1_50[49],stage1_49[70]}
   );
   gpc615_5 gpc606 (
      {stage0_49[142], stage0_49[143], stage0_49[144], stage0_49[145], stage0_49[146]},
      {stage0_50[134]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[31],stage1_51[43],stage1_50[50],stage1_49[71]}
   );
   gpc606_5 gpc607 (
      {stage0_50[135], stage0_50[136], stage0_50[137], stage0_50[138], stage0_50[139], stage0_50[140]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[11],stage1_52[32],stage1_51[44],stage1_50[51]}
   );
   gpc606_5 gpc608 (
      {stage0_50[141], stage0_50[142], stage0_50[143], stage0_50[144], stage0_50[145], stage0_50[146]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[12],stage1_52[33],stage1_51[45],stage1_50[52]}
   );
   gpc606_5 gpc609 (
      {stage0_50[147], stage0_50[148], stage0_50[149], stage0_50[150], stage0_50[151], stage0_50[152]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[13],stage1_52[34],stage1_51[46],stage1_50[53]}
   );
   gpc606_5 gpc610 (
      {stage0_50[153], stage0_50[154], stage0_50[155], stage0_50[156], stage0_50[157], stage0_50[158]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[14],stage1_52[35],stage1_51[47],stage1_50[54]}
   );
   gpc606_5 gpc611 (
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[4],stage1_53[15],stage1_52[36],stage1_51[48]}
   );
   gpc606_5 gpc612 (
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[5],stage1_53[16],stage1_52[37],stage1_51[49]}
   );
   gpc606_5 gpc613 (
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[6],stage1_53[17],stage1_52[38],stage1_51[50]}
   );
   gpc606_5 gpc614 (
      {stage0_51[84], stage0_51[85], stage0_51[86], stage0_51[87], stage0_51[88], stage0_51[89]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[7],stage1_53[18],stage1_52[39],stage1_51[51]}
   );
   gpc606_5 gpc615 (
      {stage0_51[90], stage0_51[91], stage0_51[92], stage0_51[93], stage0_51[94], stage0_51[95]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[8],stage1_53[19],stage1_52[40],stage1_51[52]}
   );
   gpc606_5 gpc616 (
      {stage0_51[96], stage0_51[97], stage0_51[98], stage0_51[99], stage0_51[100], stage0_51[101]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[9],stage1_53[20],stage1_52[41],stage1_51[53]}
   );
   gpc606_5 gpc617 (
      {stage0_51[102], stage0_51[103], stage0_51[104], stage0_51[105], stage0_51[106], stage0_51[107]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[10],stage1_53[21],stage1_52[42],stage1_51[54]}
   );
   gpc606_5 gpc618 (
      {stage0_51[108], stage0_51[109], stage0_51[110], stage0_51[111], stage0_51[112], stage0_51[113]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[11],stage1_53[22],stage1_52[43],stage1_51[55]}
   );
   gpc606_5 gpc619 (
      {stage0_51[114], stage0_51[115], stage0_51[116], stage0_51[117], stage0_51[118], stage0_51[119]},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[12],stage1_53[23],stage1_52[44],stage1_51[56]}
   );
   gpc606_5 gpc620 (
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124], stage0_51[125]},
      {stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57], stage0_53[58], stage0_53[59]},
      {stage1_55[9],stage1_54[13],stage1_53[24],stage1_52[45],stage1_51[57]}
   );
   gpc606_5 gpc621 (
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[10],stage1_54[14],stage1_53[25],stage1_52[46]}
   );
   gpc606_5 gpc622 (
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[11],stage1_54[15],stage1_53[26],stage1_52[47]}
   );
   gpc606_5 gpc623 (
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[12],stage1_54[16],stage1_53[27],stage1_52[48]}
   );
   gpc606_5 gpc624 (
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[13],stage1_54[17],stage1_53[28],stage1_52[49]}
   );
   gpc606_5 gpc625 (
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[14],stage1_54[18],stage1_53[29],stage1_52[50]}
   );
   gpc606_5 gpc626 (
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[15],stage1_54[19],stage1_53[30],stage1_52[51]}
   );
   gpc606_5 gpc627 (
      {stage0_52[60], stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[16],stage1_54[20],stage1_53[31],stage1_52[52]}
   );
   gpc606_5 gpc628 (
      {stage0_52[66], stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[17],stage1_54[21],stage1_53[32],stage1_52[53]}
   );
   gpc606_5 gpc629 (
      {stage0_52[72], stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[18],stage1_54[22],stage1_53[33],stage1_52[54]}
   );
   gpc606_5 gpc630 (
      {stage0_52[78], stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[19],stage1_54[23],stage1_53[34],stage1_52[55]}
   );
   gpc606_5 gpc631 (
      {stage0_52[84], stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[20],stage1_54[24],stage1_53[35],stage1_52[56]}
   );
   gpc606_5 gpc632 (
      {stage0_52[90], stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[21],stage1_54[25],stage1_53[36],stage1_52[57]}
   );
   gpc606_5 gpc633 (
      {stage0_52[96], stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[22],stage1_54[26],stage1_53[37],stage1_52[58]}
   );
   gpc606_5 gpc634 (
      {stage0_52[102], stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[23],stage1_54[27],stage1_53[38],stage1_52[59]}
   );
   gpc606_5 gpc635 (
      {stage0_52[108], stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87], stage0_54[88], stage0_54[89]},
      {stage1_56[14],stage1_55[24],stage1_54[28],stage1_53[39],stage1_52[60]}
   );
   gpc606_5 gpc636 (
      {stage0_52[114], stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119]},
      {stage0_54[90], stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95]},
      {stage1_56[15],stage1_55[25],stage1_54[29],stage1_53[40],stage1_52[61]}
   );
   gpc606_5 gpc637 (
      {stage0_52[120], stage0_52[121], stage0_52[122], stage0_52[123], stage0_52[124], stage0_52[125]},
      {stage0_54[96], stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101]},
      {stage1_56[16],stage1_55[26],stage1_54[30],stage1_53[41],stage1_52[62]}
   );
   gpc606_5 gpc638 (
      {stage0_52[126], stage0_52[127], stage0_52[128], stage0_52[129], stage0_52[130], stage0_52[131]},
      {stage0_54[102], stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage1_56[17],stage1_55[27],stage1_54[31],stage1_53[42],stage1_52[63]}
   );
   gpc606_5 gpc639 (
      {stage0_52[132], stage0_52[133], stage0_52[134], stage0_52[135], stage0_52[136], stage0_52[137]},
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112], stage0_54[113]},
      {stage1_56[18],stage1_55[28],stage1_54[32],stage1_53[43],stage1_52[64]}
   );
   gpc615_5 gpc640 (
      {stage0_52[138], stage0_52[139], stage0_52[140], stage0_52[141], stage0_52[142]},
      {stage0_53[60]},
      {stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117], stage0_54[118], stage0_54[119]},
      {stage1_56[19],stage1_55[29],stage1_54[33],stage1_53[44],stage1_52[65]}
   );
   gpc615_5 gpc641 (
      {stage0_52[143], stage0_52[144], stage0_52[145], stage0_52[146], stage0_52[147]},
      {stage0_53[61]},
      {stage0_54[120], stage0_54[121], stage0_54[122], stage0_54[123], stage0_54[124], stage0_54[125]},
      {stage1_56[20],stage1_55[30],stage1_54[34],stage1_53[45],stage1_52[66]}
   );
   gpc615_5 gpc642 (
      {stage0_52[148], stage0_52[149], stage0_52[150], stage0_52[151], stage0_52[152]},
      {stage0_53[62]},
      {stage0_54[126], stage0_54[127], stage0_54[128], stage0_54[129], stage0_54[130], stage0_54[131]},
      {stage1_56[21],stage1_55[31],stage1_54[35],stage1_53[46],stage1_52[67]}
   );
   gpc606_5 gpc643 (
      {stage0_53[63], stage0_53[64], stage0_53[65], stage0_53[66], stage0_53[67], stage0_53[68]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[22],stage1_55[32],stage1_54[36],stage1_53[47]}
   );
   gpc606_5 gpc644 (
      {stage0_53[69], stage0_53[70], stage0_53[71], stage0_53[72], stage0_53[73], stage0_53[74]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[23],stage1_55[33],stage1_54[37],stage1_53[48]}
   );
   gpc606_5 gpc645 (
      {stage0_53[75], stage0_53[76], stage0_53[77], stage0_53[78], stage0_53[79], stage0_53[80]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[24],stage1_55[34],stage1_54[38],stage1_53[49]}
   );
   gpc606_5 gpc646 (
      {stage0_53[81], stage0_53[82], stage0_53[83], stage0_53[84], stage0_53[85], stage0_53[86]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[25],stage1_55[35],stage1_54[39],stage1_53[50]}
   );
   gpc606_5 gpc647 (
      {stage0_53[87], stage0_53[88], stage0_53[89], stage0_53[90], stage0_53[91], stage0_53[92]},
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage1_57[4],stage1_56[26],stage1_55[36],stage1_54[40],stage1_53[51]}
   );
   gpc606_5 gpc648 (
      {stage0_53[93], stage0_53[94], stage0_53[95], stage0_53[96], stage0_53[97], stage0_53[98]},
      {stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33], stage0_55[34], stage0_55[35]},
      {stage1_57[5],stage1_56[27],stage1_55[37],stage1_54[41],stage1_53[52]}
   );
   gpc606_5 gpc649 (
      {stage0_53[99], stage0_53[100], stage0_53[101], stage0_53[102], stage0_53[103], stage0_53[104]},
      {stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39], stage0_55[40], stage0_55[41]},
      {stage1_57[6],stage1_56[28],stage1_55[38],stage1_54[42],stage1_53[53]}
   );
   gpc606_5 gpc650 (
      {stage0_53[105], stage0_53[106], stage0_53[107], stage0_53[108], stage0_53[109], stage0_53[110]},
      {stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45], stage0_55[46], stage0_55[47]},
      {stage1_57[7],stage1_56[29],stage1_55[39],stage1_54[43],stage1_53[54]}
   );
   gpc606_5 gpc651 (
      {stage0_53[111], stage0_53[112], stage0_53[113], stage0_53[114], stage0_53[115], stage0_53[116]},
      {stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51], stage0_55[52], stage0_55[53]},
      {stage1_57[8],stage1_56[30],stage1_55[40],stage1_54[44],stage1_53[55]}
   );
   gpc606_5 gpc652 (
      {stage0_53[117], stage0_53[118], stage0_53[119], stage0_53[120], stage0_53[121], stage0_53[122]},
      {stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57], stage0_55[58], stage0_55[59]},
      {stage1_57[9],stage1_56[31],stage1_55[41],stage1_54[45],stage1_53[56]}
   );
   gpc606_5 gpc653 (
      {stage0_53[123], stage0_53[124], stage0_53[125], stage0_53[126], stage0_53[127], stage0_53[128]},
      {stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63], stage0_55[64], stage0_55[65]},
      {stage1_57[10],stage1_56[32],stage1_55[42],stage1_54[46],stage1_53[57]}
   );
   gpc606_5 gpc654 (
      {stage0_53[129], stage0_53[130], stage0_53[131], stage0_53[132], stage0_53[133], stage0_53[134]},
      {stage0_55[66], stage0_55[67], stage0_55[68], stage0_55[69], stage0_55[70], stage0_55[71]},
      {stage1_57[11],stage1_56[33],stage1_55[43],stage1_54[47],stage1_53[58]}
   );
   gpc606_5 gpc655 (
      {stage0_53[135], stage0_53[136], stage0_53[137], stage0_53[138], stage0_53[139], stage0_53[140]},
      {stage0_55[72], stage0_55[73], stage0_55[74], stage0_55[75], stage0_55[76], stage0_55[77]},
      {stage1_57[12],stage1_56[34],stage1_55[44],stage1_54[48],stage1_53[59]}
   );
   gpc606_5 gpc656 (
      {stage0_53[141], stage0_53[142], stage0_53[143], stage0_53[144], stage0_53[145], stage0_53[146]},
      {stage0_55[78], stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83]},
      {stage1_57[13],stage1_56[35],stage1_55[45],stage1_54[49],stage1_53[60]}
   );
   gpc606_5 gpc657 (
      {stage0_53[147], stage0_53[148], stage0_53[149], stage0_53[150], stage0_53[151], stage0_53[152]},
      {stage0_55[84], stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89]},
      {stage1_57[14],stage1_56[36],stage1_55[46],stage1_54[50],stage1_53[61]}
   );
   gpc606_5 gpc658 (
      {stage0_53[153], stage0_53[154], stage0_53[155], stage0_53[156], stage0_53[157], stage0_53[158]},
      {stage0_55[90], stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95]},
      {stage1_57[15],stage1_56[37],stage1_55[47],stage1_54[51],stage1_53[62]}
   );
   gpc615_5 gpc659 (
      {stage0_54[132], stage0_54[133], stage0_54[134], stage0_54[135], stage0_54[136]},
      {stage0_55[96]},
      {stage0_56[0], stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5]},
      {stage1_58[0],stage1_57[16],stage1_56[38],stage1_55[48],stage1_54[52]}
   );
   gpc615_5 gpc660 (
      {stage0_54[137], stage0_54[138], stage0_54[139], stage0_54[140], stage0_54[141]},
      {stage0_55[97]},
      {stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11]},
      {stage1_58[1],stage1_57[17],stage1_56[39],stage1_55[49],stage1_54[53]}
   );
   gpc615_5 gpc661 (
      {stage0_54[142], stage0_54[143], stage0_54[144], stage0_54[145], stage0_54[146]},
      {stage0_55[98]},
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage1_58[2],stage1_57[18],stage1_56[40],stage1_55[50],stage1_54[54]}
   );
   gpc615_5 gpc662 (
      {stage0_54[147], stage0_54[148], stage0_54[149], stage0_54[150], stage0_54[151]},
      {stage0_55[99]},
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23]},
      {stage1_58[3],stage1_57[19],stage1_56[41],stage1_55[51],stage1_54[55]}
   );
   gpc615_5 gpc663 (
      {stage0_54[152], stage0_54[153], stage0_54[154], stage0_54[155], stage0_54[156]},
      {stage0_55[100]},
      {stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29]},
      {stage1_58[4],stage1_57[20],stage1_56[42],stage1_55[52],stage1_54[56]}
   );
   gpc615_5 gpc664 (
      {stage0_54[157], stage0_54[158], stage0_54[159], stage0_54[160], stage0_54[161]},
      {stage0_55[101]},
      {stage0_56[30], stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35]},
      {stage1_58[5],stage1_57[21],stage1_56[43],stage1_55[53],stage1_54[57]}
   );
   gpc615_5 gpc665 (
      {stage0_55[102], stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106]},
      {stage0_56[36]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[6],stage1_57[22],stage1_56[44],stage1_55[54]}
   );
   gpc615_5 gpc666 (
      {stage0_55[107], stage0_55[108], stage0_55[109], stage0_55[110], stage0_55[111]},
      {stage0_56[37]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[7],stage1_57[23],stage1_56[45],stage1_55[55]}
   );
   gpc615_5 gpc667 (
      {stage0_55[112], stage0_55[113], stage0_55[114], stage0_55[115], stage0_55[116]},
      {stage0_56[38]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[8],stage1_57[24],stage1_56[46],stage1_55[56]}
   );
   gpc615_5 gpc668 (
      {stage0_55[117], stage0_55[118], stage0_55[119], stage0_55[120], stage0_55[121]},
      {stage0_56[39]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[9],stage1_57[25],stage1_56[47],stage1_55[57]}
   );
   gpc606_5 gpc669 (
      {stage0_56[40], stage0_56[41], stage0_56[42], stage0_56[43], stage0_56[44], stage0_56[45]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[4],stage1_58[10],stage1_57[26],stage1_56[48]}
   );
   gpc606_5 gpc670 (
      {stage0_56[46], stage0_56[47], stage0_56[48], stage0_56[49], stage0_56[50], stage0_56[51]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[5],stage1_58[11],stage1_57[27],stage1_56[49]}
   );
   gpc606_5 gpc671 (
      {stage0_56[52], stage0_56[53], stage0_56[54], stage0_56[55], stage0_56[56], stage0_56[57]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[6],stage1_58[12],stage1_57[28],stage1_56[50]}
   );
   gpc606_5 gpc672 (
      {stage0_56[58], stage0_56[59], stage0_56[60], stage0_56[61], stage0_56[62], stage0_56[63]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[7],stage1_58[13],stage1_57[29],stage1_56[51]}
   );
   gpc606_5 gpc673 (
      {stage0_56[64], stage0_56[65], stage0_56[66], stage0_56[67], stage0_56[68], stage0_56[69]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[8],stage1_58[14],stage1_57[30],stage1_56[52]}
   );
   gpc606_5 gpc674 (
      {stage0_56[70], stage0_56[71], stage0_56[72], stage0_56[73], stage0_56[74], stage0_56[75]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[9],stage1_58[15],stage1_57[31],stage1_56[53]}
   );
   gpc606_5 gpc675 (
      {stage0_56[76], stage0_56[77], stage0_56[78], stage0_56[79], stage0_56[80], stage0_56[81]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[10],stage1_58[16],stage1_57[32],stage1_56[54]}
   );
   gpc606_5 gpc676 (
      {stage0_56[82], stage0_56[83], stage0_56[84], stage0_56[85], stage0_56[86], stage0_56[87]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[11],stage1_58[17],stage1_57[33],stage1_56[55]}
   );
   gpc606_5 gpc677 (
      {stage0_56[88], stage0_56[89], stage0_56[90], stage0_56[91], stage0_56[92], stage0_56[93]},
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage1_60[8],stage1_59[12],stage1_58[18],stage1_57[34],stage1_56[56]}
   );
   gpc606_5 gpc678 (
      {stage0_56[94], stage0_56[95], stage0_56[96], stage0_56[97], stage0_56[98], stage0_56[99]},
      {stage0_58[54], stage0_58[55], stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59]},
      {stage1_60[9],stage1_59[13],stage1_58[19],stage1_57[35],stage1_56[57]}
   );
   gpc606_5 gpc679 (
      {stage0_56[100], stage0_56[101], stage0_56[102], stage0_56[103], stage0_56[104], stage0_56[105]},
      {stage0_58[60], stage0_58[61], stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65]},
      {stage1_60[10],stage1_59[14],stage1_58[20],stage1_57[36],stage1_56[58]}
   );
   gpc606_5 gpc680 (
      {stage0_56[106], stage0_56[107], stage0_56[108], stage0_56[109], stage0_56[110], stage0_56[111]},
      {stage0_58[66], stage0_58[67], stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71]},
      {stage1_60[11],stage1_59[15],stage1_58[21],stage1_57[37],stage1_56[59]}
   );
   gpc606_5 gpc681 (
      {stage0_56[112], stage0_56[113], stage0_56[114], stage0_56[115], stage0_56[116], stage0_56[117]},
      {stage0_58[72], stage0_58[73], stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77]},
      {stage1_60[12],stage1_59[16],stage1_58[22],stage1_57[38],stage1_56[60]}
   );
   gpc606_5 gpc682 (
      {stage0_56[118], stage0_56[119], stage0_56[120], stage0_56[121], stage0_56[122], stage0_56[123]},
      {stage0_58[78], stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage1_60[13],stage1_59[17],stage1_58[23],stage1_57[39],stage1_56[61]}
   );
   gpc606_5 gpc683 (
      {stage0_56[124], stage0_56[125], stage0_56[126], stage0_56[127], stage0_56[128], stage0_56[129]},
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88], stage0_58[89]},
      {stage1_60[14],stage1_59[18],stage1_58[24],stage1_57[40],stage1_56[62]}
   );
   gpc606_5 gpc684 (
      {stage0_56[130], stage0_56[131], stage0_56[132], stage0_56[133], stage0_56[134], stage0_56[135]},
      {stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93], stage0_58[94], stage0_58[95]},
      {stage1_60[15],stage1_59[19],stage1_58[25],stage1_57[41],stage1_56[63]}
   );
   gpc606_5 gpc685 (
      {stage0_56[136], stage0_56[137], stage0_56[138], stage0_56[139], stage0_56[140], stage0_56[141]},
      {stage0_58[96], stage0_58[97], stage0_58[98], stage0_58[99], stage0_58[100], stage0_58[101]},
      {stage1_60[16],stage1_59[20],stage1_58[26],stage1_57[42],stage1_56[64]}
   );
   gpc606_5 gpc686 (
      {stage0_56[142], stage0_56[143], stage0_56[144], stage0_56[145], stage0_56[146], stage0_56[147]},
      {stage0_58[102], stage0_58[103], stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107]},
      {stage1_60[17],stage1_59[21],stage1_58[27],stage1_57[43],stage1_56[65]}
   );
   gpc606_5 gpc687 (
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[18],stage1_59[22],stage1_58[28],stage1_57[44]}
   );
   gpc606_5 gpc688 (
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[19],stage1_59[23],stage1_58[29],stage1_57[45]}
   );
   gpc606_5 gpc689 (
      {stage0_57[36], stage0_57[37], stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[20],stage1_59[24],stage1_58[30],stage1_57[46]}
   );
   gpc606_5 gpc690 (
      {stage0_57[42], stage0_57[43], stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[21],stage1_59[25],stage1_58[31],stage1_57[47]}
   );
   gpc606_5 gpc691 (
      {stage0_57[48], stage0_57[49], stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[22],stage1_59[26],stage1_58[32],stage1_57[48]}
   );
   gpc606_5 gpc692 (
      {stage0_57[54], stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[23],stage1_59[27],stage1_58[33],stage1_57[49]}
   );
   gpc606_5 gpc693 (
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[24],stage1_59[28],stage1_58[34],stage1_57[50]}
   );
   gpc606_5 gpc694 (
      {stage0_57[66], stage0_57[67], stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[25],stage1_59[29],stage1_58[35],stage1_57[51]}
   );
   gpc606_5 gpc695 (
      {stage0_57[72], stage0_57[73], stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[26],stage1_59[30],stage1_58[36],stage1_57[52]}
   );
   gpc606_5 gpc696 (
      {stage0_57[78], stage0_57[79], stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[27],stage1_59[31],stage1_58[37],stage1_57[53]}
   );
   gpc606_5 gpc697 (
      {stage0_57[84], stage0_57[85], stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[28],stage1_59[32],stage1_58[38],stage1_57[54]}
   );
   gpc606_5 gpc698 (
      {stage0_57[90], stage0_57[91], stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[29],stage1_59[33],stage1_58[39],stage1_57[55]}
   );
   gpc606_5 gpc699 (
      {stage0_57[96], stage0_57[97], stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[30],stage1_59[34],stage1_58[40],stage1_57[56]}
   );
   gpc606_5 gpc700 (
      {stage0_57[102], stage0_57[103], stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[31],stage1_59[35],stage1_58[41],stage1_57[57]}
   );
   gpc606_5 gpc701 (
      {stage0_57[108], stage0_57[109], stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[32],stage1_59[36],stage1_58[42],stage1_57[58]}
   );
   gpc606_5 gpc702 (
      {stage0_57[114], stage0_57[115], stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119]},
      {stage0_59[90], stage0_59[91], stage0_59[92], stage0_59[93], stage0_59[94], stage0_59[95]},
      {stage1_61[15],stage1_60[33],stage1_59[37],stage1_58[43],stage1_57[59]}
   );
   gpc606_5 gpc703 (
      {stage0_57[120], stage0_57[121], stage0_57[122], stage0_57[123], stage0_57[124], stage0_57[125]},
      {stage0_59[96], stage0_59[97], stage0_59[98], stage0_59[99], stage0_59[100], stage0_59[101]},
      {stage1_61[16],stage1_60[34],stage1_59[38],stage1_58[44],stage1_57[60]}
   );
   gpc606_5 gpc704 (
      {stage0_57[126], stage0_57[127], stage0_57[128], stage0_57[129], stage0_57[130], stage0_57[131]},
      {stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105], stage0_59[106], stage0_59[107]},
      {stage1_61[17],stage1_60[35],stage1_59[39],stage1_58[45],stage1_57[61]}
   );
   gpc606_5 gpc705 (
      {stage0_57[132], stage0_57[133], stage0_57[134], stage0_57[135], stage0_57[136], stage0_57[137]},
      {stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111], stage0_59[112], stage0_59[113]},
      {stage1_61[18],stage1_60[36],stage1_59[40],stage1_58[46],stage1_57[62]}
   );
   gpc606_5 gpc706 (
      {stage0_57[138], stage0_57[139], stage0_57[140], stage0_57[141], stage0_57[142], stage0_57[143]},
      {stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117], stage0_59[118], stage0_59[119]},
      {stage1_61[19],stage1_60[37],stage1_59[41],stage1_58[47],stage1_57[63]}
   );
   gpc606_5 gpc707 (
      {stage0_57[144], stage0_57[145], stage0_57[146], stage0_57[147], stage0_57[148], stage0_57[149]},
      {stage0_59[120], stage0_59[121], stage0_59[122], stage0_59[123], stage0_59[124], stage0_59[125]},
      {stage1_61[20],stage1_60[38],stage1_59[42],stage1_58[48],stage1_57[64]}
   );
   gpc606_5 gpc708 (
      {stage0_57[150], stage0_57[151], stage0_57[152], stage0_57[153], stage0_57[154], stage0_57[155]},
      {stage0_59[126], stage0_59[127], stage0_59[128], stage0_59[129], stage0_59[130], stage0_59[131]},
      {stage1_61[21],stage1_60[39],stage1_59[43],stage1_58[49],stage1_57[65]}
   );
   gpc606_5 gpc709 (
      {stage0_58[108], stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[22],stage1_60[40],stage1_59[44],stage1_58[50]}
   );
   gpc606_5 gpc710 (
      {stage0_58[114], stage0_58[115], stage0_58[116], stage0_58[117], stage0_58[118], stage0_58[119]},
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage1_62[1],stage1_61[23],stage1_60[41],stage1_59[45],stage1_58[51]}
   );
   gpc606_5 gpc711 (
      {stage0_58[120], stage0_58[121], stage0_58[122], stage0_58[123], stage0_58[124], stage0_58[125]},
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage1_62[2],stage1_61[24],stage1_60[42],stage1_59[46],stage1_58[52]}
   );
   gpc606_5 gpc712 (
      {stage0_58[126], stage0_58[127], stage0_58[128], stage0_58[129], stage0_58[130], stage0_58[131]},
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage1_62[3],stage1_61[25],stage1_60[43],stage1_59[47],stage1_58[53]}
   );
   gpc606_5 gpc713 (
      {stage0_58[132], stage0_58[133], stage0_58[134], stage0_58[135], stage0_58[136], stage0_58[137]},
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage1_62[4],stage1_61[26],stage1_60[44],stage1_59[48],stage1_58[54]}
   );
   gpc606_5 gpc714 (
      {stage0_58[138], stage0_58[139], stage0_58[140], stage0_58[141], stage0_58[142], stage0_58[143]},
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage1_62[5],stage1_61[27],stage1_60[45],stage1_59[49],stage1_58[55]}
   );
   gpc606_5 gpc715 (
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[0],stage1_62[6],stage1_61[28],stage1_60[46]}
   );
   gpc606_5 gpc716 (
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[1],stage1_62[7],stage1_61[29],stage1_60[47]}
   );
   gpc606_5 gpc717 (
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[2],stage1_62[8],stage1_61[30],stage1_60[48]}
   );
   gpc606_5 gpc718 (
      {stage0_60[54], stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[3],stage1_62[9],stage1_61[31],stage1_60[49]}
   );
   gpc606_5 gpc719 (
      {stage0_60[60], stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[4],stage1_62[10],stage1_61[32],stage1_60[50]}
   );
   gpc606_5 gpc720 (
      {stage0_60[66], stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[5],stage1_62[11],stage1_61[33],stage1_60[51]}
   );
   gpc606_5 gpc721 (
      {stage0_60[72], stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[6],stage1_62[12],stage1_61[34],stage1_60[52]}
   );
   gpc606_5 gpc722 (
      {stage0_60[78], stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[7],stage1_62[13],stage1_61[35],stage1_60[53]}
   );
   gpc606_5 gpc723 (
      {stage0_60[84], stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89]},
      {stage0_62[48], stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53]},
      {stage1_64[8],stage1_63[8],stage1_62[14],stage1_61[36],stage1_60[54]}
   );
   gpc606_5 gpc724 (
      {stage0_60[90], stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95]},
      {stage0_62[54], stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59]},
      {stage1_64[9],stage1_63[9],stage1_62[15],stage1_61[37],stage1_60[55]}
   );
   gpc606_5 gpc725 (
      {stage0_60[96], stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101]},
      {stage0_62[60], stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65]},
      {stage1_64[10],stage1_63[10],stage1_62[16],stage1_61[38],stage1_60[56]}
   );
   gpc606_5 gpc726 (
      {stage0_60[102], stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107]},
      {stage0_62[66], stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71]},
      {stage1_64[11],stage1_63[11],stage1_62[17],stage1_61[39],stage1_60[57]}
   );
   gpc606_5 gpc727 (
      {stage0_60[108], stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113]},
      {stage0_62[72], stage0_62[73], stage0_62[74], stage0_62[75], stage0_62[76], stage0_62[77]},
      {stage1_64[12],stage1_63[12],stage1_62[18],stage1_61[40],stage1_60[58]}
   );
   gpc606_5 gpc728 (
      {stage0_60[114], stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119]},
      {stage0_62[78], stage0_62[79], stage0_62[80], stage0_62[81], stage0_62[82], stage0_62[83]},
      {stage1_64[13],stage1_63[13],stage1_62[19],stage1_61[41],stage1_60[59]}
   );
   gpc606_5 gpc729 (
      {stage0_60[120], stage0_60[121], stage0_60[122], stage0_60[123], stage0_60[124], stage0_60[125]},
      {stage0_62[84], stage0_62[85], stage0_62[86], stage0_62[87], stage0_62[88], stage0_62[89]},
      {stage1_64[14],stage1_63[14],stage1_62[20],stage1_61[42],stage1_60[60]}
   );
   gpc606_5 gpc730 (
      {stage0_60[126], stage0_60[127], stage0_60[128], stage0_60[129], stage0_60[130], stage0_60[131]},
      {stage0_62[90], stage0_62[91], stage0_62[92], stage0_62[93], stage0_62[94], stage0_62[95]},
      {stage1_64[15],stage1_63[15],stage1_62[21],stage1_61[43],stage1_60[61]}
   );
   gpc606_5 gpc731 (
      {stage0_60[132], stage0_60[133], stage0_60[134], stage0_60[135], stage0_60[136], stage0_60[137]},
      {stage0_62[96], stage0_62[97], stage0_62[98], stage0_62[99], stage0_62[100], stage0_62[101]},
      {stage1_64[16],stage1_63[16],stage1_62[22],stage1_61[44],stage1_60[62]}
   );
   gpc606_5 gpc732 (
      {stage0_60[138], stage0_60[139], stage0_60[140], stage0_60[141], stage0_60[142], stage0_60[143]},
      {stage0_62[102], stage0_62[103], stage0_62[104], stage0_62[105], stage0_62[106], stage0_62[107]},
      {stage1_64[17],stage1_63[17],stage1_62[23],stage1_61[45],stage1_60[63]}
   );
   gpc606_5 gpc733 (
      {stage0_60[144], stage0_60[145], stage0_60[146], stage0_60[147], stage0_60[148], stage0_60[149]},
      {stage0_62[108], stage0_62[109], stage0_62[110], stage0_62[111], stage0_62[112], stage0_62[113]},
      {stage1_64[18],stage1_63[18],stage1_62[24],stage1_61[46],stage1_60[64]}
   );
   gpc606_5 gpc734 (
      {stage0_60[150], stage0_60[151], stage0_60[152], stage0_60[153], stage0_60[154], stage0_60[155]},
      {stage0_62[114], stage0_62[115], stage0_62[116], stage0_62[117], stage0_62[118], stage0_62[119]},
      {stage1_64[19],stage1_63[19],stage1_62[25],stage1_61[47],stage1_60[65]}
   );
   gpc606_5 gpc735 (
      {stage0_60[156], stage0_60[157], stage0_60[158], stage0_60[159], stage0_60[160], stage0_60[161]},
      {stage0_62[120], stage0_62[121], stage0_62[122], stage0_62[123], stage0_62[124], stage0_62[125]},
      {stage1_64[20],stage1_63[20],stage1_62[26],stage1_61[48],stage1_60[66]}
   );
   gpc606_5 gpc736 (
      {stage0_61[0], stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[21],stage1_63[21],stage1_62[27],stage1_61[49]}
   );
   gpc606_5 gpc737 (
      {stage0_61[6], stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[22],stage1_63[22],stage1_62[28],stage1_61[50]}
   );
   gpc606_5 gpc738 (
      {stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16], stage0_61[17]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[23],stage1_63[23],stage1_62[29],stage1_61[51]}
   );
   gpc606_5 gpc739 (
      {stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21], stage0_61[22], stage0_61[23]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[24],stage1_63[24],stage1_62[30],stage1_61[52]}
   );
   gpc606_5 gpc740 (
      {stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27], stage0_61[28], stage0_61[29]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[25],stage1_63[25],stage1_62[31],stage1_61[53]}
   );
   gpc606_5 gpc741 (
      {stage0_61[30], stage0_61[31], stage0_61[32], stage0_61[33], stage0_61[34], stage0_61[35]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[26],stage1_63[26],stage1_62[32],stage1_61[54]}
   );
   gpc606_5 gpc742 (
      {stage0_61[36], stage0_61[37], stage0_61[38], stage0_61[39], stage0_61[40], stage0_61[41]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[27],stage1_63[27],stage1_62[33],stage1_61[55]}
   );
   gpc606_5 gpc743 (
      {stage0_61[42], stage0_61[43], stage0_61[44], stage0_61[45], stage0_61[46], stage0_61[47]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[28],stage1_63[28],stage1_62[34],stage1_61[56]}
   );
   gpc606_5 gpc744 (
      {stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51], stage0_61[52], stage0_61[53]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[29],stage1_63[29],stage1_62[35],stage1_61[57]}
   );
   gpc606_5 gpc745 (
      {stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57], stage0_61[58], stage0_61[59]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[30],stage1_63[30],stage1_62[36],stage1_61[58]}
   );
   gpc606_5 gpc746 (
      {stage0_61[60], stage0_61[61], stage0_61[62], stage0_61[63], stage0_61[64], stage0_61[65]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[31],stage1_63[31],stage1_62[37],stage1_61[59]}
   );
   gpc606_5 gpc747 (
      {stage0_61[66], stage0_61[67], stage0_61[68], stage0_61[69], stage0_61[70], stage0_61[71]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[32],stage1_63[32],stage1_62[38],stage1_61[60]}
   );
   gpc606_5 gpc748 (
      {stage0_61[72], stage0_61[73], stage0_61[74], stage0_61[75], stage0_61[76], stage0_61[77]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[33],stage1_63[33],stage1_62[39],stage1_61[61]}
   );
   gpc606_5 gpc749 (
      {stage0_61[78], stage0_61[79], stage0_61[80], stage0_61[81], stage0_61[82], stage0_61[83]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[34],stage1_63[34],stage1_62[40],stage1_61[62]}
   );
   gpc606_5 gpc750 (
      {stage0_61[84], stage0_61[85], stage0_61[86], stage0_61[87], stage0_61[88], stage0_61[89]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[35],stage1_63[35],stage1_62[41],stage1_61[63]}
   );
   gpc606_5 gpc751 (
      {stage0_61[90], stage0_61[91], stage0_61[92], stage0_61[93], stage0_61[94], stage0_61[95]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[36],stage1_63[36],stage1_62[42],stage1_61[64]}
   );
   gpc606_5 gpc752 (
      {stage0_61[96], stage0_61[97], stage0_61[98], stage0_61[99], stage0_61[100], stage0_61[101]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[37],stage1_63[37],stage1_62[43],stage1_61[65]}
   );
   gpc606_5 gpc753 (
      {stage0_61[102], stage0_61[103], stage0_61[104], stage0_61[105], stage0_61[106], stage0_61[107]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[38],stage1_63[38],stage1_62[44],stage1_61[66]}
   );
   gpc606_5 gpc754 (
      {stage0_61[108], stage0_61[109], stage0_61[110], stage0_61[111], stage0_61[112], stage0_61[113]},
      {stage0_63[108], stage0_63[109], stage0_63[110], stage0_63[111], stage0_63[112], stage0_63[113]},
      {stage1_65[18],stage1_64[39],stage1_63[39],stage1_62[45],stage1_61[67]}
   );
   gpc606_5 gpc755 (
      {stage0_61[114], stage0_61[115], stage0_61[116], stage0_61[117], stage0_61[118], stage0_61[119]},
      {stage0_63[114], stage0_63[115], stage0_63[116], stage0_63[117], stage0_63[118], stage0_63[119]},
      {stage1_65[19],stage1_64[40],stage1_63[40],stage1_62[46],stage1_61[68]}
   );
   gpc606_5 gpc756 (
      {stage0_61[120], stage0_61[121], stage0_61[122], stage0_61[123], stage0_61[124], stage0_61[125]},
      {stage0_63[120], stage0_63[121], stage0_63[122], stage0_63[123], stage0_63[124], stage0_63[125]},
      {stage1_65[20],stage1_64[41],stage1_63[41],stage1_62[47],stage1_61[69]}
   );
   gpc606_5 gpc757 (
      {stage0_61[126], stage0_61[127], stage0_61[128], stage0_61[129], stage0_61[130], stage0_61[131]},
      {stage0_63[126], stage0_63[127], stage0_63[128], stage0_63[129], stage0_63[130], stage0_63[131]},
      {stage1_65[21],stage1_64[42],stage1_63[42],stage1_62[48],stage1_61[70]}
   );
   gpc606_5 gpc758 (
      {stage0_61[132], stage0_61[133], stage0_61[134], stage0_61[135], stage0_61[136], stage0_61[137]},
      {stage0_63[132], stage0_63[133], stage0_63[134], stage0_63[135], stage0_63[136], stage0_63[137]},
      {stage1_65[22],stage1_64[43],stage1_63[43],stage1_62[49],stage1_61[71]}
   );
   gpc606_5 gpc759 (
      {stage0_61[138], stage0_61[139], stage0_61[140], stage0_61[141], stage0_61[142], stage0_61[143]},
      {stage0_63[138], stage0_63[139], stage0_63[140], stage0_63[141], stage0_63[142], stage0_63[143]},
      {stage1_65[23],stage1_64[44],stage1_63[44],stage1_62[50],stage1_61[72]}
   );
   gpc1_1 gpc760 (
      {stage0_2[160]},
      {stage1_2[53]}
   );
   gpc1_1 gpc761 (
      {stage0_2[161]},
      {stage1_2[54]}
   );
   gpc1_1 gpc762 (
      {stage0_3[139]},
      {stage1_3[61]}
   );
   gpc1_1 gpc763 (
      {stage0_3[140]},
      {stage1_3[62]}
   );
   gpc1_1 gpc764 (
      {stage0_3[141]},
      {stage1_3[63]}
   );
   gpc1_1 gpc765 (
      {stage0_3[142]},
      {stage1_3[64]}
   );
   gpc1_1 gpc766 (
      {stage0_3[143]},
      {stage1_3[65]}
   );
   gpc1_1 gpc767 (
      {stage0_3[144]},
      {stage1_3[66]}
   );
   gpc1_1 gpc768 (
      {stage0_3[145]},
      {stage1_3[67]}
   );
   gpc1_1 gpc769 (
      {stage0_3[146]},
      {stage1_3[68]}
   );
   gpc1_1 gpc770 (
      {stage0_3[147]},
      {stage1_3[69]}
   );
   gpc1_1 gpc771 (
      {stage0_3[148]},
      {stage1_3[70]}
   );
   gpc1_1 gpc772 (
      {stage0_3[149]},
      {stage1_3[71]}
   );
   gpc1_1 gpc773 (
      {stage0_3[150]},
      {stage1_3[72]}
   );
   gpc1_1 gpc774 (
      {stage0_3[151]},
      {stage1_3[73]}
   );
   gpc1_1 gpc775 (
      {stage0_3[152]},
      {stage1_3[74]}
   );
   gpc1_1 gpc776 (
      {stage0_3[153]},
      {stage1_3[75]}
   );
   gpc1_1 gpc777 (
      {stage0_3[154]},
      {stage1_3[76]}
   );
   gpc1_1 gpc778 (
      {stage0_3[155]},
      {stage1_3[77]}
   );
   gpc1_1 gpc779 (
      {stage0_3[156]},
      {stage1_3[78]}
   );
   gpc1_1 gpc780 (
      {stage0_3[157]},
      {stage1_3[79]}
   );
   gpc1_1 gpc781 (
      {stage0_3[158]},
      {stage1_3[80]}
   );
   gpc1_1 gpc782 (
      {stage0_3[159]},
      {stage1_3[81]}
   );
   gpc1_1 gpc783 (
      {stage0_3[160]},
      {stage1_3[82]}
   );
   gpc1_1 gpc784 (
      {stage0_3[161]},
      {stage1_3[83]}
   );
   gpc1_1 gpc785 (
      {stage0_4[158]},
      {stage1_4[79]}
   );
   gpc1_1 gpc786 (
      {stage0_4[159]},
      {stage1_4[80]}
   );
   gpc1_1 gpc787 (
      {stage0_4[160]},
      {stage1_4[81]}
   );
   gpc1_1 gpc788 (
      {stage0_4[161]},
      {stage1_4[82]}
   );
   gpc1_1 gpc789 (
      {stage0_5[102]},
      {stage1_5[55]}
   );
   gpc1_1 gpc790 (
      {stage0_5[103]},
      {stage1_5[56]}
   );
   gpc1_1 gpc791 (
      {stage0_5[104]},
      {stage1_5[57]}
   );
   gpc1_1 gpc792 (
      {stage0_5[105]},
      {stage1_5[58]}
   );
   gpc1_1 gpc793 (
      {stage0_5[106]},
      {stage1_5[59]}
   );
   gpc1_1 gpc794 (
      {stage0_5[107]},
      {stage1_5[60]}
   );
   gpc1_1 gpc795 (
      {stage0_5[108]},
      {stage1_5[61]}
   );
   gpc1_1 gpc796 (
      {stage0_5[109]},
      {stage1_5[62]}
   );
   gpc1_1 gpc797 (
      {stage0_5[110]},
      {stage1_5[63]}
   );
   gpc1_1 gpc798 (
      {stage0_5[111]},
      {stage1_5[64]}
   );
   gpc1_1 gpc799 (
      {stage0_5[112]},
      {stage1_5[65]}
   );
   gpc1_1 gpc800 (
      {stage0_5[113]},
      {stage1_5[66]}
   );
   gpc1_1 gpc801 (
      {stage0_5[114]},
      {stage1_5[67]}
   );
   gpc1_1 gpc802 (
      {stage0_5[115]},
      {stage1_5[68]}
   );
   gpc1_1 gpc803 (
      {stage0_5[116]},
      {stage1_5[69]}
   );
   gpc1_1 gpc804 (
      {stage0_5[117]},
      {stage1_5[70]}
   );
   gpc1_1 gpc805 (
      {stage0_5[118]},
      {stage1_5[71]}
   );
   gpc1_1 gpc806 (
      {stage0_5[119]},
      {stage1_5[72]}
   );
   gpc1_1 gpc807 (
      {stage0_5[120]},
      {stage1_5[73]}
   );
   gpc1_1 gpc808 (
      {stage0_5[121]},
      {stage1_5[74]}
   );
   gpc1_1 gpc809 (
      {stage0_5[122]},
      {stage1_5[75]}
   );
   gpc1_1 gpc810 (
      {stage0_5[123]},
      {stage1_5[76]}
   );
   gpc1_1 gpc811 (
      {stage0_5[124]},
      {stage1_5[77]}
   );
   gpc1_1 gpc812 (
      {stage0_5[125]},
      {stage1_5[78]}
   );
   gpc1_1 gpc813 (
      {stage0_5[126]},
      {stage1_5[79]}
   );
   gpc1_1 gpc814 (
      {stage0_5[127]},
      {stage1_5[80]}
   );
   gpc1_1 gpc815 (
      {stage0_5[128]},
      {stage1_5[81]}
   );
   gpc1_1 gpc816 (
      {stage0_5[129]},
      {stage1_5[82]}
   );
   gpc1_1 gpc817 (
      {stage0_5[130]},
      {stage1_5[83]}
   );
   gpc1_1 gpc818 (
      {stage0_5[131]},
      {stage1_5[84]}
   );
   gpc1_1 gpc819 (
      {stage0_5[132]},
      {stage1_5[85]}
   );
   gpc1_1 gpc820 (
      {stage0_5[133]},
      {stage1_5[86]}
   );
   gpc1_1 gpc821 (
      {stage0_5[134]},
      {stage1_5[87]}
   );
   gpc1_1 gpc822 (
      {stage0_5[135]},
      {stage1_5[88]}
   );
   gpc1_1 gpc823 (
      {stage0_5[136]},
      {stage1_5[89]}
   );
   gpc1_1 gpc824 (
      {stage0_5[137]},
      {stage1_5[90]}
   );
   gpc1_1 gpc825 (
      {stage0_5[138]},
      {stage1_5[91]}
   );
   gpc1_1 gpc826 (
      {stage0_5[139]},
      {stage1_5[92]}
   );
   gpc1_1 gpc827 (
      {stage0_5[140]},
      {stage1_5[93]}
   );
   gpc1_1 gpc828 (
      {stage0_5[141]},
      {stage1_5[94]}
   );
   gpc1_1 gpc829 (
      {stage0_5[142]},
      {stage1_5[95]}
   );
   gpc1_1 gpc830 (
      {stage0_5[143]},
      {stage1_5[96]}
   );
   gpc1_1 gpc831 (
      {stage0_5[144]},
      {stage1_5[97]}
   );
   gpc1_1 gpc832 (
      {stage0_5[145]},
      {stage1_5[98]}
   );
   gpc1_1 gpc833 (
      {stage0_5[146]},
      {stage1_5[99]}
   );
   gpc1_1 gpc834 (
      {stage0_5[147]},
      {stage1_5[100]}
   );
   gpc1_1 gpc835 (
      {stage0_5[148]},
      {stage1_5[101]}
   );
   gpc1_1 gpc836 (
      {stage0_5[149]},
      {stage1_5[102]}
   );
   gpc1_1 gpc837 (
      {stage0_5[150]},
      {stage1_5[103]}
   );
   gpc1_1 gpc838 (
      {stage0_5[151]},
      {stage1_5[104]}
   );
   gpc1_1 gpc839 (
      {stage0_5[152]},
      {stage1_5[105]}
   );
   gpc1_1 gpc840 (
      {stage0_5[153]},
      {stage1_5[106]}
   );
   gpc1_1 gpc841 (
      {stage0_5[154]},
      {stage1_5[107]}
   );
   gpc1_1 gpc842 (
      {stage0_5[155]},
      {stage1_5[108]}
   );
   gpc1_1 gpc843 (
      {stage0_5[156]},
      {stage1_5[109]}
   );
   gpc1_1 gpc844 (
      {stage0_5[157]},
      {stage1_5[110]}
   );
   gpc1_1 gpc845 (
      {stage0_5[158]},
      {stage1_5[111]}
   );
   gpc1_1 gpc846 (
      {stage0_5[159]},
      {stage1_5[112]}
   );
   gpc1_1 gpc847 (
      {stage0_5[160]},
      {stage1_5[113]}
   );
   gpc1_1 gpc848 (
      {stage0_5[161]},
      {stage1_5[114]}
   );
   gpc1_1 gpc849 (
      {stage0_6[154]},
      {stage1_6[50]}
   );
   gpc1_1 gpc850 (
      {stage0_6[155]},
      {stage1_6[51]}
   );
   gpc1_1 gpc851 (
      {stage0_6[156]},
      {stage1_6[52]}
   );
   gpc1_1 gpc852 (
      {stage0_6[157]},
      {stage1_6[53]}
   );
   gpc1_1 gpc853 (
      {stage0_6[158]},
      {stage1_6[54]}
   );
   gpc1_1 gpc854 (
      {stage0_6[159]},
      {stage1_6[55]}
   );
   gpc1_1 gpc855 (
      {stage0_6[160]},
      {stage1_6[56]}
   );
   gpc1_1 gpc856 (
      {stage0_6[161]},
      {stage1_6[57]}
   );
   gpc1_1 gpc857 (
      {stage0_7[153]},
      {stage1_7[62]}
   );
   gpc1_1 gpc858 (
      {stage0_7[154]},
      {stage1_7[63]}
   );
   gpc1_1 gpc859 (
      {stage0_7[155]},
      {stage1_7[64]}
   );
   gpc1_1 gpc860 (
      {stage0_7[156]},
      {stage1_7[65]}
   );
   gpc1_1 gpc861 (
      {stage0_7[157]},
      {stage1_7[66]}
   );
   gpc1_1 gpc862 (
      {stage0_7[158]},
      {stage1_7[67]}
   );
   gpc1_1 gpc863 (
      {stage0_7[159]},
      {stage1_7[68]}
   );
   gpc1_1 gpc864 (
      {stage0_7[160]},
      {stage1_7[69]}
   );
   gpc1_1 gpc865 (
      {stage0_7[161]},
      {stage1_7[70]}
   );
   gpc1_1 gpc866 (
      {stage0_8[149]},
      {stage1_8[68]}
   );
   gpc1_1 gpc867 (
      {stage0_8[150]},
      {stage1_8[69]}
   );
   gpc1_1 gpc868 (
      {stage0_8[151]},
      {stage1_8[70]}
   );
   gpc1_1 gpc869 (
      {stage0_8[152]},
      {stage1_8[71]}
   );
   gpc1_1 gpc870 (
      {stage0_8[153]},
      {stage1_8[72]}
   );
   gpc1_1 gpc871 (
      {stage0_8[154]},
      {stage1_8[73]}
   );
   gpc1_1 gpc872 (
      {stage0_8[155]},
      {stage1_8[74]}
   );
   gpc1_1 gpc873 (
      {stage0_8[156]},
      {stage1_8[75]}
   );
   gpc1_1 gpc874 (
      {stage0_8[157]},
      {stage1_8[76]}
   );
   gpc1_1 gpc875 (
      {stage0_8[158]},
      {stage1_8[77]}
   );
   gpc1_1 gpc876 (
      {stage0_8[159]},
      {stage1_8[78]}
   );
   gpc1_1 gpc877 (
      {stage0_8[160]},
      {stage1_8[79]}
   );
   gpc1_1 gpc878 (
      {stage0_8[161]},
      {stage1_8[80]}
   );
   gpc1_1 gpc879 (
      {stage0_10[124]},
      {stage1_10[57]}
   );
   gpc1_1 gpc880 (
      {stage0_10[125]},
      {stage1_10[58]}
   );
   gpc1_1 gpc881 (
      {stage0_10[126]},
      {stage1_10[59]}
   );
   gpc1_1 gpc882 (
      {stage0_10[127]},
      {stage1_10[60]}
   );
   gpc1_1 gpc883 (
      {stage0_10[128]},
      {stage1_10[61]}
   );
   gpc1_1 gpc884 (
      {stage0_10[129]},
      {stage1_10[62]}
   );
   gpc1_1 gpc885 (
      {stage0_10[130]},
      {stage1_10[63]}
   );
   gpc1_1 gpc886 (
      {stage0_10[131]},
      {stage1_10[64]}
   );
   gpc1_1 gpc887 (
      {stage0_10[132]},
      {stage1_10[65]}
   );
   gpc1_1 gpc888 (
      {stage0_10[133]},
      {stage1_10[66]}
   );
   gpc1_1 gpc889 (
      {stage0_10[134]},
      {stage1_10[67]}
   );
   gpc1_1 gpc890 (
      {stage0_10[135]},
      {stage1_10[68]}
   );
   gpc1_1 gpc891 (
      {stage0_10[136]},
      {stage1_10[69]}
   );
   gpc1_1 gpc892 (
      {stage0_10[137]},
      {stage1_10[70]}
   );
   gpc1_1 gpc893 (
      {stage0_10[138]},
      {stage1_10[71]}
   );
   gpc1_1 gpc894 (
      {stage0_10[139]},
      {stage1_10[72]}
   );
   gpc1_1 gpc895 (
      {stage0_10[140]},
      {stage1_10[73]}
   );
   gpc1_1 gpc896 (
      {stage0_10[141]},
      {stage1_10[74]}
   );
   gpc1_1 gpc897 (
      {stage0_10[142]},
      {stage1_10[75]}
   );
   gpc1_1 gpc898 (
      {stage0_10[143]},
      {stage1_10[76]}
   );
   gpc1_1 gpc899 (
      {stage0_10[144]},
      {stage1_10[77]}
   );
   gpc1_1 gpc900 (
      {stage0_10[145]},
      {stage1_10[78]}
   );
   gpc1_1 gpc901 (
      {stage0_10[146]},
      {stage1_10[79]}
   );
   gpc1_1 gpc902 (
      {stage0_10[147]},
      {stage1_10[80]}
   );
   gpc1_1 gpc903 (
      {stage0_10[148]},
      {stage1_10[81]}
   );
   gpc1_1 gpc904 (
      {stage0_10[149]},
      {stage1_10[82]}
   );
   gpc1_1 gpc905 (
      {stage0_10[150]},
      {stage1_10[83]}
   );
   gpc1_1 gpc906 (
      {stage0_10[151]},
      {stage1_10[84]}
   );
   gpc1_1 gpc907 (
      {stage0_10[152]},
      {stage1_10[85]}
   );
   gpc1_1 gpc908 (
      {stage0_10[153]},
      {stage1_10[86]}
   );
   gpc1_1 gpc909 (
      {stage0_10[154]},
      {stage1_10[87]}
   );
   gpc1_1 gpc910 (
      {stage0_10[155]},
      {stage1_10[88]}
   );
   gpc1_1 gpc911 (
      {stage0_10[156]},
      {stage1_10[89]}
   );
   gpc1_1 gpc912 (
      {stage0_10[157]},
      {stage1_10[90]}
   );
   gpc1_1 gpc913 (
      {stage0_10[158]},
      {stage1_10[91]}
   );
   gpc1_1 gpc914 (
      {stage0_10[159]},
      {stage1_10[92]}
   );
   gpc1_1 gpc915 (
      {stage0_10[160]},
      {stage1_10[93]}
   );
   gpc1_1 gpc916 (
      {stage0_10[161]},
      {stage1_10[94]}
   );
   gpc1_1 gpc917 (
      {stage0_11[144]},
      {stage1_11[63]}
   );
   gpc1_1 gpc918 (
      {stage0_11[145]},
      {stage1_11[64]}
   );
   gpc1_1 gpc919 (
      {stage0_11[146]},
      {stage1_11[65]}
   );
   gpc1_1 gpc920 (
      {stage0_11[147]},
      {stage1_11[66]}
   );
   gpc1_1 gpc921 (
      {stage0_11[148]},
      {stage1_11[67]}
   );
   gpc1_1 gpc922 (
      {stage0_11[149]},
      {stage1_11[68]}
   );
   gpc1_1 gpc923 (
      {stage0_11[150]},
      {stage1_11[69]}
   );
   gpc1_1 gpc924 (
      {stage0_11[151]},
      {stage1_11[70]}
   );
   gpc1_1 gpc925 (
      {stage0_11[152]},
      {stage1_11[71]}
   );
   gpc1_1 gpc926 (
      {stage0_11[153]},
      {stage1_11[72]}
   );
   gpc1_1 gpc927 (
      {stage0_11[154]},
      {stage1_11[73]}
   );
   gpc1_1 gpc928 (
      {stage0_11[155]},
      {stage1_11[74]}
   );
   gpc1_1 gpc929 (
      {stage0_11[156]},
      {stage1_11[75]}
   );
   gpc1_1 gpc930 (
      {stage0_11[157]},
      {stage1_11[76]}
   );
   gpc1_1 gpc931 (
      {stage0_11[158]},
      {stage1_11[77]}
   );
   gpc1_1 gpc932 (
      {stage0_11[159]},
      {stage1_11[78]}
   );
   gpc1_1 gpc933 (
      {stage0_11[160]},
      {stage1_11[79]}
   );
   gpc1_1 gpc934 (
      {stage0_11[161]},
      {stage1_11[80]}
   );
   gpc1_1 gpc935 (
      {stage0_12[158]},
      {stage1_12[63]}
   );
   gpc1_1 gpc936 (
      {stage0_12[159]},
      {stage1_12[64]}
   );
   gpc1_1 gpc937 (
      {stage0_12[160]},
      {stage1_12[65]}
   );
   gpc1_1 gpc938 (
      {stage0_12[161]},
      {stage1_12[66]}
   );
   gpc1_1 gpc939 (
      {stage0_13[132]},
      {stage1_13[57]}
   );
   gpc1_1 gpc940 (
      {stage0_13[133]},
      {stage1_13[58]}
   );
   gpc1_1 gpc941 (
      {stage0_13[134]},
      {stage1_13[59]}
   );
   gpc1_1 gpc942 (
      {stage0_13[135]},
      {stage1_13[60]}
   );
   gpc1_1 gpc943 (
      {stage0_13[136]},
      {stage1_13[61]}
   );
   gpc1_1 gpc944 (
      {stage0_13[137]},
      {stage1_13[62]}
   );
   gpc1_1 gpc945 (
      {stage0_13[138]},
      {stage1_13[63]}
   );
   gpc1_1 gpc946 (
      {stage0_13[139]},
      {stage1_13[64]}
   );
   gpc1_1 gpc947 (
      {stage0_13[140]},
      {stage1_13[65]}
   );
   gpc1_1 gpc948 (
      {stage0_13[141]},
      {stage1_13[66]}
   );
   gpc1_1 gpc949 (
      {stage0_13[142]},
      {stage1_13[67]}
   );
   gpc1_1 gpc950 (
      {stage0_13[143]},
      {stage1_13[68]}
   );
   gpc1_1 gpc951 (
      {stage0_13[144]},
      {stage1_13[69]}
   );
   gpc1_1 gpc952 (
      {stage0_13[145]},
      {stage1_13[70]}
   );
   gpc1_1 gpc953 (
      {stage0_13[146]},
      {stage1_13[71]}
   );
   gpc1_1 gpc954 (
      {stage0_13[147]},
      {stage1_13[72]}
   );
   gpc1_1 gpc955 (
      {stage0_13[148]},
      {stage1_13[73]}
   );
   gpc1_1 gpc956 (
      {stage0_13[149]},
      {stage1_13[74]}
   );
   gpc1_1 gpc957 (
      {stage0_13[150]},
      {stage1_13[75]}
   );
   gpc1_1 gpc958 (
      {stage0_13[151]},
      {stage1_13[76]}
   );
   gpc1_1 gpc959 (
      {stage0_13[152]},
      {stage1_13[77]}
   );
   gpc1_1 gpc960 (
      {stage0_13[153]},
      {stage1_13[78]}
   );
   gpc1_1 gpc961 (
      {stage0_13[154]},
      {stage1_13[79]}
   );
   gpc1_1 gpc962 (
      {stage0_13[155]},
      {stage1_13[80]}
   );
   gpc1_1 gpc963 (
      {stage0_13[156]},
      {stage1_13[81]}
   );
   gpc1_1 gpc964 (
      {stage0_13[157]},
      {stage1_13[82]}
   );
   gpc1_1 gpc965 (
      {stage0_13[158]},
      {stage1_13[83]}
   );
   gpc1_1 gpc966 (
      {stage0_13[159]},
      {stage1_13[84]}
   );
   gpc1_1 gpc967 (
      {stage0_13[160]},
      {stage1_13[85]}
   );
   gpc1_1 gpc968 (
      {stage0_13[161]},
      {stage1_13[86]}
   );
   gpc1_1 gpc969 (
      {stage0_14[158]},
      {stage1_14[58]}
   );
   gpc1_1 gpc970 (
      {stage0_14[159]},
      {stage1_14[59]}
   );
   gpc1_1 gpc971 (
      {stage0_14[160]},
      {stage1_14[60]}
   );
   gpc1_1 gpc972 (
      {stage0_14[161]},
      {stage1_14[61]}
   );
   gpc1_1 gpc973 (
      {stage0_15[128]},
      {stage1_15[64]}
   );
   gpc1_1 gpc974 (
      {stage0_15[129]},
      {stage1_15[65]}
   );
   gpc1_1 gpc975 (
      {stage0_15[130]},
      {stage1_15[66]}
   );
   gpc1_1 gpc976 (
      {stage0_15[131]},
      {stage1_15[67]}
   );
   gpc1_1 gpc977 (
      {stage0_15[132]},
      {stage1_15[68]}
   );
   gpc1_1 gpc978 (
      {stage0_15[133]},
      {stage1_15[69]}
   );
   gpc1_1 gpc979 (
      {stage0_15[134]},
      {stage1_15[70]}
   );
   gpc1_1 gpc980 (
      {stage0_15[135]},
      {stage1_15[71]}
   );
   gpc1_1 gpc981 (
      {stage0_15[136]},
      {stage1_15[72]}
   );
   gpc1_1 gpc982 (
      {stage0_15[137]},
      {stage1_15[73]}
   );
   gpc1_1 gpc983 (
      {stage0_15[138]},
      {stage1_15[74]}
   );
   gpc1_1 gpc984 (
      {stage0_15[139]},
      {stage1_15[75]}
   );
   gpc1_1 gpc985 (
      {stage0_15[140]},
      {stage1_15[76]}
   );
   gpc1_1 gpc986 (
      {stage0_15[141]},
      {stage1_15[77]}
   );
   gpc1_1 gpc987 (
      {stage0_15[142]},
      {stage1_15[78]}
   );
   gpc1_1 gpc988 (
      {stage0_15[143]},
      {stage1_15[79]}
   );
   gpc1_1 gpc989 (
      {stage0_15[144]},
      {stage1_15[80]}
   );
   gpc1_1 gpc990 (
      {stage0_15[145]},
      {stage1_15[81]}
   );
   gpc1_1 gpc991 (
      {stage0_15[146]},
      {stage1_15[82]}
   );
   gpc1_1 gpc992 (
      {stage0_15[147]},
      {stage1_15[83]}
   );
   gpc1_1 gpc993 (
      {stage0_15[148]},
      {stage1_15[84]}
   );
   gpc1_1 gpc994 (
      {stage0_15[149]},
      {stage1_15[85]}
   );
   gpc1_1 gpc995 (
      {stage0_15[150]},
      {stage1_15[86]}
   );
   gpc1_1 gpc996 (
      {stage0_15[151]},
      {stage1_15[87]}
   );
   gpc1_1 gpc997 (
      {stage0_15[152]},
      {stage1_15[88]}
   );
   gpc1_1 gpc998 (
      {stage0_15[153]},
      {stage1_15[89]}
   );
   gpc1_1 gpc999 (
      {stage0_15[154]},
      {stage1_15[90]}
   );
   gpc1_1 gpc1000 (
      {stage0_15[155]},
      {stage1_15[91]}
   );
   gpc1_1 gpc1001 (
      {stage0_15[156]},
      {stage1_15[92]}
   );
   gpc1_1 gpc1002 (
      {stage0_15[157]},
      {stage1_15[93]}
   );
   gpc1_1 gpc1003 (
      {stage0_15[158]},
      {stage1_15[94]}
   );
   gpc1_1 gpc1004 (
      {stage0_15[159]},
      {stage1_15[95]}
   );
   gpc1_1 gpc1005 (
      {stage0_15[160]},
      {stage1_15[96]}
   );
   gpc1_1 gpc1006 (
      {stage0_15[161]},
      {stage1_15[97]}
   );
   gpc1_1 gpc1007 (
      {stage0_16[158]},
      {stage1_16[64]}
   );
   gpc1_1 gpc1008 (
      {stage0_16[159]},
      {stage1_16[65]}
   );
   gpc1_1 gpc1009 (
      {stage0_16[160]},
      {stage1_16[66]}
   );
   gpc1_1 gpc1010 (
      {stage0_16[161]},
      {stage1_16[67]}
   );
   gpc1_1 gpc1011 (
      {stage0_17[96]},
      {stage1_17[48]}
   );
   gpc1_1 gpc1012 (
      {stage0_17[97]},
      {stage1_17[49]}
   );
   gpc1_1 gpc1013 (
      {stage0_17[98]},
      {stage1_17[50]}
   );
   gpc1_1 gpc1014 (
      {stage0_17[99]},
      {stage1_17[51]}
   );
   gpc1_1 gpc1015 (
      {stage0_17[100]},
      {stage1_17[52]}
   );
   gpc1_1 gpc1016 (
      {stage0_17[101]},
      {stage1_17[53]}
   );
   gpc1_1 gpc1017 (
      {stage0_17[102]},
      {stage1_17[54]}
   );
   gpc1_1 gpc1018 (
      {stage0_17[103]},
      {stage1_17[55]}
   );
   gpc1_1 gpc1019 (
      {stage0_17[104]},
      {stage1_17[56]}
   );
   gpc1_1 gpc1020 (
      {stage0_17[105]},
      {stage1_17[57]}
   );
   gpc1_1 gpc1021 (
      {stage0_17[106]},
      {stage1_17[58]}
   );
   gpc1_1 gpc1022 (
      {stage0_17[107]},
      {stage1_17[59]}
   );
   gpc1_1 gpc1023 (
      {stage0_17[108]},
      {stage1_17[60]}
   );
   gpc1_1 gpc1024 (
      {stage0_17[109]},
      {stage1_17[61]}
   );
   gpc1_1 gpc1025 (
      {stage0_17[110]},
      {stage1_17[62]}
   );
   gpc1_1 gpc1026 (
      {stage0_17[111]},
      {stage1_17[63]}
   );
   gpc1_1 gpc1027 (
      {stage0_17[112]},
      {stage1_17[64]}
   );
   gpc1_1 gpc1028 (
      {stage0_17[113]},
      {stage1_17[65]}
   );
   gpc1_1 gpc1029 (
      {stage0_17[114]},
      {stage1_17[66]}
   );
   gpc1_1 gpc1030 (
      {stage0_17[115]},
      {stage1_17[67]}
   );
   gpc1_1 gpc1031 (
      {stage0_17[116]},
      {stage1_17[68]}
   );
   gpc1_1 gpc1032 (
      {stage0_17[117]},
      {stage1_17[69]}
   );
   gpc1_1 gpc1033 (
      {stage0_17[118]},
      {stage1_17[70]}
   );
   gpc1_1 gpc1034 (
      {stage0_17[119]},
      {stage1_17[71]}
   );
   gpc1_1 gpc1035 (
      {stage0_17[120]},
      {stage1_17[72]}
   );
   gpc1_1 gpc1036 (
      {stage0_17[121]},
      {stage1_17[73]}
   );
   gpc1_1 gpc1037 (
      {stage0_17[122]},
      {stage1_17[74]}
   );
   gpc1_1 gpc1038 (
      {stage0_17[123]},
      {stage1_17[75]}
   );
   gpc1_1 gpc1039 (
      {stage0_17[124]},
      {stage1_17[76]}
   );
   gpc1_1 gpc1040 (
      {stage0_17[125]},
      {stage1_17[77]}
   );
   gpc1_1 gpc1041 (
      {stage0_17[126]},
      {stage1_17[78]}
   );
   gpc1_1 gpc1042 (
      {stage0_17[127]},
      {stage1_17[79]}
   );
   gpc1_1 gpc1043 (
      {stage0_17[128]},
      {stage1_17[80]}
   );
   gpc1_1 gpc1044 (
      {stage0_17[129]},
      {stage1_17[81]}
   );
   gpc1_1 gpc1045 (
      {stage0_17[130]},
      {stage1_17[82]}
   );
   gpc1_1 gpc1046 (
      {stage0_17[131]},
      {stage1_17[83]}
   );
   gpc1_1 gpc1047 (
      {stage0_17[132]},
      {stage1_17[84]}
   );
   gpc1_1 gpc1048 (
      {stage0_17[133]},
      {stage1_17[85]}
   );
   gpc1_1 gpc1049 (
      {stage0_17[134]},
      {stage1_17[86]}
   );
   gpc1_1 gpc1050 (
      {stage0_17[135]},
      {stage1_17[87]}
   );
   gpc1_1 gpc1051 (
      {stage0_17[136]},
      {stage1_17[88]}
   );
   gpc1_1 gpc1052 (
      {stage0_17[137]},
      {stage1_17[89]}
   );
   gpc1_1 gpc1053 (
      {stage0_17[138]},
      {stage1_17[90]}
   );
   gpc1_1 gpc1054 (
      {stage0_17[139]},
      {stage1_17[91]}
   );
   gpc1_1 gpc1055 (
      {stage0_17[140]},
      {stage1_17[92]}
   );
   gpc1_1 gpc1056 (
      {stage0_17[141]},
      {stage1_17[93]}
   );
   gpc1_1 gpc1057 (
      {stage0_17[142]},
      {stage1_17[94]}
   );
   gpc1_1 gpc1058 (
      {stage0_17[143]},
      {stage1_17[95]}
   );
   gpc1_1 gpc1059 (
      {stage0_17[144]},
      {stage1_17[96]}
   );
   gpc1_1 gpc1060 (
      {stage0_17[145]},
      {stage1_17[97]}
   );
   gpc1_1 gpc1061 (
      {stage0_17[146]},
      {stage1_17[98]}
   );
   gpc1_1 gpc1062 (
      {stage0_17[147]},
      {stage1_17[99]}
   );
   gpc1_1 gpc1063 (
      {stage0_17[148]},
      {stage1_17[100]}
   );
   gpc1_1 gpc1064 (
      {stage0_17[149]},
      {stage1_17[101]}
   );
   gpc1_1 gpc1065 (
      {stage0_17[150]},
      {stage1_17[102]}
   );
   gpc1_1 gpc1066 (
      {stage0_17[151]},
      {stage1_17[103]}
   );
   gpc1_1 gpc1067 (
      {stage0_17[152]},
      {stage1_17[104]}
   );
   gpc1_1 gpc1068 (
      {stage0_17[153]},
      {stage1_17[105]}
   );
   gpc1_1 gpc1069 (
      {stage0_17[154]},
      {stage1_17[106]}
   );
   gpc1_1 gpc1070 (
      {stage0_17[155]},
      {stage1_17[107]}
   );
   gpc1_1 gpc1071 (
      {stage0_17[156]},
      {stage1_17[108]}
   );
   gpc1_1 gpc1072 (
      {stage0_17[157]},
      {stage1_17[109]}
   );
   gpc1_1 gpc1073 (
      {stage0_17[158]},
      {stage1_17[110]}
   );
   gpc1_1 gpc1074 (
      {stage0_17[159]},
      {stage1_17[111]}
   );
   gpc1_1 gpc1075 (
      {stage0_17[160]},
      {stage1_17[112]}
   );
   gpc1_1 gpc1076 (
      {stage0_17[161]},
      {stage1_17[113]}
   );
   gpc1_1 gpc1077 (
      {stage0_18[151]},
      {stage1_18[52]}
   );
   gpc1_1 gpc1078 (
      {stage0_18[152]},
      {stage1_18[53]}
   );
   gpc1_1 gpc1079 (
      {stage0_18[153]},
      {stage1_18[54]}
   );
   gpc1_1 gpc1080 (
      {stage0_18[154]},
      {stage1_18[55]}
   );
   gpc1_1 gpc1081 (
      {stage0_18[155]},
      {stage1_18[56]}
   );
   gpc1_1 gpc1082 (
      {stage0_18[156]},
      {stage1_18[57]}
   );
   gpc1_1 gpc1083 (
      {stage0_18[157]},
      {stage1_18[58]}
   );
   gpc1_1 gpc1084 (
      {stage0_18[158]},
      {stage1_18[59]}
   );
   gpc1_1 gpc1085 (
      {stage0_18[159]},
      {stage1_18[60]}
   );
   gpc1_1 gpc1086 (
      {stage0_18[160]},
      {stage1_18[61]}
   );
   gpc1_1 gpc1087 (
      {stage0_18[161]},
      {stage1_18[62]}
   );
   gpc1_1 gpc1088 (
      {stage0_19[156]},
      {stage1_19[65]}
   );
   gpc1_1 gpc1089 (
      {stage0_19[157]},
      {stage1_19[66]}
   );
   gpc1_1 gpc1090 (
      {stage0_19[158]},
      {stage1_19[67]}
   );
   gpc1_1 gpc1091 (
      {stage0_19[159]},
      {stage1_19[68]}
   );
   gpc1_1 gpc1092 (
      {stage0_19[160]},
      {stage1_19[69]}
   );
   gpc1_1 gpc1093 (
      {stage0_19[161]},
      {stage1_19[70]}
   );
   gpc1_1 gpc1094 (
      {stage0_20[159]},
      {stage1_20[65]}
   );
   gpc1_1 gpc1095 (
      {stage0_20[160]},
      {stage1_20[66]}
   );
   gpc1_1 gpc1096 (
      {stage0_20[161]},
      {stage1_20[67]}
   );
   gpc1_1 gpc1097 (
      {stage0_21[147]},
      {stage1_21[56]}
   );
   gpc1_1 gpc1098 (
      {stage0_21[148]},
      {stage1_21[57]}
   );
   gpc1_1 gpc1099 (
      {stage0_21[149]},
      {stage1_21[58]}
   );
   gpc1_1 gpc1100 (
      {stage0_21[150]},
      {stage1_21[59]}
   );
   gpc1_1 gpc1101 (
      {stage0_21[151]},
      {stage1_21[60]}
   );
   gpc1_1 gpc1102 (
      {stage0_21[152]},
      {stage1_21[61]}
   );
   gpc1_1 gpc1103 (
      {stage0_21[153]},
      {stage1_21[62]}
   );
   gpc1_1 gpc1104 (
      {stage0_21[154]},
      {stage1_21[63]}
   );
   gpc1_1 gpc1105 (
      {stage0_21[155]},
      {stage1_21[64]}
   );
   gpc1_1 gpc1106 (
      {stage0_21[156]},
      {stage1_21[65]}
   );
   gpc1_1 gpc1107 (
      {stage0_21[157]},
      {stage1_21[66]}
   );
   gpc1_1 gpc1108 (
      {stage0_21[158]},
      {stage1_21[67]}
   );
   gpc1_1 gpc1109 (
      {stage0_21[159]},
      {stage1_21[68]}
   );
   gpc1_1 gpc1110 (
      {stage0_21[160]},
      {stage1_21[69]}
   );
   gpc1_1 gpc1111 (
      {stage0_21[161]},
      {stage1_21[70]}
   );
   gpc1_1 gpc1112 (
      {stage0_23[77]},
      {stage1_23[58]}
   );
   gpc1_1 gpc1113 (
      {stage0_23[78]},
      {stage1_23[59]}
   );
   gpc1_1 gpc1114 (
      {stage0_23[79]},
      {stage1_23[60]}
   );
   gpc1_1 gpc1115 (
      {stage0_23[80]},
      {stage1_23[61]}
   );
   gpc1_1 gpc1116 (
      {stage0_23[81]},
      {stage1_23[62]}
   );
   gpc1_1 gpc1117 (
      {stage0_23[82]},
      {stage1_23[63]}
   );
   gpc1_1 gpc1118 (
      {stage0_23[83]},
      {stage1_23[64]}
   );
   gpc1_1 gpc1119 (
      {stage0_23[84]},
      {stage1_23[65]}
   );
   gpc1_1 gpc1120 (
      {stage0_23[85]},
      {stage1_23[66]}
   );
   gpc1_1 gpc1121 (
      {stage0_23[86]},
      {stage1_23[67]}
   );
   gpc1_1 gpc1122 (
      {stage0_23[87]},
      {stage1_23[68]}
   );
   gpc1_1 gpc1123 (
      {stage0_23[88]},
      {stage1_23[69]}
   );
   gpc1_1 gpc1124 (
      {stage0_23[89]},
      {stage1_23[70]}
   );
   gpc1_1 gpc1125 (
      {stage0_23[90]},
      {stage1_23[71]}
   );
   gpc1_1 gpc1126 (
      {stage0_23[91]},
      {stage1_23[72]}
   );
   gpc1_1 gpc1127 (
      {stage0_23[92]},
      {stage1_23[73]}
   );
   gpc1_1 gpc1128 (
      {stage0_23[93]},
      {stage1_23[74]}
   );
   gpc1_1 gpc1129 (
      {stage0_23[94]},
      {stage1_23[75]}
   );
   gpc1_1 gpc1130 (
      {stage0_23[95]},
      {stage1_23[76]}
   );
   gpc1_1 gpc1131 (
      {stage0_23[96]},
      {stage1_23[77]}
   );
   gpc1_1 gpc1132 (
      {stage0_23[97]},
      {stage1_23[78]}
   );
   gpc1_1 gpc1133 (
      {stage0_23[98]},
      {stage1_23[79]}
   );
   gpc1_1 gpc1134 (
      {stage0_23[99]},
      {stage1_23[80]}
   );
   gpc1_1 gpc1135 (
      {stage0_23[100]},
      {stage1_23[81]}
   );
   gpc1_1 gpc1136 (
      {stage0_23[101]},
      {stage1_23[82]}
   );
   gpc1_1 gpc1137 (
      {stage0_23[102]},
      {stage1_23[83]}
   );
   gpc1_1 gpc1138 (
      {stage0_23[103]},
      {stage1_23[84]}
   );
   gpc1_1 gpc1139 (
      {stage0_23[104]},
      {stage1_23[85]}
   );
   gpc1_1 gpc1140 (
      {stage0_23[105]},
      {stage1_23[86]}
   );
   gpc1_1 gpc1141 (
      {stage0_23[106]},
      {stage1_23[87]}
   );
   gpc1_1 gpc1142 (
      {stage0_23[107]},
      {stage1_23[88]}
   );
   gpc1_1 gpc1143 (
      {stage0_23[108]},
      {stage1_23[89]}
   );
   gpc1_1 gpc1144 (
      {stage0_23[109]},
      {stage1_23[90]}
   );
   gpc1_1 gpc1145 (
      {stage0_23[110]},
      {stage1_23[91]}
   );
   gpc1_1 gpc1146 (
      {stage0_23[111]},
      {stage1_23[92]}
   );
   gpc1_1 gpc1147 (
      {stage0_23[112]},
      {stage1_23[93]}
   );
   gpc1_1 gpc1148 (
      {stage0_23[113]},
      {stage1_23[94]}
   );
   gpc1_1 gpc1149 (
      {stage0_23[114]},
      {stage1_23[95]}
   );
   gpc1_1 gpc1150 (
      {stage0_23[115]},
      {stage1_23[96]}
   );
   gpc1_1 gpc1151 (
      {stage0_23[116]},
      {stage1_23[97]}
   );
   gpc1_1 gpc1152 (
      {stage0_23[117]},
      {stage1_23[98]}
   );
   gpc1_1 gpc1153 (
      {stage0_23[118]},
      {stage1_23[99]}
   );
   gpc1_1 gpc1154 (
      {stage0_23[119]},
      {stage1_23[100]}
   );
   gpc1_1 gpc1155 (
      {stage0_23[120]},
      {stage1_23[101]}
   );
   gpc1_1 gpc1156 (
      {stage0_23[121]},
      {stage1_23[102]}
   );
   gpc1_1 gpc1157 (
      {stage0_23[122]},
      {stage1_23[103]}
   );
   gpc1_1 gpc1158 (
      {stage0_23[123]},
      {stage1_23[104]}
   );
   gpc1_1 gpc1159 (
      {stage0_23[124]},
      {stage1_23[105]}
   );
   gpc1_1 gpc1160 (
      {stage0_23[125]},
      {stage1_23[106]}
   );
   gpc1_1 gpc1161 (
      {stage0_23[126]},
      {stage1_23[107]}
   );
   gpc1_1 gpc1162 (
      {stage0_23[127]},
      {stage1_23[108]}
   );
   gpc1_1 gpc1163 (
      {stage0_23[128]},
      {stage1_23[109]}
   );
   gpc1_1 gpc1164 (
      {stage0_23[129]},
      {stage1_23[110]}
   );
   gpc1_1 gpc1165 (
      {stage0_23[130]},
      {stage1_23[111]}
   );
   gpc1_1 gpc1166 (
      {stage0_23[131]},
      {stage1_23[112]}
   );
   gpc1_1 gpc1167 (
      {stage0_23[132]},
      {stage1_23[113]}
   );
   gpc1_1 gpc1168 (
      {stage0_23[133]},
      {stage1_23[114]}
   );
   gpc1_1 gpc1169 (
      {stage0_23[134]},
      {stage1_23[115]}
   );
   gpc1_1 gpc1170 (
      {stage0_23[135]},
      {stage1_23[116]}
   );
   gpc1_1 gpc1171 (
      {stage0_23[136]},
      {stage1_23[117]}
   );
   gpc1_1 gpc1172 (
      {stage0_23[137]},
      {stage1_23[118]}
   );
   gpc1_1 gpc1173 (
      {stage0_23[138]},
      {stage1_23[119]}
   );
   gpc1_1 gpc1174 (
      {stage0_23[139]},
      {stage1_23[120]}
   );
   gpc1_1 gpc1175 (
      {stage0_23[140]},
      {stage1_23[121]}
   );
   gpc1_1 gpc1176 (
      {stage0_23[141]},
      {stage1_23[122]}
   );
   gpc1_1 gpc1177 (
      {stage0_23[142]},
      {stage1_23[123]}
   );
   gpc1_1 gpc1178 (
      {stage0_23[143]},
      {stage1_23[124]}
   );
   gpc1_1 gpc1179 (
      {stage0_23[144]},
      {stage1_23[125]}
   );
   gpc1_1 gpc1180 (
      {stage0_23[145]},
      {stage1_23[126]}
   );
   gpc1_1 gpc1181 (
      {stage0_23[146]},
      {stage1_23[127]}
   );
   gpc1_1 gpc1182 (
      {stage0_23[147]},
      {stage1_23[128]}
   );
   gpc1_1 gpc1183 (
      {stage0_23[148]},
      {stage1_23[129]}
   );
   gpc1_1 gpc1184 (
      {stage0_23[149]},
      {stage1_23[130]}
   );
   gpc1_1 gpc1185 (
      {stage0_23[150]},
      {stage1_23[131]}
   );
   gpc1_1 gpc1186 (
      {stage0_23[151]},
      {stage1_23[132]}
   );
   gpc1_1 gpc1187 (
      {stage0_23[152]},
      {stage1_23[133]}
   );
   gpc1_1 gpc1188 (
      {stage0_23[153]},
      {stage1_23[134]}
   );
   gpc1_1 gpc1189 (
      {stage0_23[154]},
      {stage1_23[135]}
   );
   gpc1_1 gpc1190 (
      {stage0_23[155]},
      {stage1_23[136]}
   );
   gpc1_1 gpc1191 (
      {stage0_23[156]},
      {stage1_23[137]}
   );
   gpc1_1 gpc1192 (
      {stage0_23[157]},
      {stage1_23[138]}
   );
   gpc1_1 gpc1193 (
      {stage0_23[158]},
      {stage1_23[139]}
   );
   gpc1_1 gpc1194 (
      {stage0_23[159]},
      {stage1_23[140]}
   );
   gpc1_1 gpc1195 (
      {stage0_23[160]},
      {stage1_23[141]}
   );
   gpc1_1 gpc1196 (
      {stage0_23[161]},
      {stage1_23[142]}
   );
   gpc1_1 gpc1197 (
      {stage0_24[126]},
      {stage1_24[47]}
   );
   gpc1_1 gpc1198 (
      {stage0_24[127]},
      {stage1_24[48]}
   );
   gpc1_1 gpc1199 (
      {stage0_24[128]},
      {stage1_24[49]}
   );
   gpc1_1 gpc1200 (
      {stage0_24[129]},
      {stage1_24[50]}
   );
   gpc1_1 gpc1201 (
      {stage0_24[130]},
      {stage1_24[51]}
   );
   gpc1_1 gpc1202 (
      {stage0_24[131]},
      {stage1_24[52]}
   );
   gpc1_1 gpc1203 (
      {stage0_24[132]},
      {stage1_24[53]}
   );
   gpc1_1 gpc1204 (
      {stage0_24[133]},
      {stage1_24[54]}
   );
   gpc1_1 gpc1205 (
      {stage0_24[134]},
      {stage1_24[55]}
   );
   gpc1_1 gpc1206 (
      {stage0_24[135]},
      {stage1_24[56]}
   );
   gpc1_1 gpc1207 (
      {stage0_24[136]},
      {stage1_24[57]}
   );
   gpc1_1 gpc1208 (
      {stage0_24[137]},
      {stage1_24[58]}
   );
   gpc1_1 gpc1209 (
      {stage0_24[138]},
      {stage1_24[59]}
   );
   gpc1_1 gpc1210 (
      {stage0_24[139]},
      {stage1_24[60]}
   );
   gpc1_1 gpc1211 (
      {stage0_24[140]},
      {stage1_24[61]}
   );
   gpc1_1 gpc1212 (
      {stage0_24[141]},
      {stage1_24[62]}
   );
   gpc1_1 gpc1213 (
      {stage0_24[142]},
      {stage1_24[63]}
   );
   gpc1_1 gpc1214 (
      {stage0_24[143]},
      {stage1_24[64]}
   );
   gpc1_1 gpc1215 (
      {stage0_24[144]},
      {stage1_24[65]}
   );
   gpc1_1 gpc1216 (
      {stage0_24[145]},
      {stage1_24[66]}
   );
   gpc1_1 gpc1217 (
      {stage0_24[146]},
      {stage1_24[67]}
   );
   gpc1_1 gpc1218 (
      {stage0_24[147]},
      {stage1_24[68]}
   );
   gpc1_1 gpc1219 (
      {stage0_24[148]},
      {stage1_24[69]}
   );
   gpc1_1 gpc1220 (
      {stage0_24[149]},
      {stage1_24[70]}
   );
   gpc1_1 gpc1221 (
      {stage0_24[150]},
      {stage1_24[71]}
   );
   gpc1_1 gpc1222 (
      {stage0_24[151]},
      {stage1_24[72]}
   );
   gpc1_1 gpc1223 (
      {stage0_24[152]},
      {stage1_24[73]}
   );
   gpc1_1 gpc1224 (
      {stage0_24[153]},
      {stage1_24[74]}
   );
   gpc1_1 gpc1225 (
      {stage0_24[154]},
      {stage1_24[75]}
   );
   gpc1_1 gpc1226 (
      {stage0_24[155]},
      {stage1_24[76]}
   );
   gpc1_1 gpc1227 (
      {stage0_24[156]},
      {stage1_24[77]}
   );
   gpc1_1 gpc1228 (
      {stage0_24[157]},
      {stage1_24[78]}
   );
   gpc1_1 gpc1229 (
      {stage0_24[158]},
      {stage1_24[79]}
   );
   gpc1_1 gpc1230 (
      {stage0_24[159]},
      {stage1_24[80]}
   );
   gpc1_1 gpc1231 (
      {stage0_24[160]},
      {stage1_24[81]}
   );
   gpc1_1 gpc1232 (
      {stage0_24[161]},
      {stage1_24[82]}
   );
   gpc1_1 gpc1233 (
      {stage0_25[127]},
      {stage1_25[50]}
   );
   gpc1_1 gpc1234 (
      {stage0_25[128]},
      {stage1_25[51]}
   );
   gpc1_1 gpc1235 (
      {stage0_25[129]},
      {stage1_25[52]}
   );
   gpc1_1 gpc1236 (
      {stage0_25[130]},
      {stage1_25[53]}
   );
   gpc1_1 gpc1237 (
      {stage0_25[131]},
      {stage1_25[54]}
   );
   gpc1_1 gpc1238 (
      {stage0_25[132]},
      {stage1_25[55]}
   );
   gpc1_1 gpc1239 (
      {stage0_25[133]},
      {stage1_25[56]}
   );
   gpc1_1 gpc1240 (
      {stage0_25[134]},
      {stage1_25[57]}
   );
   gpc1_1 gpc1241 (
      {stage0_25[135]},
      {stage1_25[58]}
   );
   gpc1_1 gpc1242 (
      {stage0_25[136]},
      {stage1_25[59]}
   );
   gpc1_1 gpc1243 (
      {stage0_25[137]},
      {stage1_25[60]}
   );
   gpc1_1 gpc1244 (
      {stage0_25[138]},
      {stage1_25[61]}
   );
   gpc1_1 gpc1245 (
      {stage0_25[139]},
      {stage1_25[62]}
   );
   gpc1_1 gpc1246 (
      {stage0_25[140]},
      {stage1_25[63]}
   );
   gpc1_1 gpc1247 (
      {stage0_25[141]},
      {stage1_25[64]}
   );
   gpc1_1 gpc1248 (
      {stage0_25[142]},
      {stage1_25[65]}
   );
   gpc1_1 gpc1249 (
      {stage0_25[143]},
      {stage1_25[66]}
   );
   gpc1_1 gpc1250 (
      {stage0_25[144]},
      {stage1_25[67]}
   );
   gpc1_1 gpc1251 (
      {stage0_25[145]},
      {stage1_25[68]}
   );
   gpc1_1 gpc1252 (
      {stage0_25[146]},
      {stage1_25[69]}
   );
   gpc1_1 gpc1253 (
      {stage0_25[147]},
      {stage1_25[70]}
   );
   gpc1_1 gpc1254 (
      {stage0_25[148]},
      {stage1_25[71]}
   );
   gpc1_1 gpc1255 (
      {stage0_25[149]},
      {stage1_25[72]}
   );
   gpc1_1 gpc1256 (
      {stage0_25[150]},
      {stage1_25[73]}
   );
   gpc1_1 gpc1257 (
      {stage0_25[151]},
      {stage1_25[74]}
   );
   gpc1_1 gpc1258 (
      {stage0_25[152]},
      {stage1_25[75]}
   );
   gpc1_1 gpc1259 (
      {stage0_25[153]},
      {stage1_25[76]}
   );
   gpc1_1 gpc1260 (
      {stage0_25[154]},
      {stage1_25[77]}
   );
   gpc1_1 gpc1261 (
      {stage0_25[155]},
      {stage1_25[78]}
   );
   gpc1_1 gpc1262 (
      {stage0_25[156]},
      {stage1_25[79]}
   );
   gpc1_1 gpc1263 (
      {stage0_25[157]},
      {stage1_25[80]}
   );
   gpc1_1 gpc1264 (
      {stage0_25[158]},
      {stage1_25[81]}
   );
   gpc1_1 gpc1265 (
      {stage0_25[159]},
      {stage1_25[82]}
   );
   gpc1_1 gpc1266 (
      {stage0_25[160]},
      {stage1_25[83]}
   );
   gpc1_1 gpc1267 (
      {stage0_25[161]},
      {stage1_25[84]}
   );
   gpc1_1 gpc1268 (
      {stage0_26[149]},
      {stage1_26[59]}
   );
   gpc1_1 gpc1269 (
      {stage0_26[150]},
      {stage1_26[60]}
   );
   gpc1_1 gpc1270 (
      {stage0_26[151]},
      {stage1_26[61]}
   );
   gpc1_1 gpc1271 (
      {stage0_26[152]},
      {stage1_26[62]}
   );
   gpc1_1 gpc1272 (
      {stage0_26[153]},
      {stage1_26[63]}
   );
   gpc1_1 gpc1273 (
      {stage0_26[154]},
      {stage1_26[64]}
   );
   gpc1_1 gpc1274 (
      {stage0_26[155]},
      {stage1_26[65]}
   );
   gpc1_1 gpc1275 (
      {stage0_26[156]},
      {stage1_26[66]}
   );
   gpc1_1 gpc1276 (
      {stage0_26[157]},
      {stage1_26[67]}
   );
   gpc1_1 gpc1277 (
      {stage0_26[158]},
      {stage1_26[68]}
   );
   gpc1_1 gpc1278 (
      {stage0_26[159]},
      {stage1_26[69]}
   );
   gpc1_1 gpc1279 (
      {stage0_26[160]},
      {stage1_26[70]}
   );
   gpc1_1 gpc1280 (
      {stage0_26[161]},
      {stage1_26[71]}
   );
   gpc1_1 gpc1281 (
      {stage0_27[142]},
      {stage1_27[54]}
   );
   gpc1_1 gpc1282 (
      {stage0_27[143]},
      {stage1_27[55]}
   );
   gpc1_1 gpc1283 (
      {stage0_27[144]},
      {stage1_27[56]}
   );
   gpc1_1 gpc1284 (
      {stage0_27[145]},
      {stage1_27[57]}
   );
   gpc1_1 gpc1285 (
      {stage0_27[146]},
      {stage1_27[58]}
   );
   gpc1_1 gpc1286 (
      {stage0_27[147]},
      {stage1_27[59]}
   );
   gpc1_1 gpc1287 (
      {stage0_27[148]},
      {stage1_27[60]}
   );
   gpc1_1 gpc1288 (
      {stage0_27[149]},
      {stage1_27[61]}
   );
   gpc1_1 gpc1289 (
      {stage0_27[150]},
      {stage1_27[62]}
   );
   gpc1_1 gpc1290 (
      {stage0_27[151]},
      {stage1_27[63]}
   );
   gpc1_1 gpc1291 (
      {stage0_27[152]},
      {stage1_27[64]}
   );
   gpc1_1 gpc1292 (
      {stage0_27[153]},
      {stage1_27[65]}
   );
   gpc1_1 gpc1293 (
      {stage0_27[154]},
      {stage1_27[66]}
   );
   gpc1_1 gpc1294 (
      {stage0_27[155]},
      {stage1_27[67]}
   );
   gpc1_1 gpc1295 (
      {stage0_27[156]},
      {stage1_27[68]}
   );
   gpc1_1 gpc1296 (
      {stage0_27[157]},
      {stage1_27[69]}
   );
   gpc1_1 gpc1297 (
      {stage0_27[158]},
      {stage1_27[70]}
   );
   gpc1_1 gpc1298 (
      {stage0_27[159]},
      {stage1_27[71]}
   );
   gpc1_1 gpc1299 (
      {stage0_27[160]},
      {stage1_27[72]}
   );
   gpc1_1 gpc1300 (
      {stage0_27[161]},
      {stage1_27[73]}
   );
   gpc1_1 gpc1301 (
      {stage0_28[140]},
      {stage1_28[55]}
   );
   gpc1_1 gpc1302 (
      {stage0_28[141]},
      {stage1_28[56]}
   );
   gpc1_1 gpc1303 (
      {stage0_28[142]},
      {stage1_28[57]}
   );
   gpc1_1 gpc1304 (
      {stage0_28[143]},
      {stage1_28[58]}
   );
   gpc1_1 gpc1305 (
      {stage0_28[144]},
      {stage1_28[59]}
   );
   gpc1_1 gpc1306 (
      {stage0_28[145]},
      {stage1_28[60]}
   );
   gpc1_1 gpc1307 (
      {stage0_28[146]},
      {stage1_28[61]}
   );
   gpc1_1 gpc1308 (
      {stage0_28[147]},
      {stage1_28[62]}
   );
   gpc1_1 gpc1309 (
      {stage0_28[148]},
      {stage1_28[63]}
   );
   gpc1_1 gpc1310 (
      {stage0_28[149]},
      {stage1_28[64]}
   );
   gpc1_1 gpc1311 (
      {stage0_28[150]},
      {stage1_28[65]}
   );
   gpc1_1 gpc1312 (
      {stage0_28[151]},
      {stage1_28[66]}
   );
   gpc1_1 gpc1313 (
      {stage0_28[152]},
      {stage1_28[67]}
   );
   gpc1_1 gpc1314 (
      {stage0_28[153]},
      {stage1_28[68]}
   );
   gpc1_1 gpc1315 (
      {stage0_28[154]},
      {stage1_28[69]}
   );
   gpc1_1 gpc1316 (
      {stage0_28[155]},
      {stage1_28[70]}
   );
   gpc1_1 gpc1317 (
      {stage0_28[156]},
      {stage1_28[71]}
   );
   gpc1_1 gpc1318 (
      {stage0_28[157]},
      {stage1_28[72]}
   );
   gpc1_1 gpc1319 (
      {stage0_28[158]},
      {stage1_28[73]}
   );
   gpc1_1 gpc1320 (
      {stage0_28[159]},
      {stage1_28[74]}
   );
   gpc1_1 gpc1321 (
      {stage0_28[160]},
      {stage1_28[75]}
   );
   gpc1_1 gpc1322 (
      {stage0_28[161]},
      {stage1_28[76]}
   );
   gpc1_1 gpc1323 (
      {stage0_29[144]},
      {stage1_29[63]}
   );
   gpc1_1 gpc1324 (
      {stage0_29[145]},
      {stage1_29[64]}
   );
   gpc1_1 gpc1325 (
      {stage0_29[146]},
      {stage1_29[65]}
   );
   gpc1_1 gpc1326 (
      {stage0_29[147]},
      {stage1_29[66]}
   );
   gpc1_1 gpc1327 (
      {stage0_29[148]},
      {stage1_29[67]}
   );
   gpc1_1 gpc1328 (
      {stage0_29[149]},
      {stage1_29[68]}
   );
   gpc1_1 gpc1329 (
      {stage0_29[150]},
      {stage1_29[69]}
   );
   gpc1_1 gpc1330 (
      {stage0_29[151]},
      {stage1_29[70]}
   );
   gpc1_1 gpc1331 (
      {stage0_29[152]},
      {stage1_29[71]}
   );
   gpc1_1 gpc1332 (
      {stage0_29[153]},
      {stage1_29[72]}
   );
   gpc1_1 gpc1333 (
      {stage0_29[154]},
      {stage1_29[73]}
   );
   gpc1_1 gpc1334 (
      {stage0_29[155]},
      {stage1_29[74]}
   );
   gpc1_1 gpc1335 (
      {stage0_29[156]},
      {stage1_29[75]}
   );
   gpc1_1 gpc1336 (
      {stage0_29[157]},
      {stage1_29[76]}
   );
   gpc1_1 gpc1337 (
      {stage0_29[158]},
      {stage1_29[77]}
   );
   gpc1_1 gpc1338 (
      {stage0_29[159]},
      {stage1_29[78]}
   );
   gpc1_1 gpc1339 (
      {stage0_29[160]},
      {stage1_29[79]}
   );
   gpc1_1 gpc1340 (
      {stage0_29[161]},
      {stage1_29[80]}
   );
   gpc1_1 gpc1341 (
      {stage0_30[111]},
      {stage1_30[56]}
   );
   gpc1_1 gpc1342 (
      {stage0_30[112]},
      {stage1_30[57]}
   );
   gpc1_1 gpc1343 (
      {stage0_30[113]},
      {stage1_30[58]}
   );
   gpc1_1 gpc1344 (
      {stage0_30[114]},
      {stage1_30[59]}
   );
   gpc1_1 gpc1345 (
      {stage0_30[115]},
      {stage1_30[60]}
   );
   gpc1_1 gpc1346 (
      {stage0_30[116]},
      {stage1_30[61]}
   );
   gpc1_1 gpc1347 (
      {stage0_30[117]},
      {stage1_30[62]}
   );
   gpc1_1 gpc1348 (
      {stage0_30[118]},
      {stage1_30[63]}
   );
   gpc1_1 gpc1349 (
      {stage0_30[119]},
      {stage1_30[64]}
   );
   gpc1_1 gpc1350 (
      {stage0_30[120]},
      {stage1_30[65]}
   );
   gpc1_1 gpc1351 (
      {stage0_30[121]},
      {stage1_30[66]}
   );
   gpc1_1 gpc1352 (
      {stage0_30[122]},
      {stage1_30[67]}
   );
   gpc1_1 gpc1353 (
      {stage0_30[123]},
      {stage1_30[68]}
   );
   gpc1_1 gpc1354 (
      {stage0_30[124]},
      {stage1_30[69]}
   );
   gpc1_1 gpc1355 (
      {stage0_30[125]},
      {stage1_30[70]}
   );
   gpc1_1 gpc1356 (
      {stage0_30[126]},
      {stage1_30[71]}
   );
   gpc1_1 gpc1357 (
      {stage0_30[127]},
      {stage1_30[72]}
   );
   gpc1_1 gpc1358 (
      {stage0_30[128]},
      {stage1_30[73]}
   );
   gpc1_1 gpc1359 (
      {stage0_30[129]},
      {stage1_30[74]}
   );
   gpc1_1 gpc1360 (
      {stage0_30[130]},
      {stage1_30[75]}
   );
   gpc1_1 gpc1361 (
      {stage0_30[131]},
      {stage1_30[76]}
   );
   gpc1_1 gpc1362 (
      {stage0_30[132]},
      {stage1_30[77]}
   );
   gpc1_1 gpc1363 (
      {stage0_30[133]},
      {stage1_30[78]}
   );
   gpc1_1 gpc1364 (
      {stage0_30[134]},
      {stage1_30[79]}
   );
   gpc1_1 gpc1365 (
      {stage0_30[135]},
      {stage1_30[80]}
   );
   gpc1_1 gpc1366 (
      {stage0_30[136]},
      {stage1_30[81]}
   );
   gpc1_1 gpc1367 (
      {stage0_30[137]},
      {stage1_30[82]}
   );
   gpc1_1 gpc1368 (
      {stage0_30[138]},
      {stage1_30[83]}
   );
   gpc1_1 gpc1369 (
      {stage0_30[139]},
      {stage1_30[84]}
   );
   gpc1_1 gpc1370 (
      {stage0_30[140]},
      {stage1_30[85]}
   );
   gpc1_1 gpc1371 (
      {stage0_30[141]},
      {stage1_30[86]}
   );
   gpc1_1 gpc1372 (
      {stage0_30[142]},
      {stage1_30[87]}
   );
   gpc1_1 gpc1373 (
      {stage0_30[143]},
      {stage1_30[88]}
   );
   gpc1_1 gpc1374 (
      {stage0_30[144]},
      {stage1_30[89]}
   );
   gpc1_1 gpc1375 (
      {stage0_30[145]},
      {stage1_30[90]}
   );
   gpc1_1 gpc1376 (
      {stage0_30[146]},
      {stage1_30[91]}
   );
   gpc1_1 gpc1377 (
      {stage0_30[147]},
      {stage1_30[92]}
   );
   gpc1_1 gpc1378 (
      {stage0_30[148]},
      {stage1_30[93]}
   );
   gpc1_1 gpc1379 (
      {stage0_30[149]},
      {stage1_30[94]}
   );
   gpc1_1 gpc1380 (
      {stage0_30[150]},
      {stage1_30[95]}
   );
   gpc1_1 gpc1381 (
      {stage0_30[151]},
      {stage1_30[96]}
   );
   gpc1_1 gpc1382 (
      {stage0_30[152]},
      {stage1_30[97]}
   );
   gpc1_1 gpc1383 (
      {stage0_30[153]},
      {stage1_30[98]}
   );
   gpc1_1 gpc1384 (
      {stage0_30[154]},
      {stage1_30[99]}
   );
   gpc1_1 gpc1385 (
      {stage0_30[155]},
      {stage1_30[100]}
   );
   gpc1_1 gpc1386 (
      {stage0_30[156]},
      {stage1_30[101]}
   );
   gpc1_1 gpc1387 (
      {stage0_30[157]},
      {stage1_30[102]}
   );
   gpc1_1 gpc1388 (
      {stage0_30[158]},
      {stage1_30[103]}
   );
   gpc1_1 gpc1389 (
      {stage0_30[159]},
      {stage1_30[104]}
   );
   gpc1_1 gpc1390 (
      {stage0_30[160]},
      {stage1_30[105]}
   );
   gpc1_1 gpc1391 (
      {stage0_30[161]},
      {stage1_30[106]}
   );
   gpc1_1 gpc1392 (
      {stage0_31[109]},
      {stage1_31[44]}
   );
   gpc1_1 gpc1393 (
      {stage0_31[110]},
      {stage1_31[45]}
   );
   gpc1_1 gpc1394 (
      {stage0_31[111]},
      {stage1_31[46]}
   );
   gpc1_1 gpc1395 (
      {stage0_31[112]},
      {stage1_31[47]}
   );
   gpc1_1 gpc1396 (
      {stage0_31[113]},
      {stage1_31[48]}
   );
   gpc1_1 gpc1397 (
      {stage0_31[114]},
      {stage1_31[49]}
   );
   gpc1_1 gpc1398 (
      {stage0_31[115]},
      {stage1_31[50]}
   );
   gpc1_1 gpc1399 (
      {stage0_31[116]},
      {stage1_31[51]}
   );
   gpc1_1 gpc1400 (
      {stage0_31[117]},
      {stage1_31[52]}
   );
   gpc1_1 gpc1401 (
      {stage0_31[118]},
      {stage1_31[53]}
   );
   gpc1_1 gpc1402 (
      {stage0_31[119]},
      {stage1_31[54]}
   );
   gpc1_1 gpc1403 (
      {stage0_31[120]},
      {stage1_31[55]}
   );
   gpc1_1 gpc1404 (
      {stage0_31[121]},
      {stage1_31[56]}
   );
   gpc1_1 gpc1405 (
      {stage0_31[122]},
      {stage1_31[57]}
   );
   gpc1_1 gpc1406 (
      {stage0_31[123]},
      {stage1_31[58]}
   );
   gpc1_1 gpc1407 (
      {stage0_31[124]},
      {stage1_31[59]}
   );
   gpc1_1 gpc1408 (
      {stage0_31[125]},
      {stage1_31[60]}
   );
   gpc1_1 gpc1409 (
      {stage0_31[126]},
      {stage1_31[61]}
   );
   gpc1_1 gpc1410 (
      {stage0_31[127]},
      {stage1_31[62]}
   );
   gpc1_1 gpc1411 (
      {stage0_31[128]},
      {stage1_31[63]}
   );
   gpc1_1 gpc1412 (
      {stage0_31[129]},
      {stage1_31[64]}
   );
   gpc1_1 gpc1413 (
      {stage0_31[130]},
      {stage1_31[65]}
   );
   gpc1_1 gpc1414 (
      {stage0_31[131]},
      {stage1_31[66]}
   );
   gpc1_1 gpc1415 (
      {stage0_31[132]},
      {stage1_31[67]}
   );
   gpc1_1 gpc1416 (
      {stage0_31[133]},
      {stage1_31[68]}
   );
   gpc1_1 gpc1417 (
      {stage0_31[134]},
      {stage1_31[69]}
   );
   gpc1_1 gpc1418 (
      {stage0_31[135]},
      {stage1_31[70]}
   );
   gpc1_1 gpc1419 (
      {stage0_31[136]},
      {stage1_31[71]}
   );
   gpc1_1 gpc1420 (
      {stage0_31[137]},
      {stage1_31[72]}
   );
   gpc1_1 gpc1421 (
      {stage0_31[138]},
      {stage1_31[73]}
   );
   gpc1_1 gpc1422 (
      {stage0_31[139]},
      {stage1_31[74]}
   );
   gpc1_1 gpc1423 (
      {stage0_31[140]},
      {stage1_31[75]}
   );
   gpc1_1 gpc1424 (
      {stage0_31[141]},
      {stage1_31[76]}
   );
   gpc1_1 gpc1425 (
      {stage0_31[142]},
      {stage1_31[77]}
   );
   gpc1_1 gpc1426 (
      {stage0_31[143]},
      {stage1_31[78]}
   );
   gpc1_1 gpc1427 (
      {stage0_31[144]},
      {stage1_31[79]}
   );
   gpc1_1 gpc1428 (
      {stage0_31[145]},
      {stage1_31[80]}
   );
   gpc1_1 gpc1429 (
      {stage0_31[146]},
      {stage1_31[81]}
   );
   gpc1_1 gpc1430 (
      {stage0_31[147]},
      {stage1_31[82]}
   );
   gpc1_1 gpc1431 (
      {stage0_31[148]},
      {stage1_31[83]}
   );
   gpc1_1 gpc1432 (
      {stage0_31[149]},
      {stage1_31[84]}
   );
   gpc1_1 gpc1433 (
      {stage0_31[150]},
      {stage1_31[85]}
   );
   gpc1_1 gpc1434 (
      {stage0_31[151]},
      {stage1_31[86]}
   );
   gpc1_1 gpc1435 (
      {stage0_31[152]},
      {stage1_31[87]}
   );
   gpc1_1 gpc1436 (
      {stage0_31[153]},
      {stage1_31[88]}
   );
   gpc1_1 gpc1437 (
      {stage0_31[154]},
      {stage1_31[89]}
   );
   gpc1_1 gpc1438 (
      {stage0_31[155]},
      {stage1_31[90]}
   );
   gpc1_1 gpc1439 (
      {stage0_31[156]},
      {stage1_31[91]}
   );
   gpc1_1 gpc1440 (
      {stage0_31[157]},
      {stage1_31[92]}
   );
   gpc1_1 gpc1441 (
      {stage0_31[158]},
      {stage1_31[93]}
   );
   gpc1_1 gpc1442 (
      {stage0_31[159]},
      {stage1_31[94]}
   );
   gpc1_1 gpc1443 (
      {stage0_31[160]},
      {stage1_31[95]}
   );
   gpc1_1 gpc1444 (
      {stage0_31[161]},
      {stage1_31[96]}
   );
   gpc1_1 gpc1445 (
      {stage0_32[129]},
      {stage1_32[54]}
   );
   gpc1_1 gpc1446 (
      {stage0_32[130]},
      {stage1_32[55]}
   );
   gpc1_1 gpc1447 (
      {stage0_32[131]},
      {stage1_32[56]}
   );
   gpc1_1 gpc1448 (
      {stage0_32[132]},
      {stage1_32[57]}
   );
   gpc1_1 gpc1449 (
      {stage0_32[133]},
      {stage1_32[58]}
   );
   gpc1_1 gpc1450 (
      {stage0_32[134]},
      {stage1_32[59]}
   );
   gpc1_1 gpc1451 (
      {stage0_32[135]},
      {stage1_32[60]}
   );
   gpc1_1 gpc1452 (
      {stage0_32[136]},
      {stage1_32[61]}
   );
   gpc1_1 gpc1453 (
      {stage0_32[137]},
      {stage1_32[62]}
   );
   gpc1_1 gpc1454 (
      {stage0_32[138]},
      {stage1_32[63]}
   );
   gpc1_1 gpc1455 (
      {stage0_32[139]},
      {stage1_32[64]}
   );
   gpc1_1 gpc1456 (
      {stage0_32[140]},
      {stage1_32[65]}
   );
   gpc1_1 gpc1457 (
      {stage0_32[141]},
      {stage1_32[66]}
   );
   gpc1_1 gpc1458 (
      {stage0_32[142]},
      {stage1_32[67]}
   );
   gpc1_1 gpc1459 (
      {stage0_32[143]},
      {stage1_32[68]}
   );
   gpc1_1 gpc1460 (
      {stage0_32[144]},
      {stage1_32[69]}
   );
   gpc1_1 gpc1461 (
      {stage0_32[145]},
      {stage1_32[70]}
   );
   gpc1_1 gpc1462 (
      {stage0_32[146]},
      {stage1_32[71]}
   );
   gpc1_1 gpc1463 (
      {stage0_32[147]},
      {stage1_32[72]}
   );
   gpc1_1 gpc1464 (
      {stage0_32[148]},
      {stage1_32[73]}
   );
   gpc1_1 gpc1465 (
      {stage0_32[149]},
      {stage1_32[74]}
   );
   gpc1_1 gpc1466 (
      {stage0_32[150]},
      {stage1_32[75]}
   );
   gpc1_1 gpc1467 (
      {stage0_32[151]},
      {stage1_32[76]}
   );
   gpc1_1 gpc1468 (
      {stage0_32[152]},
      {stage1_32[77]}
   );
   gpc1_1 gpc1469 (
      {stage0_32[153]},
      {stage1_32[78]}
   );
   gpc1_1 gpc1470 (
      {stage0_32[154]},
      {stage1_32[79]}
   );
   gpc1_1 gpc1471 (
      {stage0_32[155]},
      {stage1_32[80]}
   );
   gpc1_1 gpc1472 (
      {stage0_32[156]},
      {stage1_32[81]}
   );
   gpc1_1 gpc1473 (
      {stage0_32[157]},
      {stage1_32[82]}
   );
   gpc1_1 gpc1474 (
      {stage0_32[158]},
      {stage1_32[83]}
   );
   gpc1_1 gpc1475 (
      {stage0_32[159]},
      {stage1_32[84]}
   );
   gpc1_1 gpc1476 (
      {stage0_32[160]},
      {stage1_32[85]}
   );
   gpc1_1 gpc1477 (
      {stage0_32[161]},
      {stage1_32[86]}
   );
   gpc1_1 gpc1478 (
      {stage0_33[136]},
      {stage1_33[64]}
   );
   gpc1_1 gpc1479 (
      {stage0_33[137]},
      {stage1_33[65]}
   );
   gpc1_1 gpc1480 (
      {stage0_33[138]},
      {stage1_33[66]}
   );
   gpc1_1 gpc1481 (
      {stage0_33[139]},
      {stage1_33[67]}
   );
   gpc1_1 gpc1482 (
      {stage0_33[140]},
      {stage1_33[68]}
   );
   gpc1_1 gpc1483 (
      {stage0_33[141]},
      {stage1_33[69]}
   );
   gpc1_1 gpc1484 (
      {stage0_33[142]},
      {stage1_33[70]}
   );
   gpc1_1 gpc1485 (
      {stage0_33[143]},
      {stage1_33[71]}
   );
   gpc1_1 gpc1486 (
      {stage0_33[144]},
      {stage1_33[72]}
   );
   gpc1_1 gpc1487 (
      {stage0_33[145]},
      {stage1_33[73]}
   );
   gpc1_1 gpc1488 (
      {stage0_33[146]},
      {stage1_33[74]}
   );
   gpc1_1 gpc1489 (
      {stage0_33[147]},
      {stage1_33[75]}
   );
   gpc1_1 gpc1490 (
      {stage0_33[148]},
      {stage1_33[76]}
   );
   gpc1_1 gpc1491 (
      {stage0_33[149]},
      {stage1_33[77]}
   );
   gpc1_1 gpc1492 (
      {stage0_33[150]},
      {stage1_33[78]}
   );
   gpc1_1 gpc1493 (
      {stage0_33[151]},
      {stage1_33[79]}
   );
   gpc1_1 gpc1494 (
      {stage0_33[152]},
      {stage1_33[80]}
   );
   gpc1_1 gpc1495 (
      {stage0_33[153]},
      {stage1_33[81]}
   );
   gpc1_1 gpc1496 (
      {stage0_33[154]},
      {stage1_33[82]}
   );
   gpc1_1 gpc1497 (
      {stage0_33[155]},
      {stage1_33[83]}
   );
   gpc1_1 gpc1498 (
      {stage0_33[156]},
      {stage1_33[84]}
   );
   gpc1_1 gpc1499 (
      {stage0_33[157]},
      {stage1_33[85]}
   );
   gpc1_1 gpc1500 (
      {stage0_33[158]},
      {stage1_33[86]}
   );
   gpc1_1 gpc1501 (
      {stage0_33[159]},
      {stage1_33[87]}
   );
   gpc1_1 gpc1502 (
      {stage0_33[160]},
      {stage1_33[88]}
   );
   gpc1_1 gpc1503 (
      {stage0_33[161]},
      {stage1_33[89]}
   );
   gpc1_1 gpc1504 (
      {stage0_34[158]},
      {stage1_34[52]}
   );
   gpc1_1 gpc1505 (
      {stage0_34[159]},
      {stage1_34[53]}
   );
   gpc1_1 gpc1506 (
      {stage0_34[160]},
      {stage1_34[54]}
   );
   gpc1_1 gpc1507 (
      {stage0_34[161]},
      {stage1_34[55]}
   );
   gpc1_1 gpc1508 (
      {stage0_35[158]},
      {stage1_35[56]}
   );
   gpc1_1 gpc1509 (
      {stage0_35[159]},
      {stage1_35[57]}
   );
   gpc1_1 gpc1510 (
      {stage0_35[160]},
      {stage1_35[58]}
   );
   gpc1_1 gpc1511 (
      {stage0_35[161]},
      {stage1_35[59]}
   );
   gpc1_1 gpc1512 (
      {stage0_36[146]},
      {stage1_36[67]}
   );
   gpc1_1 gpc1513 (
      {stage0_36[147]},
      {stage1_36[68]}
   );
   gpc1_1 gpc1514 (
      {stage0_36[148]},
      {stage1_36[69]}
   );
   gpc1_1 gpc1515 (
      {stage0_36[149]},
      {stage1_36[70]}
   );
   gpc1_1 gpc1516 (
      {stage0_36[150]},
      {stage1_36[71]}
   );
   gpc1_1 gpc1517 (
      {stage0_36[151]},
      {stage1_36[72]}
   );
   gpc1_1 gpc1518 (
      {stage0_36[152]},
      {stage1_36[73]}
   );
   gpc1_1 gpc1519 (
      {stage0_36[153]},
      {stage1_36[74]}
   );
   gpc1_1 gpc1520 (
      {stage0_36[154]},
      {stage1_36[75]}
   );
   gpc1_1 gpc1521 (
      {stage0_36[155]},
      {stage1_36[76]}
   );
   gpc1_1 gpc1522 (
      {stage0_36[156]},
      {stage1_36[77]}
   );
   gpc1_1 gpc1523 (
      {stage0_36[157]},
      {stage1_36[78]}
   );
   gpc1_1 gpc1524 (
      {stage0_36[158]},
      {stage1_36[79]}
   );
   gpc1_1 gpc1525 (
      {stage0_36[159]},
      {stage1_36[80]}
   );
   gpc1_1 gpc1526 (
      {stage0_36[160]},
      {stage1_36[81]}
   );
   gpc1_1 gpc1527 (
      {stage0_36[161]},
      {stage1_36[82]}
   );
   gpc1_1 gpc1528 (
      {stage0_37[90]},
      {stage1_37[56]}
   );
   gpc1_1 gpc1529 (
      {stage0_37[91]},
      {stage1_37[57]}
   );
   gpc1_1 gpc1530 (
      {stage0_37[92]},
      {stage1_37[58]}
   );
   gpc1_1 gpc1531 (
      {stage0_37[93]},
      {stage1_37[59]}
   );
   gpc1_1 gpc1532 (
      {stage0_37[94]},
      {stage1_37[60]}
   );
   gpc1_1 gpc1533 (
      {stage0_37[95]},
      {stage1_37[61]}
   );
   gpc1_1 gpc1534 (
      {stage0_37[96]},
      {stage1_37[62]}
   );
   gpc1_1 gpc1535 (
      {stage0_37[97]},
      {stage1_37[63]}
   );
   gpc1_1 gpc1536 (
      {stage0_37[98]},
      {stage1_37[64]}
   );
   gpc1_1 gpc1537 (
      {stage0_37[99]},
      {stage1_37[65]}
   );
   gpc1_1 gpc1538 (
      {stage0_37[100]},
      {stage1_37[66]}
   );
   gpc1_1 gpc1539 (
      {stage0_37[101]},
      {stage1_37[67]}
   );
   gpc1_1 gpc1540 (
      {stage0_37[102]},
      {stage1_37[68]}
   );
   gpc1_1 gpc1541 (
      {stage0_37[103]},
      {stage1_37[69]}
   );
   gpc1_1 gpc1542 (
      {stage0_37[104]},
      {stage1_37[70]}
   );
   gpc1_1 gpc1543 (
      {stage0_37[105]},
      {stage1_37[71]}
   );
   gpc1_1 gpc1544 (
      {stage0_37[106]},
      {stage1_37[72]}
   );
   gpc1_1 gpc1545 (
      {stage0_37[107]},
      {stage1_37[73]}
   );
   gpc1_1 gpc1546 (
      {stage0_37[108]},
      {stage1_37[74]}
   );
   gpc1_1 gpc1547 (
      {stage0_37[109]},
      {stage1_37[75]}
   );
   gpc1_1 gpc1548 (
      {stage0_37[110]},
      {stage1_37[76]}
   );
   gpc1_1 gpc1549 (
      {stage0_37[111]},
      {stage1_37[77]}
   );
   gpc1_1 gpc1550 (
      {stage0_37[112]},
      {stage1_37[78]}
   );
   gpc1_1 gpc1551 (
      {stage0_37[113]},
      {stage1_37[79]}
   );
   gpc1_1 gpc1552 (
      {stage0_37[114]},
      {stage1_37[80]}
   );
   gpc1_1 gpc1553 (
      {stage0_37[115]},
      {stage1_37[81]}
   );
   gpc1_1 gpc1554 (
      {stage0_37[116]},
      {stage1_37[82]}
   );
   gpc1_1 gpc1555 (
      {stage0_37[117]},
      {stage1_37[83]}
   );
   gpc1_1 gpc1556 (
      {stage0_37[118]},
      {stage1_37[84]}
   );
   gpc1_1 gpc1557 (
      {stage0_37[119]},
      {stage1_37[85]}
   );
   gpc1_1 gpc1558 (
      {stage0_37[120]},
      {stage1_37[86]}
   );
   gpc1_1 gpc1559 (
      {stage0_37[121]},
      {stage1_37[87]}
   );
   gpc1_1 gpc1560 (
      {stage0_37[122]},
      {stage1_37[88]}
   );
   gpc1_1 gpc1561 (
      {stage0_37[123]},
      {stage1_37[89]}
   );
   gpc1_1 gpc1562 (
      {stage0_37[124]},
      {stage1_37[90]}
   );
   gpc1_1 gpc1563 (
      {stage0_37[125]},
      {stage1_37[91]}
   );
   gpc1_1 gpc1564 (
      {stage0_37[126]},
      {stage1_37[92]}
   );
   gpc1_1 gpc1565 (
      {stage0_37[127]},
      {stage1_37[93]}
   );
   gpc1_1 gpc1566 (
      {stage0_37[128]},
      {stage1_37[94]}
   );
   gpc1_1 gpc1567 (
      {stage0_37[129]},
      {stage1_37[95]}
   );
   gpc1_1 gpc1568 (
      {stage0_37[130]},
      {stage1_37[96]}
   );
   gpc1_1 gpc1569 (
      {stage0_37[131]},
      {stage1_37[97]}
   );
   gpc1_1 gpc1570 (
      {stage0_37[132]},
      {stage1_37[98]}
   );
   gpc1_1 gpc1571 (
      {stage0_37[133]},
      {stage1_37[99]}
   );
   gpc1_1 gpc1572 (
      {stage0_37[134]},
      {stage1_37[100]}
   );
   gpc1_1 gpc1573 (
      {stage0_37[135]},
      {stage1_37[101]}
   );
   gpc1_1 gpc1574 (
      {stage0_37[136]},
      {stage1_37[102]}
   );
   gpc1_1 gpc1575 (
      {stage0_37[137]},
      {stage1_37[103]}
   );
   gpc1_1 gpc1576 (
      {stage0_37[138]},
      {stage1_37[104]}
   );
   gpc1_1 gpc1577 (
      {stage0_37[139]},
      {stage1_37[105]}
   );
   gpc1_1 gpc1578 (
      {stage0_37[140]},
      {stage1_37[106]}
   );
   gpc1_1 gpc1579 (
      {stage0_37[141]},
      {stage1_37[107]}
   );
   gpc1_1 gpc1580 (
      {stage0_37[142]},
      {stage1_37[108]}
   );
   gpc1_1 gpc1581 (
      {stage0_37[143]},
      {stage1_37[109]}
   );
   gpc1_1 gpc1582 (
      {stage0_37[144]},
      {stage1_37[110]}
   );
   gpc1_1 gpc1583 (
      {stage0_37[145]},
      {stage1_37[111]}
   );
   gpc1_1 gpc1584 (
      {stage0_37[146]},
      {stage1_37[112]}
   );
   gpc1_1 gpc1585 (
      {stage0_37[147]},
      {stage1_37[113]}
   );
   gpc1_1 gpc1586 (
      {stage0_37[148]},
      {stage1_37[114]}
   );
   gpc1_1 gpc1587 (
      {stage0_37[149]},
      {stage1_37[115]}
   );
   gpc1_1 gpc1588 (
      {stage0_37[150]},
      {stage1_37[116]}
   );
   gpc1_1 gpc1589 (
      {stage0_37[151]},
      {stage1_37[117]}
   );
   gpc1_1 gpc1590 (
      {stage0_37[152]},
      {stage1_37[118]}
   );
   gpc1_1 gpc1591 (
      {stage0_37[153]},
      {stage1_37[119]}
   );
   gpc1_1 gpc1592 (
      {stage0_37[154]},
      {stage1_37[120]}
   );
   gpc1_1 gpc1593 (
      {stage0_37[155]},
      {stage1_37[121]}
   );
   gpc1_1 gpc1594 (
      {stage0_37[156]},
      {stage1_37[122]}
   );
   gpc1_1 gpc1595 (
      {stage0_37[157]},
      {stage1_37[123]}
   );
   gpc1_1 gpc1596 (
      {stage0_37[158]},
      {stage1_37[124]}
   );
   gpc1_1 gpc1597 (
      {stage0_37[159]},
      {stage1_37[125]}
   );
   gpc1_1 gpc1598 (
      {stage0_37[160]},
      {stage1_37[126]}
   );
   gpc1_1 gpc1599 (
      {stage0_37[161]},
      {stage1_37[127]}
   );
   gpc1_1 gpc1600 (
      {stage0_38[148]},
      {stage1_38[52]}
   );
   gpc1_1 gpc1601 (
      {stage0_38[149]},
      {stage1_38[53]}
   );
   gpc1_1 gpc1602 (
      {stage0_38[150]},
      {stage1_38[54]}
   );
   gpc1_1 gpc1603 (
      {stage0_38[151]},
      {stage1_38[55]}
   );
   gpc1_1 gpc1604 (
      {stage0_38[152]},
      {stage1_38[56]}
   );
   gpc1_1 gpc1605 (
      {stage0_38[153]},
      {stage1_38[57]}
   );
   gpc1_1 gpc1606 (
      {stage0_38[154]},
      {stage1_38[58]}
   );
   gpc1_1 gpc1607 (
      {stage0_38[155]},
      {stage1_38[59]}
   );
   gpc1_1 gpc1608 (
      {stage0_38[156]},
      {stage1_38[60]}
   );
   gpc1_1 gpc1609 (
      {stage0_38[157]},
      {stage1_38[61]}
   );
   gpc1_1 gpc1610 (
      {stage0_38[158]},
      {stage1_38[62]}
   );
   gpc1_1 gpc1611 (
      {stage0_38[159]},
      {stage1_38[63]}
   );
   gpc1_1 gpc1612 (
      {stage0_38[160]},
      {stage1_38[64]}
   );
   gpc1_1 gpc1613 (
      {stage0_38[161]},
      {stage1_38[65]}
   );
   gpc1_1 gpc1614 (
      {stage0_39[156]},
      {stage1_39[62]}
   );
   gpc1_1 gpc1615 (
      {stage0_39[157]},
      {stage1_39[63]}
   );
   gpc1_1 gpc1616 (
      {stage0_39[158]},
      {stage1_39[64]}
   );
   gpc1_1 gpc1617 (
      {stage0_39[159]},
      {stage1_39[65]}
   );
   gpc1_1 gpc1618 (
      {stage0_39[160]},
      {stage1_39[66]}
   );
   gpc1_1 gpc1619 (
      {stage0_39[161]},
      {stage1_39[67]}
   );
   gpc1_1 gpc1620 (
      {stage0_40[140]},
      {stage1_40[60]}
   );
   gpc1_1 gpc1621 (
      {stage0_40[141]},
      {stage1_40[61]}
   );
   gpc1_1 gpc1622 (
      {stage0_40[142]},
      {stage1_40[62]}
   );
   gpc1_1 gpc1623 (
      {stage0_40[143]},
      {stage1_40[63]}
   );
   gpc1_1 gpc1624 (
      {stage0_40[144]},
      {stage1_40[64]}
   );
   gpc1_1 gpc1625 (
      {stage0_40[145]},
      {stage1_40[65]}
   );
   gpc1_1 gpc1626 (
      {stage0_40[146]},
      {stage1_40[66]}
   );
   gpc1_1 gpc1627 (
      {stage0_40[147]},
      {stage1_40[67]}
   );
   gpc1_1 gpc1628 (
      {stage0_40[148]},
      {stage1_40[68]}
   );
   gpc1_1 gpc1629 (
      {stage0_40[149]},
      {stage1_40[69]}
   );
   gpc1_1 gpc1630 (
      {stage0_40[150]},
      {stage1_40[70]}
   );
   gpc1_1 gpc1631 (
      {stage0_40[151]},
      {stage1_40[71]}
   );
   gpc1_1 gpc1632 (
      {stage0_40[152]},
      {stage1_40[72]}
   );
   gpc1_1 gpc1633 (
      {stage0_40[153]},
      {stage1_40[73]}
   );
   gpc1_1 gpc1634 (
      {stage0_40[154]},
      {stage1_40[74]}
   );
   gpc1_1 gpc1635 (
      {stage0_40[155]},
      {stage1_40[75]}
   );
   gpc1_1 gpc1636 (
      {stage0_40[156]},
      {stage1_40[76]}
   );
   gpc1_1 gpc1637 (
      {stage0_40[157]},
      {stage1_40[77]}
   );
   gpc1_1 gpc1638 (
      {stage0_40[158]},
      {stage1_40[78]}
   );
   gpc1_1 gpc1639 (
      {stage0_40[159]},
      {stage1_40[79]}
   );
   gpc1_1 gpc1640 (
      {stage0_40[160]},
      {stage1_40[80]}
   );
   gpc1_1 gpc1641 (
      {stage0_40[161]},
      {stage1_40[81]}
   );
   gpc1_1 gpc1642 (
      {stage0_41[138]},
      {stage1_41[50]}
   );
   gpc1_1 gpc1643 (
      {stage0_41[139]},
      {stage1_41[51]}
   );
   gpc1_1 gpc1644 (
      {stage0_41[140]},
      {stage1_41[52]}
   );
   gpc1_1 gpc1645 (
      {stage0_41[141]},
      {stage1_41[53]}
   );
   gpc1_1 gpc1646 (
      {stage0_41[142]},
      {stage1_41[54]}
   );
   gpc1_1 gpc1647 (
      {stage0_41[143]},
      {stage1_41[55]}
   );
   gpc1_1 gpc1648 (
      {stage0_41[144]},
      {stage1_41[56]}
   );
   gpc1_1 gpc1649 (
      {stage0_41[145]},
      {stage1_41[57]}
   );
   gpc1_1 gpc1650 (
      {stage0_41[146]},
      {stage1_41[58]}
   );
   gpc1_1 gpc1651 (
      {stage0_41[147]},
      {stage1_41[59]}
   );
   gpc1_1 gpc1652 (
      {stage0_41[148]},
      {stage1_41[60]}
   );
   gpc1_1 gpc1653 (
      {stage0_41[149]},
      {stage1_41[61]}
   );
   gpc1_1 gpc1654 (
      {stage0_41[150]},
      {stage1_41[62]}
   );
   gpc1_1 gpc1655 (
      {stage0_41[151]},
      {stage1_41[63]}
   );
   gpc1_1 gpc1656 (
      {stage0_41[152]},
      {stage1_41[64]}
   );
   gpc1_1 gpc1657 (
      {stage0_41[153]},
      {stage1_41[65]}
   );
   gpc1_1 gpc1658 (
      {stage0_41[154]},
      {stage1_41[66]}
   );
   gpc1_1 gpc1659 (
      {stage0_41[155]},
      {stage1_41[67]}
   );
   gpc1_1 gpc1660 (
      {stage0_41[156]},
      {stage1_41[68]}
   );
   gpc1_1 gpc1661 (
      {stage0_41[157]},
      {stage1_41[69]}
   );
   gpc1_1 gpc1662 (
      {stage0_41[158]},
      {stage1_41[70]}
   );
   gpc1_1 gpc1663 (
      {stage0_41[159]},
      {stage1_41[71]}
   );
   gpc1_1 gpc1664 (
      {stage0_41[160]},
      {stage1_41[72]}
   );
   gpc1_1 gpc1665 (
      {stage0_41[161]},
      {stage1_41[73]}
   );
   gpc1_1 gpc1666 (
      {stage0_42[126]},
      {stage1_42[60]}
   );
   gpc1_1 gpc1667 (
      {stage0_42[127]},
      {stage1_42[61]}
   );
   gpc1_1 gpc1668 (
      {stage0_42[128]},
      {stage1_42[62]}
   );
   gpc1_1 gpc1669 (
      {stage0_42[129]},
      {stage1_42[63]}
   );
   gpc1_1 gpc1670 (
      {stage0_42[130]},
      {stage1_42[64]}
   );
   gpc1_1 gpc1671 (
      {stage0_42[131]},
      {stage1_42[65]}
   );
   gpc1_1 gpc1672 (
      {stage0_42[132]},
      {stage1_42[66]}
   );
   gpc1_1 gpc1673 (
      {stage0_42[133]},
      {stage1_42[67]}
   );
   gpc1_1 gpc1674 (
      {stage0_42[134]},
      {stage1_42[68]}
   );
   gpc1_1 gpc1675 (
      {stage0_42[135]},
      {stage1_42[69]}
   );
   gpc1_1 gpc1676 (
      {stage0_42[136]},
      {stage1_42[70]}
   );
   gpc1_1 gpc1677 (
      {stage0_42[137]},
      {stage1_42[71]}
   );
   gpc1_1 gpc1678 (
      {stage0_42[138]},
      {stage1_42[72]}
   );
   gpc1_1 gpc1679 (
      {stage0_42[139]},
      {stage1_42[73]}
   );
   gpc1_1 gpc1680 (
      {stage0_42[140]},
      {stage1_42[74]}
   );
   gpc1_1 gpc1681 (
      {stage0_42[141]},
      {stage1_42[75]}
   );
   gpc1_1 gpc1682 (
      {stage0_42[142]},
      {stage1_42[76]}
   );
   gpc1_1 gpc1683 (
      {stage0_42[143]},
      {stage1_42[77]}
   );
   gpc1_1 gpc1684 (
      {stage0_42[144]},
      {stage1_42[78]}
   );
   gpc1_1 gpc1685 (
      {stage0_42[145]},
      {stage1_42[79]}
   );
   gpc1_1 gpc1686 (
      {stage0_42[146]},
      {stage1_42[80]}
   );
   gpc1_1 gpc1687 (
      {stage0_42[147]},
      {stage1_42[81]}
   );
   gpc1_1 gpc1688 (
      {stage0_42[148]},
      {stage1_42[82]}
   );
   gpc1_1 gpc1689 (
      {stage0_42[149]},
      {stage1_42[83]}
   );
   gpc1_1 gpc1690 (
      {stage0_42[150]},
      {stage1_42[84]}
   );
   gpc1_1 gpc1691 (
      {stage0_42[151]},
      {stage1_42[85]}
   );
   gpc1_1 gpc1692 (
      {stage0_42[152]},
      {stage1_42[86]}
   );
   gpc1_1 gpc1693 (
      {stage0_42[153]},
      {stage1_42[87]}
   );
   gpc1_1 gpc1694 (
      {stage0_42[154]},
      {stage1_42[88]}
   );
   gpc1_1 gpc1695 (
      {stage0_42[155]},
      {stage1_42[89]}
   );
   gpc1_1 gpc1696 (
      {stage0_42[156]},
      {stage1_42[90]}
   );
   gpc1_1 gpc1697 (
      {stage0_42[157]},
      {stage1_42[91]}
   );
   gpc1_1 gpc1698 (
      {stage0_42[158]},
      {stage1_42[92]}
   );
   gpc1_1 gpc1699 (
      {stage0_42[159]},
      {stage1_42[93]}
   );
   gpc1_1 gpc1700 (
      {stage0_42[160]},
      {stage1_42[94]}
   );
   gpc1_1 gpc1701 (
      {stage0_42[161]},
      {stage1_42[95]}
   );
   gpc1_1 gpc1702 (
      {stage0_43[78]},
      {stage1_43[54]}
   );
   gpc1_1 gpc1703 (
      {stage0_43[79]},
      {stage1_43[55]}
   );
   gpc1_1 gpc1704 (
      {stage0_43[80]},
      {stage1_43[56]}
   );
   gpc1_1 gpc1705 (
      {stage0_43[81]},
      {stage1_43[57]}
   );
   gpc1_1 gpc1706 (
      {stage0_43[82]},
      {stage1_43[58]}
   );
   gpc1_1 gpc1707 (
      {stage0_43[83]},
      {stage1_43[59]}
   );
   gpc1_1 gpc1708 (
      {stage0_43[84]},
      {stage1_43[60]}
   );
   gpc1_1 gpc1709 (
      {stage0_43[85]},
      {stage1_43[61]}
   );
   gpc1_1 gpc1710 (
      {stage0_43[86]},
      {stage1_43[62]}
   );
   gpc1_1 gpc1711 (
      {stage0_43[87]},
      {stage1_43[63]}
   );
   gpc1_1 gpc1712 (
      {stage0_43[88]},
      {stage1_43[64]}
   );
   gpc1_1 gpc1713 (
      {stage0_43[89]},
      {stage1_43[65]}
   );
   gpc1_1 gpc1714 (
      {stage0_43[90]},
      {stage1_43[66]}
   );
   gpc1_1 gpc1715 (
      {stage0_43[91]},
      {stage1_43[67]}
   );
   gpc1_1 gpc1716 (
      {stage0_43[92]},
      {stage1_43[68]}
   );
   gpc1_1 gpc1717 (
      {stage0_43[93]},
      {stage1_43[69]}
   );
   gpc1_1 gpc1718 (
      {stage0_43[94]},
      {stage1_43[70]}
   );
   gpc1_1 gpc1719 (
      {stage0_43[95]},
      {stage1_43[71]}
   );
   gpc1_1 gpc1720 (
      {stage0_43[96]},
      {stage1_43[72]}
   );
   gpc1_1 gpc1721 (
      {stage0_43[97]},
      {stage1_43[73]}
   );
   gpc1_1 gpc1722 (
      {stage0_43[98]},
      {stage1_43[74]}
   );
   gpc1_1 gpc1723 (
      {stage0_43[99]},
      {stage1_43[75]}
   );
   gpc1_1 gpc1724 (
      {stage0_43[100]},
      {stage1_43[76]}
   );
   gpc1_1 gpc1725 (
      {stage0_43[101]},
      {stage1_43[77]}
   );
   gpc1_1 gpc1726 (
      {stage0_43[102]},
      {stage1_43[78]}
   );
   gpc1_1 gpc1727 (
      {stage0_43[103]},
      {stage1_43[79]}
   );
   gpc1_1 gpc1728 (
      {stage0_43[104]},
      {stage1_43[80]}
   );
   gpc1_1 gpc1729 (
      {stage0_43[105]},
      {stage1_43[81]}
   );
   gpc1_1 gpc1730 (
      {stage0_43[106]},
      {stage1_43[82]}
   );
   gpc1_1 gpc1731 (
      {stage0_43[107]},
      {stage1_43[83]}
   );
   gpc1_1 gpc1732 (
      {stage0_43[108]},
      {stage1_43[84]}
   );
   gpc1_1 gpc1733 (
      {stage0_43[109]},
      {stage1_43[85]}
   );
   gpc1_1 gpc1734 (
      {stage0_43[110]},
      {stage1_43[86]}
   );
   gpc1_1 gpc1735 (
      {stage0_43[111]},
      {stage1_43[87]}
   );
   gpc1_1 gpc1736 (
      {stage0_43[112]},
      {stage1_43[88]}
   );
   gpc1_1 gpc1737 (
      {stage0_43[113]},
      {stage1_43[89]}
   );
   gpc1_1 gpc1738 (
      {stage0_43[114]},
      {stage1_43[90]}
   );
   gpc1_1 gpc1739 (
      {stage0_43[115]},
      {stage1_43[91]}
   );
   gpc1_1 gpc1740 (
      {stage0_43[116]},
      {stage1_43[92]}
   );
   gpc1_1 gpc1741 (
      {stage0_43[117]},
      {stage1_43[93]}
   );
   gpc1_1 gpc1742 (
      {stage0_43[118]},
      {stage1_43[94]}
   );
   gpc1_1 gpc1743 (
      {stage0_43[119]},
      {stage1_43[95]}
   );
   gpc1_1 gpc1744 (
      {stage0_43[120]},
      {stage1_43[96]}
   );
   gpc1_1 gpc1745 (
      {stage0_43[121]},
      {stage1_43[97]}
   );
   gpc1_1 gpc1746 (
      {stage0_43[122]},
      {stage1_43[98]}
   );
   gpc1_1 gpc1747 (
      {stage0_43[123]},
      {stage1_43[99]}
   );
   gpc1_1 gpc1748 (
      {stage0_43[124]},
      {stage1_43[100]}
   );
   gpc1_1 gpc1749 (
      {stage0_43[125]},
      {stage1_43[101]}
   );
   gpc1_1 gpc1750 (
      {stage0_43[126]},
      {stage1_43[102]}
   );
   gpc1_1 gpc1751 (
      {stage0_43[127]},
      {stage1_43[103]}
   );
   gpc1_1 gpc1752 (
      {stage0_43[128]},
      {stage1_43[104]}
   );
   gpc1_1 gpc1753 (
      {stage0_43[129]},
      {stage1_43[105]}
   );
   gpc1_1 gpc1754 (
      {stage0_43[130]},
      {stage1_43[106]}
   );
   gpc1_1 gpc1755 (
      {stage0_43[131]},
      {stage1_43[107]}
   );
   gpc1_1 gpc1756 (
      {stage0_43[132]},
      {stage1_43[108]}
   );
   gpc1_1 gpc1757 (
      {stage0_43[133]},
      {stage1_43[109]}
   );
   gpc1_1 gpc1758 (
      {stage0_43[134]},
      {stage1_43[110]}
   );
   gpc1_1 gpc1759 (
      {stage0_43[135]},
      {stage1_43[111]}
   );
   gpc1_1 gpc1760 (
      {stage0_43[136]},
      {stage1_43[112]}
   );
   gpc1_1 gpc1761 (
      {stage0_43[137]},
      {stage1_43[113]}
   );
   gpc1_1 gpc1762 (
      {stage0_43[138]},
      {stage1_43[114]}
   );
   gpc1_1 gpc1763 (
      {stage0_43[139]},
      {stage1_43[115]}
   );
   gpc1_1 gpc1764 (
      {stage0_43[140]},
      {stage1_43[116]}
   );
   gpc1_1 gpc1765 (
      {stage0_43[141]},
      {stage1_43[117]}
   );
   gpc1_1 gpc1766 (
      {stage0_43[142]},
      {stage1_43[118]}
   );
   gpc1_1 gpc1767 (
      {stage0_43[143]},
      {stage1_43[119]}
   );
   gpc1_1 gpc1768 (
      {stage0_43[144]},
      {stage1_43[120]}
   );
   gpc1_1 gpc1769 (
      {stage0_43[145]},
      {stage1_43[121]}
   );
   gpc1_1 gpc1770 (
      {stage0_43[146]},
      {stage1_43[122]}
   );
   gpc1_1 gpc1771 (
      {stage0_43[147]},
      {stage1_43[123]}
   );
   gpc1_1 gpc1772 (
      {stage0_43[148]},
      {stage1_43[124]}
   );
   gpc1_1 gpc1773 (
      {stage0_43[149]},
      {stage1_43[125]}
   );
   gpc1_1 gpc1774 (
      {stage0_43[150]},
      {stage1_43[126]}
   );
   gpc1_1 gpc1775 (
      {stage0_43[151]},
      {stage1_43[127]}
   );
   gpc1_1 gpc1776 (
      {stage0_43[152]},
      {stage1_43[128]}
   );
   gpc1_1 gpc1777 (
      {stage0_43[153]},
      {stage1_43[129]}
   );
   gpc1_1 gpc1778 (
      {stage0_43[154]},
      {stage1_43[130]}
   );
   gpc1_1 gpc1779 (
      {stage0_43[155]},
      {stage1_43[131]}
   );
   gpc1_1 gpc1780 (
      {stage0_43[156]},
      {stage1_43[132]}
   );
   gpc1_1 gpc1781 (
      {stage0_43[157]},
      {stage1_43[133]}
   );
   gpc1_1 gpc1782 (
      {stage0_43[158]},
      {stage1_43[134]}
   );
   gpc1_1 gpc1783 (
      {stage0_43[159]},
      {stage1_43[135]}
   );
   gpc1_1 gpc1784 (
      {stage0_43[160]},
      {stage1_43[136]}
   );
   gpc1_1 gpc1785 (
      {stage0_43[161]},
      {stage1_43[137]}
   );
   gpc1_1 gpc1786 (
      {stage0_44[160]},
      {stage1_44[44]}
   );
   gpc1_1 gpc1787 (
      {stage0_44[161]},
      {stage1_44[45]}
   );
   gpc1_1 gpc1788 (
      {stage0_45[121]},
      {stage1_45[52]}
   );
   gpc1_1 gpc1789 (
      {stage0_45[122]},
      {stage1_45[53]}
   );
   gpc1_1 gpc1790 (
      {stage0_45[123]},
      {stage1_45[54]}
   );
   gpc1_1 gpc1791 (
      {stage0_45[124]},
      {stage1_45[55]}
   );
   gpc1_1 gpc1792 (
      {stage0_45[125]},
      {stage1_45[56]}
   );
   gpc1_1 gpc1793 (
      {stage0_45[126]},
      {stage1_45[57]}
   );
   gpc1_1 gpc1794 (
      {stage0_45[127]},
      {stage1_45[58]}
   );
   gpc1_1 gpc1795 (
      {stage0_45[128]},
      {stage1_45[59]}
   );
   gpc1_1 gpc1796 (
      {stage0_45[129]},
      {stage1_45[60]}
   );
   gpc1_1 gpc1797 (
      {stage0_45[130]},
      {stage1_45[61]}
   );
   gpc1_1 gpc1798 (
      {stage0_45[131]},
      {stage1_45[62]}
   );
   gpc1_1 gpc1799 (
      {stage0_45[132]},
      {stage1_45[63]}
   );
   gpc1_1 gpc1800 (
      {stage0_45[133]},
      {stage1_45[64]}
   );
   gpc1_1 gpc1801 (
      {stage0_45[134]},
      {stage1_45[65]}
   );
   gpc1_1 gpc1802 (
      {stage0_45[135]},
      {stage1_45[66]}
   );
   gpc1_1 gpc1803 (
      {stage0_45[136]},
      {stage1_45[67]}
   );
   gpc1_1 gpc1804 (
      {stage0_45[137]},
      {stage1_45[68]}
   );
   gpc1_1 gpc1805 (
      {stage0_45[138]},
      {stage1_45[69]}
   );
   gpc1_1 gpc1806 (
      {stage0_45[139]},
      {stage1_45[70]}
   );
   gpc1_1 gpc1807 (
      {stage0_45[140]},
      {stage1_45[71]}
   );
   gpc1_1 gpc1808 (
      {stage0_45[141]},
      {stage1_45[72]}
   );
   gpc1_1 gpc1809 (
      {stage0_45[142]},
      {stage1_45[73]}
   );
   gpc1_1 gpc1810 (
      {stage0_45[143]},
      {stage1_45[74]}
   );
   gpc1_1 gpc1811 (
      {stage0_45[144]},
      {stage1_45[75]}
   );
   gpc1_1 gpc1812 (
      {stage0_45[145]},
      {stage1_45[76]}
   );
   gpc1_1 gpc1813 (
      {stage0_45[146]},
      {stage1_45[77]}
   );
   gpc1_1 gpc1814 (
      {stage0_45[147]},
      {stage1_45[78]}
   );
   gpc1_1 gpc1815 (
      {stage0_45[148]},
      {stage1_45[79]}
   );
   gpc1_1 gpc1816 (
      {stage0_45[149]},
      {stage1_45[80]}
   );
   gpc1_1 gpc1817 (
      {stage0_45[150]},
      {stage1_45[81]}
   );
   gpc1_1 gpc1818 (
      {stage0_45[151]},
      {stage1_45[82]}
   );
   gpc1_1 gpc1819 (
      {stage0_45[152]},
      {stage1_45[83]}
   );
   gpc1_1 gpc1820 (
      {stage0_45[153]},
      {stage1_45[84]}
   );
   gpc1_1 gpc1821 (
      {stage0_45[154]},
      {stage1_45[85]}
   );
   gpc1_1 gpc1822 (
      {stage0_45[155]},
      {stage1_45[86]}
   );
   gpc1_1 gpc1823 (
      {stage0_45[156]},
      {stage1_45[87]}
   );
   gpc1_1 gpc1824 (
      {stage0_45[157]},
      {stage1_45[88]}
   );
   gpc1_1 gpc1825 (
      {stage0_45[158]},
      {stage1_45[89]}
   );
   gpc1_1 gpc1826 (
      {stage0_45[159]},
      {stage1_45[90]}
   );
   gpc1_1 gpc1827 (
      {stage0_45[160]},
      {stage1_45[91]}
   );
   gpc1_1 gpc1828 (
      {stage0_45[161]},
      {stage1_45[92]}
   );
   gpc1_1 gpc1829 (
      {stage0_46[161]},
      {stage1_46[63]}
   );
   gpc1_1 gpc1830 (
      {stage0_48[161]},
      {stage1_48[71]}
   );
   gpc1_1 gpc1831 (
      {stage0_49[147]},
      {stage1_49[72]}
   );
   gpc1_1 gpc1832 (
      {stage0_49[148]},
      {stage1_49[73]}
   );
   gpc1_1 gpc1833 (
      {stage0_49[149]},
      {stage1_49[74]}
   );
   gpc1_1 gpc1834 (
      {stage0_49[150]},
      {stage1_49[75]}
   );
   gpc1_1 gpc1835 (
      {stage0_49[151]},
      {stage1_49[76]}
   );
   gpc1_1 gpc1836 (
      {stage0_49[152]},
      {stage1_49[77]}
   );
   gpc1_1 gpc1837 (
      {stage0_49[153]},
      {stage1_49[78]}
   );
   gpc1_1 gpc1838 (
      {stage0_49[154]},
      {stage1_49[79]}
   );
   gpc1_1 gpc1839 (
      {stage0_49[155]},
      {stage1_49[80]}
   );
   gpc1_1 gpc1840 (
      {stage0_49[156]},
      {stage1_49[81]}
   );
   gpc1_1 gpc1841 (
      {stage0_49[157]},
      {stage1_49[82]}
   );
   gpc1_1 gpc1842 (
      {stage0_49[158]},
      {stage1_49[83]}
   );
   gpc1_1 gpc1843 (
      {stage0_49[159]},
      {stage1_49[84]}
   );
   gpc1_1 gpc1844 (
      {stage0_49[160]},
      {stage1_49[85]}
   );
   gpc1_1 gpc1845 (
      {stage0_49[161]},
      {stage1_49[86]}
   );
   gpc1_1 gpc1846 (
      {stage0_50[159]},
      {stage1_50[55]}
   );
   gpc1_1 gpc1847 (
      {stage0_50[160]},
      {stage1_50[56]}
   );
   gpc1_1 gpc1848 (
      {stage0_50[161]},
      {stage1_50[57]}
   );
   gpc1_1 gpc1849 (
      {stage0_51[126]},
      {stage1_51[58]}
   );
   gpc1_1 gpc1850 (
      {stage0_51[127]},
      {stage1_51[59]}
   );
   gpc1_1 gpc1851 (
      {stage0_51[128]},
      {stage1_51[60]}
   );
   gpc1_1 gpc1852 (
      {stage0_51[129]},
      {stage1_51[61]}
   );
   gpc1_1 gpc1853 (
      {stage0_51[130]},
      {stage1_51[62]}
   );
   gpc1_1 gpc1854 (
      {stage0_51[131]},
      {stage1_51[63]}
   );
   gpc1_1 gpc1855 (
      {stage0_51[132]},
      {stage1_51[64]}
   );
   gpc1_1 gpc1856 (
      {stage0_51[133]},
      {stage1_51[65]}
   );
   gpc1_1 gpc1857 (
      {stage0_51[134]},
      {stage1_51[66]}
   );
   gpc1_1 gpc1858 (
      {stage0_51[135]},
      {stage1_51[67]}
   );
   gpc1_1 gpc1859 (
      {stage0_51[136]},
      {stage1_51[68]}
   );
   gpc1_1 gpc1860 (
      {stage0_51[137]},
      {stage1_51[69]}
   );
   gpc1_1 gpc1861 (
      {stage0_51[138]},
      {stage1_51[70]}
   );
   gpc1_1 gpc1862 (
      {stage0_51[139]},
      {stage1_51[71]}
   );
   gpc1_1 gpc1863 (
      {stage0_51[140]},
      {stage1_51[72]}
   );
   gpc1_1 gpc1864 (
      {stage0_51[141]},
      {stage1_51[73]}
   );
   gpc1_1 gpc1865 (
      {stage0_51[142]},
      {stage1_51[74]}
   );
   gpc1_1 gpc1866 (
      {stage0_51[143]},
      {stage1_51[75]}
   );
   gpc1_1 gpc1867 (
      {stage0_51[144]},
      {stage1_51[76]}
   );
   gpc1_1 gpc1868 (
      {stage0_51[145]},
      {stage1_51[77]}
   );
   gpc1_1 gpc1869 (
      {stage0_51[146]},
      {stage1_51[78]}
   );
   gpc1_1 gpc1870 (
      {stage0_51[147]},
      {stage1_51[79]}
   );
   gpc1_1 gpc1871 (
      {stage0_51[148]},
      {stage1_51[80]}
   );
   gpc1_1 gpc1872 (
      {stage0_51[149]},
      {stage1_51[81]}
   );
   gpc1_1 gpc1873 (
      {stage0_51[150]},
      {stage1_51[82]}
   );
   gpc1_1 gpc1874 (
      {stage0_51[151]},
      {stage1_51[83]}
   );
   gpc1_1 gpc1875 (
      {stage0_51[152]},
      {stage1_51[84]}
   );
   gpc1_1 gpc1876 (
      {stage0_51[153]},
      {stage1_51[85]}
   );
   gpc1_1 gpc1877 (
      {stage0_51[154]},
      {stage1_51[86]}
   );
   gpc1_1 gpc1878 (
      {stage0_51[155]},
      {stage1_51[87]}
   );
   gpc1_1 gpc1879 (
      {stage0_51[156]},
      {stage1_51[88]}
   );
   gpc1_1 gpc1880 (
      {stage0_51[157]},
      {stage1_51[89]}
   );
   gpc1_1 gpc1881 (
      {stage0_51[158]},
      {stage1_51[90]}
   );
   gpc1_1 gpc1882 (
      {stage0_51[159]},
      {stage1_51[91]}
   );
   gpc1_1 gpc1883 (
      {stage0_51[160]},
      {stage1_51[92]}
   );
   gpc1_1 gpc1884 (
      {stage0_51[161]},
      {stage1_51[93]}
   );
   gpc1_1 gpc1885 (
      {stage0_52[153]},
      {stage1_52[68]}
   );
   gpc1_1 gpc1886 (
      {stage0_52[154]},
      {stage1_52[69]}
   );
   gpc1_1 gpc1887 (
      {stage0_52[155]},
      {stage1_52[70]}
   );
   gpc1_1 gpc1888 (
      {stage0_52[156]},
      {stage1_52[71]}
   );
   gpc1_1 gpc1889 (
      {stage0_52[157]},
      {stage1_52[72]}
   );
   gpc1_1 gpc1890 (
      {stage0_52[158]},
      {stage1_52[73]}
   );
   gpc1_1 gpc1891 (
      {stage0_52[159]},
      {stage1_52[74]}
   );
   gpc1_1 gpc1892 (
      {stage0_52[160]},
      {stage1_52[75]}
   );
   gpc1_1 gpc1893 (
      {stage0_52[161]},
      {stage1_52[76]}
   );
   gpc1_1 gpc1894 (
      {stage0_53[159]},
      {stage1_53[63]}
   );
   gpc1_1 gpc1895 (
      {stage0_53[160]},
      {stage1_53[64]}
   );
   gpc1_1 gpc1896 (
      {stage0_53[161]},
      {stage1_53[65]}
   );
   gpc1_1 gpc1897 (
      {stage0_55[122]},
      {stage1_55[58]}
   );
   gpc1_1 gpc1898 (
      {stage0_55[123]},
      {stage1_55[59]}
   );
   gpc1_1 gpc1899 (
      {stage0_55[124]},
      {stage1_55[60]}
   );
   gpc1_1 gpc1900 (
      {stage0_55[125]},
      {stage1_55[61]}
   );
   gpc1_1 gpc1901 (
      {stage0_55[126]},
      {stage1_55[62]}
   );
   gpc1_1 gpc1902 (
      {stage0_55[127]},
      {stage1_55[63]}
   );
   gpc1_1 gpc1903 (
      {stage0_55[128]},
      {stage1_55[64]}
   );
   gpc1_1 gpc1904 (
      {stage0_55[129]},
      {stage1_55[65]}
   );
   gpc1_1 gpc1905 (
      {stage0_55[130]},
      {stage1_55[66]}
   );
   gpc1_1 gpc1906 (
      {stage0_55[131]},
      {stage1_55[67]}
   );
   gpc1_1 gpc1907 (
      {stage0_55[132]},
      {stage1_55[68]}
   );
   gpc1_1 gpc1908 (
      {stage0_55[133]},
      {stage1_55[69]}
   );
   gpc1_1 gpc1909 (
      {stage0_55[134]},
      {stage1_55[70]}
   );
   gpc1_1 gpc1910 (
      {stage0_55[135]},
      {stage1_55[71]}
   );
   gpc1_1 gpc1911 (
      {stage0_55[136]},
      {stage1_55[72]}
   );
   gpc1_1 gpc1912 (
      {stage0_55[137]},
      {stage1_55[73]}
   );
   gpc1_1 gpc1913 (
      {stage0_55[138]},
      {stage1_55[74]}
   );
   gpc1_1 gpc1914 (
      {stage0_55[139]},
      {stage1_55[75]}
   );
   gpc1_1 gpc1915 (
      {stage0_55[140]},
      {stage1_55[76]}
   );
   gpc1_1 gpc1916 (
      {stage0_55[141]},
      {stage1_55[77]}
   );
   gpc1_1 gpc1917 (
      {stage0_55[142]},
      {stage1_55[78]}
   );
   gpc1_1 gpc1918 (
      {stage0_55[143]},
      {stage1_55[79]}
   );
   gpc1_1 gpc1919 (
      {stage0_55[144]},
      {stage1_55[80]}
   );
   gpc1_1 gpc1920 (
      {stage0_55[145]},
      {stage1_55[81]}
   );
   gpc1_1 gpc1921 (
      {stage0_55[146]},
      {stage1_55[82]}
   );
   gpc1_1 gpc1922 (
      {stage0_55[147]},
      {stage1_55[83]}
   );
   gpc1_1 gpc1923 (
      {stage0_55[148]},
      {stage1_55[84]}
   );
   gpc1_1 gpc1924 (
      {stage0_55[149]},
      {stage1_55[85]}
   );
   gpc1_1 gpc1925 (
      {stage0_55[150]},
      {stage1_55[86]}
   );
   gpc1_1 gpc1926 (
      {stage0_55[151]},
      {stage1_55[87]}
   );
   gpc1_1 gpc1927 (
      {stage0_55[152]},
      {stage1_55[88]}
   );
   gpc1_1 gpc1928 (
      {stage0_55[153]},
      {stage1_55[89]}
   );
   gpc1_1 gpc1929 (
      {stage0_55[154]},
      {stage1_55[90]}
   );
   gpc1_1 gpc1930 (
      {stage0_55[155]},
      {stage1_55[91]}
   );
   gpc1_1 gpc1931 (
      {stage0_55[156]},
      {stage1_55[92]}
   );
   gpc1_1 gpc1932 (
      {stage0_55[157]},
      {stage1_55[93]}
   );
   gpc1_1 gpc1933 (
      {stage0_55[158]},
      {stage1_55[94]}
   );
   gpc1_1 gpc1934 (
      {stage0_55[159]},
      {stage1_55[95]}
   );
   gpc1_1 gpc1935 (
      {stage0_55[160]},
      {stage1_55[96]}
   );
   gpc1_1 gpc1936 (
      {stage0_55[161]},
      {stage1_55[97]}
   );
   gpc1_1 gpc1937 (
      {stage0_56[148]},
      {stage1_56[66]}
   );
   gpc1_1 gpc1938 (
      {stage0_56[149]},
      {stage1_56[67]}
   );
   gpc1_1 gpc1939 (
      {stage0_56[150]},
      {stage1_56[68]}
   );
   gpc1_1 gpc1940 (
      {stage0_56[151]},
      {stage1_56[69]}
   );
   gpc1_1 gpc1941 (
      {stage0_56[152]},
      {stage1_56[70]}
   );
   gpc1_1 gpc1942 (
      {stage0_56[153]},
      {stage1_56[71]}
   );
   gpc1_1 gpc1943 (
      {stage0_56[154]},
      {stage1_56[72]}
   );
   gpc1_1 gpc1944 (
      {stage0_56[155]},
      {stage1_56[73]}
   );
   gpc1_1 gpc1945 (
      {stage0_56[156]},
      {stage1_56[74]}
   );
   gpc1_1 gpc1946 (
      {stage0_56[157]},
      {stage1_56[75]}
   );
   gpc1_1 gpc1947 (
      {stage0_56[158]},
      {stage1_56[76]}
   );
   gpc1_1 gpc1948 (
      {stage0_56[159]},
      {stage1_56[77]}
   );
   gpc1_1 gpc1949 (
      {stage0_56[160]},
      {stage1_56[78]}
   );
   gpc1_1 gpc1950 (
      {stage0_56[161]},
      {stage1_56[79]}
   );
   gpc1_1 gpc1951 (
      {stage0_57[156]},
      {stage1_57[66]}
   );
   gpc1_1 gpc1952 (
      {stage0_57[157]},
      {stage1_57[67]}
   );
   gpc1_1 gpc1953 (
      {stage0_57[158]},
      {stage1_57[68]}
   );
   gpc1_1 gpc1954 (
      {stage0_57[159]},
      {stage1_57[69]}
   );
   gpc1_1 gpc1955 (
      {stage0_57[160]},
      {stage1_57[70]}
   );
   gpc1_1 gpc1956 (
      {stage0_57[161]},
      {stage1_57[71]}
   );
   gpc1_1 gpc1957 (
      {stage0_58[144]},
      {stage1_58[56]}
   );
   gpc1_1 gpc1958 (
      {stage0_58[145]},
      {stage1_58[57]}
   );
   gpc1_1 gpc1959 (
      {stage0_58[146]},
      {stage1_58[58]}
   );
   gpc1_1 gpc1960 (
      {stage0_58[147]},
      {stage1_58[59]}
   );
   gpc1_1 gpc1961 (
      {stage0_58[148]},
      {stage1_58[60]}
   );
   gpc1_1 gpc1962 (
      {stage0_58[149]},
      {stage1_58[61]}
   );
   gpc1_1 gpc1963 (
      {stage0_58[150]},
      {stage1_58[62]}
   );
   gpc1_1 gpc1964 (
      {stage0_58[151]},
      {stage1_58[63]}
   );
   gpc1_1 gpc1965 (
      {stage0_58[152]},
      {stage1_58[64]}
   );
   gpc1_1 gpc1966 (
      {stage0_58[153]},
      {stage1_58[65]}
   );
   gpc1_1 gpc1967 (
      {stage0_58[154]},
      {stage1_58[66]}
   );
   gpc1_1 gpc1968 (
      {stage0_58[155]},
      {stage1_58[67]}
   );
   gpc1_1 gpc1969 (
      {stage0_58[156]},
      {stage1_58[68]}
   );
   gpc1_1 gpc1970 (
      {stage0_58[157]},
      {stage1_58[69]}
   );
   gpc1_1 gpc1971 (
      {stage0_58[158]},
      {stage1_58[70]}
   );
   gpc1_1 gpc1972 (
      {stage0_58[159]},
      {stage1_58[71]}
   );
   gpc1_1 gpc1973 (
      {stage0_58[160]},
      {stage1_58[72]}
   );
   gpc1_1 gpc1974 (
      {stage0_58[161]},
      {stage1_58[73]}
   );
   gpc1_1 gpc1975 (
      {stage0_59[132]},
      {stage1_59[50]}
   );
   gpc1_1 gpc1976 (
      {stage0_59[133]},
      {stage1_59[51]}
   );
   gpc1_1 gpc1977 (
      {stage0_59[134]},
      {stage1_59[52]}
   );
   gpc1_1 gpc1978 (
      {stage0_59[135]},
      {stage1_59[53]}
   );
   gpc1_1 gpc1979 (
      {stage0_59[136]},
      {stage1_59[54]}
   );
   gpc1_1 gpc1980 (
      {stage0_59[137]},
      {stage1_59[55]}
   );
   gpc1_1 gpc1981 (
      {stage0_59[138]},
      {stage1_59[56]}
   );
   gpc1_1 gpc1982 (
      {stage0_59[139]},
      {stage1_59[57]}
   );
   gpc1_1 gpc1983 (
      {stage0_59[140]},
      {stage1_59[58]}
   );
   gpc1_1 gpc1984 (
      {stage0_59[141]},
      {stage1_59[59]}
   );
   gpc1_1 gpc1985 (
      {stage0_59[142]},
      {stage1_59[60]}
   );
   gpc1_1 gpc1986 (
      {stage0_59[143]},
      {stage1_59[61]}
   );
   gpc1_1 gpc1987 (
      {stage0_59[144]},
      {stage1_59[62]}
   );
   gpc1_1 gpc1988 (
      {stage0_59[145]},
      {stage1_59[63]}
   );
   gpc1_1 gpc1989 (
      {stage0_59[146]},
      {stage1_59[64]}
   );
   gpc1_1 gpc1990 (
      {stage0_59[147]},
      {stage1_59[65]}
   );
   gpc1_1 gpc1991 (
      {stage0_59[148]},
      {stage1_59[66]}
   );
   gpc1_1 gpc1992 (
      {stage0_59[149]},
      {stage1_59[67]}
   );
   gpc1_1 gpc1993 (
      {stage0_59[150]},
      {stage1_59[68]}
   );
   gpc1_1 gpc1994 (
      {stage0_59[151]},
      {stage1_59[69]}
   );
   gpc1_1 gpc1995 (
      {stage0_59[152]},
      {stage1_59[70]}
   );
   gpc1_1 gpc1996 (
      {stage0_59[153]},
      {stage1_59[71]}
   );
   gpc1_1 gpc1997 (
      {stage0_59[154]},
      {stage1_59[72]}
   );
   gpc1_1 gpc1998 (
      {stage0_59[155]},
      {stage1_59[73]}
   );
   gpc1_1 gpc1999 (
      {stage0_59[156]},
      {stage1_59[74]}
   );
   gpc1_1 gpc2000 (
      {stage0_59[157]},
      {stage1_59[75]}
   );
   gpc1_1 gpc2001 (
      {stage0_59[158]},
      {stage1_59[76]}
   );
   gpc1_1 gpc2002 (
      {stage0_59[159]},
      {stage1_59[77]}
   );
   gpc1_1 gpc2003 (
      {stage0_59[160]},
      {stage1_59[78]}
   );
   gpc1_1 gpc2004 (
      {stage0_59[161]},
      {stage1_59[79]}
   );
   gpc1_1 gpc2005 (
      {stage0_61[144]},
      {stage1_61[73]}
   );
   gpc1_1 gpc2006 (
      {stage0_61[145]},
      {stage1_61[74]}
   );
   gpc1_1 gpc2007 (
      {stage0_61[146]},
      {stage1_61[75]}
   );
   gpc1_1 gpc2008 (
      {stage0_61[147]},
      {stage1_61[76]}
   );
   gpc1_1 gpc2009 (
      {stage0_61[148]},
      {stage1_61[77]}
   );
   gpc1_1 gpc2010 (
      {stage0_61[149]},
      {stage1_61[78]}
   );
   gpc1_1 gpc2011 (
      {stage0_61[150]},
      {stage1_61[79]}
   );
   gpc1_1 gpc2012 (
      {stage0_61[151]},
      {stage1_61[80]}
   );
   gpc1_1 gpc2013 (
      {stage0_61[152]},
      {stage1_61[81]}
   );
   gpc1_1 gpc2014 (
      {stage0_61[153]},
      {stage1_61[82]}
   );
   gpc1_1 gpc2015 (
      {stage0_61[154]},
      {stage1_61[83]}
   );
   gpc1_1 gpc2016 (
      {stage0_61[155]},
      {stage1_61[84]}
   );
   gpc1_1 gpc2017 (
      {stage0_61[156]},
      {stage1_61[85]}
   );
   gpc1_1 gpc2018 (
      {stage0_61[157]},
      {stage1_61[86]}
   );
   gpc1_1 gpc2019 (
      {stage0_61[158]},
      {stage1_61[87]}
   );
   gpc1_1 gpc2020 (
      {stage0_61[159]},
      {stage1_61[88]}
   );
   gpc1_1 gpc2021 (
      {stage0_61[160]},
      {stage1_61[89]}
   );
   gpc1_1 gpc2022 (
      {stage0_61[161]},
      {stage1_61[90]}
   );
   gpc1_1 gpc2023 (
      {stage0_62[126]},
      {stage1_62[51]}
   );
   gpc1_1 gpc2024 (
      {stage0_62[127]},
      {stage1_62[52]}
   );
   gpc1_1 gpc2025 (
      {stage0_62[128]},
      {stage1_62[53]}
   );
   gpc1_1 gpc2026 (
      {stage0_62[129]},
      {stage1_62[54]}
   );
   gpc1_1 gpc2027 (
      {stage0_62[130]},
      {stage1_62[55]}
   );
   gpc1_1 gpc2028 (
      {stage0_62[131]},
      {stage1_62[56]}
   );
   gpc1_1 gpc2029 (
      {stage0_62[132]},
      {stage1_62[57]}
   );
   gpc1_1 gpc2030 (
      {stage0_62[133]},
      {stage1_62[58]}
   );
   gpc1_1 gpc2031 (
      {stage0_62[134]},
      {stage1_62[59]}
   );
   gpc1_1 gpc2032 (
      {stage0_62[135]},
      {stage1_62[60]}
   );
   gpc1_1 gpc2033 (
      {stage0_62[136]},
      {stage1_62[61]}
   );
   gpc1_1 gpc2034 (
      {stage0_62[137]},
      {stage1_62[62]}
   );
   gpc1_1 gpc2035 (
      {stage0_62[138]},
      {stage1_62[63]}
   );
   gpc1_1 gpc2036 (
      {stage0_62[139]},
      {stage1_62[64]}
   );
   gpc1_1 gpc2037 (
      {stage0_62[140]},
      {stage1_62[65]}
   );
   gpc1_1 gpc2038 (
      {stage0_62[141]},
      {stage1_62[66]}
   );
   gpc1_1 gpc2039 (
      {stage0_62[142]},
      {stage1_62[67]}
   );
   gpc1_1 gpc2040 (
      {stage0_62[143]},
      {stage1_62[68]}
   );
   gpc1_1 gpc2041 (
      {stage0_62[144]},
      {stage1_62[69]}
   );
   gpc1_1 gpc2042 (
      {stage0_62[145]},
      {stage1_62[70]}
   );
   gpc1_1 gpc2043 (
      {stage0_62[146]},
      {stage1_62[71]}
   );
   gpc1_1 gpc2044 (
      {stage0_62[147]},
      {stage1_62[72]}
   );
   gpc1_1 gpc2045 (
      {stage0_62[148]},
      {stage1_62[73]}
   );
   gpc1_1 gpc2046 (
      {stage0_62[149]},
      {stage1_62[74]}
   );
   gpc1_1 gpc2047 (
      {stage0_62[150]},
      {stage1_62[75]}
   );
   gpc1_1 gpc2048 (
      {stage0_62[151]},
      {stage1_62[76]}
   );
   gpc1_1 gpc2049 (
      {stage0_62[152]},
      {stage1_62[77]}
   );
   gpc1_1 gpc2050 (
      {stage0_62[153]},
      {stage1_62[78]}
   );
   gpc1_1 gpc2051 (
      {stage0_62[154]},
      {stage1_62[79]}
   );
   gpc1_1 gpc2052 (
      {stage0_62[155]},
      {stage1_62[80]}
   );
   gpc1_1 gpc2053 (
      {stage0_62[156]},
      {stage1_62[81]}
   );
   gpc1_1 gpc2054 (
      {stage0_62[157]},
      {stage1_62[82]}
   );
   gpc1_1 gpc2055 (
      {stage0_62[158]},
      {stage1_62[83]}
   );
   gpc1_1 gpc2056 (
      {stage0_62[159]},
      {stage1_62[84]}
   );
   gpc1_1 gpc2057 (
      {stage0_62[160]},
      {stage1_62[85]}
   );
   gpc1_1 gpc2058 (
      {stage0_62[161]},
      {stage1_62[86]}
   );
   gpc1_1 gpc2059 (
      {stage0_63[144]},
      {stage1_63[45]}
   );
   gpc1_1 gpc2060 (
      {stage0_63[145]},
      {stage1_63[46]}
   );
   gpc1_1 gpc2061 (
      {stage0_63[146]},
      {stage1_63[47]}
   );
   gpc1_1 gpc2062 (
      {stage0_63[147]},
      {stage1_63[48]}
   );
   gpc1_1 gpc2063 (
      {stage0_63[148]},
      {stage1_63[49]}
   );
   gpc1_1 gpc2064 (
      {stage0_63[149]},
      {stage1_63[50]}
   );
   gpc1_1 gpc2065 (
      {stage0_63[150]},
      {stage1_63[51]}
   );
   gpc1_1 gpc2066 (
      {stage0_63[151]},
      {stage1_63[52]}
   );
   gpc1_1 gpc2067 (
      {stage0_63[152]},
      {stage1_63[53]}
   );
   gpc1_1 gpc2068 (
      {stage0_63[153]},
      {stage1_63[54]}
   );
   gpc1_1 gpc2069 (
      {stage0_63[154]},
      {stage1_63[55]}
   );
   gpc1_1 gpc2070 (
      {stage0_63[155]},
      {stage1_63[56]}
   );
   gpc1_1 gpc2071 (
      {stage0_63[156]},
      {stage1_63[57]}
   );
   gpc1_1 gpc2072 (
      {stage0_63[157]},
      {stage1_63[58]}
   );
   gpc1_1 gpc2073 (
      {stage0_63[158]},
      {stage1_63[59]}
   );
   gpc1_1 gpc2074 (
      {stage0_63[159]},
      {stage1_63[60]}
   );
   gpc1_1 gpc2075 (
      {stage0_63[160]},
      {stage1_63[61]}
   );
   gpc1_1 gpc2076 (
      {stage0_63[161]},
      {stage1_63[62]}
   );
   gpc1163_5 gpc2077 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc2078 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc2079 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc2080 (
      {stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc606_5 gpc2081 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc615_5 gpc2082 (
      {stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24], stage1_0[25]},
      {stage1_1[18]},
      {stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc615_5 gpc2083 (
      {stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29], stage1_0[30]},
      {stage1_1[19]},
      {stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc606_5 gpc2084 (
      {stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25]},
      {stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8]},
      {stage2_5[0],stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7]}
   );
   gpc606_5 gpc2085 (
      {stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31]},
      {stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14]},
      {stage2_5[1],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc606_5 gpc2086 (
      {stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37]},
      {stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20]},
      {stage2_5[2],stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9]}
   );
   gpc1163_5 gpc2087 (
      {stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_5[0]},
      {stage1_6[0]},
      {stage2_7[0],stage2_6[0],stage2_5[3],stage2_4[10],stage2_3[10]}
   );
   gpc615_5 gpc2088 (
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28]},
      {stage1_4[6]},
      {stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5], stage1_5[6]},
      {stage2_7[1],stage2_6[1],stage2_5[4],stage2_4[11],stage2_3[11]}
   );
   gpc615_5 gpc2089 (
      {stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage1_4[7]},
      {stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11], stage1_5[12]},
      {stage2_7[2],stage2_6[2],stage2_5[5],stage2_4[12],stage2_3[12]}
   );
   gpc615_5 gpc2090 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38]},
      {stage1_4[8]},
      {stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17], stage1_5[18]},
      {stage2_7[3],stage2_6[3],stage2_5[6],stage2_4[13],stage2_3[13]}
   );
   gpc615_5 gpc2091 (
      {stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage1_4[9]},
      {stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23], stage1_5[24]},
      {stage2_7[4],stage2_6[4],stage2_5[7],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc2092 (
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48]},
      {stage1_4[10]},
      {stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29], stage1_5[30]},
      {stage2_7[5],stage2_6[5],stage2_5[8],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc2093 (
      {stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage1_4[11]},
      {stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36]},
      {stage2_7[6],stage2_6[6],stage2_5[9],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc2094 (
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58]},
      {stage1_4[12]},
      {stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42]},
      {stage2_7[7],stage2_6[7],stage2_5[10],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc2095 (
      {stage1_3[59], stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63]},
      {stage1_4[13]},
      {stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48]},
      {stage2_7[8],stage2_6[8],stage2_5[11],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc2096 (
      {stage1_3[64], stage1_3[65], stage1_3[66], stage1_3[67], stage1_3[68]},
      {stage1_4[14]},
      {stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53], stage1_5[54]},
      {stage2_7[9],stage2_6[9],stage2_5[12],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc2097 (
      {stage1_3[69], stage1_3[70], stage1_3[71], stage1_3[72], stage1_3[73]},
      {stage1_4[15]},
      {stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59], stage1_5[60]},
      {stage2_7[10],stage2_6[10],stage2_5[13],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc2098 (
      {stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77], stage1_3[78]},
      {stage1_4[16]},
      {stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66]},
      {stage2_7[11],stage2_6[11],stage2_5[14],stage2_4[21],stage2_3[21]}
   );
   gpc615_5 gpc2099 (
      {stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83]},
      {stage1_4[17]},
      {stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71], stage1_5[72]},
      {stage2_7[12],stage2_6[12],stage2_5[15],stage2_4[22],stage2_3[22]}
   );
   gpc606_5 gpc2100 (
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[0],stage2_7[13],stage2_6[13],stage2_5[16],stage2_4[23]}
   );
   gpc606_5 gpc2101 (
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[1],stage2_7[14],stage2_6[14],stage2_5[17],stage2_4[24]}
   );
   gpc606_5 gpc2102 (
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[2],stage2_7[15],stage2_6[15],stage2_5[18],stage2_4[25]}
   );
   gpc606_5 gpc2103 (
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[3],stage2_7[16],stage2_6[16],stage2_5[19],stage2_4[26]}
   );
   gpc606_5 gpc2104 (
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[4],stage2_7[17],stage2_6[17],stage2_5[20],stage2_4[27]}
   );
   gpc606_5 gpc2105 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[5],stage2_7[18],stage2_6[18],stage2_5[21],stage2_4[28]}
   );
   gpc606_5 gpc2106 (
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[6],stage2_7[19],stage2_6[19],stage2_5[22],stage2_4[29]}
   );
   gpc606_5 gpc2107 (
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage2_8[7],stage2_7[20],stage2_6[20],stage2_5[23],stage2_4[30]}
   );
   gpc606_5 gpc2108 (
      {stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77], stage1_5[78]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[8],stage2_7[21],stage2_6[21],stage2_5[24]}
   );
   gpc606_5 gpc2109 (
      {stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83], stage1_5[84]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[9],stage2_7[22],stage2_6[22],stage2_5[25]}
   );
   gpc606_5 gpc2110 (
      {stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89], stage1_5[90]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[10],stage2_7[23],stage2_6[23],stage2_5[26]}
   );
   gpc606_5 gpc2111 (
      {stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95], stage1_5[96]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[11],stage2_7[24],stage2_6[24],stage2_5[27]}
   );
   gpc606_5 gpc2112 (
      {stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101], stage1_5[102]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[12],stage2_7[25],stage2_6[25],stage2_5[28]}
   );
   gpc606_5 gpc2113 (
      {stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107], stage1_5[108]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[13],stage2_7[26],stage2_6[26],stage2_5[29]}
   );
   gpc615_5 gpc2114 (
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage1_7[36]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[6],stage2_8[14],stage2_7[27],stage2_6[27]}
   );
   gpc615_5 gpc2115 (
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], 1'b0},
      {stage1_7[37]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[7],stage2_8[15],stage2_7[28],stage2_6[28]}
   );
   gpc606_5 gpc2116 (
      {stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[2],stage2_9[8],stage2_8[16],stage2_7[29]}
   );
   gpc615_5 gpc2117 (
      {stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47], stage1_7[48]},
      {stage1_8[12]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[3],stage2_9[9],stage2_8[17],stage2_7[30]}
   );
   gpc615_5 gpc2118 (
      {stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage1_8[13]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[4],stage2_9[10],stage2_8[18],stage2_7[31]}
   );
   gpc615_5 gpc2119 (
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58]},
      {stage1_8[14]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[5],stage2_9[11],stage2_8[19],stage2_7[32]}
   );
   gpc615_5 gpc2120 (
      {stage1_7[59], stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63]},
      {stage1_8[15]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[6],stage2_9[12],stage2_8[20],stage2_7[33]}
   );
   gpc606_5 gpc2121 (
      {stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[5],stage2_10[7],stage2_9[13],stage2_8[21]}
   );
   gpc606_5 gpc2122 (
      {stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[6],stage2_10[8],stage2_9[14],stage2_8[22]}
   );
   gpc606_5 gpc2123 (
      {stage1_8[28], stage1_8[29], stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[7],stage2_10[9],stage2_9[15],stage2_8[23]}
   );
   gpc606_5 gpc2124 (
      {stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[8],stage2_10[10],stage2_9[16],stage2_8[24]}
   );
   gpc606_5 gpc2125 (
      {stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[9],stage2_10[11],stage2_9[17],stage2_8[25]}
   );
   gpc606_5 gpc2126 (
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[5],stage2_11[10],stage2_10[12],stage2_9[18]}
   );
   gpc606_5 gpc2127 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[6],stage2_11[11],stage2_10[13],stage2_9[19]}
   );
   gpc606_5 gpc2128 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[7],stage2_11[12],stage2_10[14],stage2_9[20]}
   );
   gpc606_5 gpc2129 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[8],stage2_11[13],stage2_10[15],stage2_9[21]}
   );
   gpc606_5 gpc2130 (
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[4],stage2_12[9],stage2_11[14],stage2_10[16]}
   );
   gpc606_5 gpc2131 (
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[5],stage2_12[10],stage2_11[15],stage2_10[17]}
   );
   gpc606_5 gpc2132 (
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[6],stage2_12[11],stage2_11[16],stage2_10[18]}
   );
   gpc606_5 gpc2133 (
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[7],stage2_12[12],stage2_11[17],stage2_10[19]}
   );
   gpc615_5 gpc2134 (
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58]},
      {stage1_11[24]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[8],stage2_12[13],stage2_11[18],stage2_10[20]}
   );
   gpc615_5 gpc2135 (
      {stage1_10[59], stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63]},
      {stage1_11[25]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[9],stage2_12[14],stage2_11[19],stage2_10[21]}
   );
   gpc615_5 gpc2136 (
      {stage1_10[64], stage1_10[65], stage1_10[66], stage1_10[67], stage1_10[68]},
      {stage1_11[26]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[10],stage2_12[15],stage2_11[20],stage2_10[22]}
   );
   gpc615_5 gpc2137 (
      {stage1_10[69], stage1_10[70], stage1_10[71], stage1_10[72], stage1_10[73]},
      {stage1_11[27]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[11],stage2_12[16],stage2_11[21],stage2_10[23]}
   );
   gpc615_5 gpc2138 (
      {stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77], stage1_10[78]},
      {stage1_11[28]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[12],stage2_12[17],stage2_11[22],stage2_10[24]}
   );
   gpc615_5 gpc2139 (
      {stage1_11[29], stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33]},
      {stage1_12[54]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[9],stage2_13[13],stage2_12[18],stage2_11[23]}
   );
   gpc615_5 gpc2140 (
      {stage1_11[34], stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38]},
      {stage1_12[55]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[10],stage2_13[14],stage2_12[19],stage2_11[24]}
   );
   gpc615_5 gpc2141 (
      {stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43]},
      {stage1_12[56]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[11],stage2_13[15],stage2_12[20],stage2_11[25]}
   );
   gpc615_5 gpc2142 (
      {stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_12[57]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[12],stage2_13[16],stage2_12[21],stage2_11[26]}
   );
   gpc615_5 gpc2143 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage1_12[58]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[13],stage2_13[17],stage2_12[22],stage2_11[27]}
   );
   gpc615_5 gpc2144 (
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58]},
      {stage1_12[59]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[14],stage2_13[18],stage2_12[23],stage2_11[28]}
   );
   gpc615_5 gpc2145 (
      {stage1_11[59], stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63]},
      {stage1_12[60]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[15],stage2_13[19],stage2_12[24],stage2_11[29]}
   );
   gpc615_5 gpc2146 (
      {stage1_11[64], stage1_11[65], stage1_11[66], stage1_11[67], stage1_11[68]},
      {stage1_12[61]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[16],stage2_13[20],stage2_12[25],stage2_11[30]}
   );
   gpc615_5 gpc2147 (
      {stage1_11[69], stage1_11[70], stage1_11[71], stage1_11[72], stage1_11[73]},
      {stage1_12[62]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[17],stage2_13[21],stage2_12[26],stage2_11[31]}
   );
   gpc606_5 gpc2148 (
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[9],stage2_14[18],stage2_13[22]}
   );
   gpc606_5 gpc2149 (
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[1],stage2_15[10],stage2_14[19],stage2_13[23]}
   );
   gpc615_5 gpc2150 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4]},
      {stage1_15[12]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[2],stage2_16[2],stage2_15[11],stage2_14[20]}
   );
   gpc615_5 gpc2151 (
      {stage1_14[5], stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9]},
      {stage1_15[13]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[3],stage2_16[3],stage2_15[12],stage2_14[21]}
   );
   gpc606_5 gpc2152 (
      {stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[4],stage2_16[4],stage2_15[13]}
   );
   gpc606_5 gpc2153 (
      {stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23], stage1_15[24], stage1_15[25]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[3],stage2_17[5],stage2_16[5],stage2_15[14]}
   );
   gpc606_5 gpc2154 (
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[4],stage2_17[6],stage2_16[6],stage2_15[15]}
   );
   gpc606_5 gpc2155 (
      {stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[5],stage2_17[7],stage2_16[7],stage2_15[16]}
   );
   gpc606_5 gpc2156 (
      {stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[6],stage2_17[8],stage2_16[8],stage2_15[17]}
   );
   gpc606_5 gpc2157 (
      {stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47], stage1_15[48], stage1_15[49]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[7],stage2_17[9],stage2_16[9],stage2_15[18]}
   );
   gpc606_5 gpc2158 (
      {stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53], stage1_15[54], stage1_15[55]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[8],stage2_17[10],stage2_16[10],stage2_15[19]}
   );
   gpc606_5 gpc2159 (
      {stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59], stage1_15[60], stage1_15[61]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[9],stage2_17[11],stage2_16[11],stage2_15[20]}
   );
   gpc606_5 gpc2160 (
      {stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65], stage1_15[66], stage1_15[67]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[10],stage2_17[12],stage2_16[12],stage2_15[21]}
   );
   gpc606_5 gpc2161 (
      {stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71], stage1_15[72], stage1_15[73]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[11],stage2_17[13],stage2_16[13],stage2_15[22]}
   );
   gpc606_5 gpc2162 (
      {stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77], stage1_15[78], stage1_15[79]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage2_19[10],stage2_18[12],stage2_17[14],stage2_16[14],stage2_15[23]}
   );
   gpc606_5 gpc2163 (
      {stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83], stage1_15[84], stage1_15[85]},
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage2_19[11],stage2_18[13],stage2_17[15],stage2_16[15],stage2_15[24]}
   );
   gpc606_5 gpc2164 (
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[12],stage2_18[14],stage2_17[16],stage2_16[16]}
   );
   gpc606_5 gpc2165 (
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[13],stage2_18[15],stage2_17[17],stage2_16[17]}
   );
   gpc606_5 gpc2166 (
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[14],stage2_18[16],stage2_17[18],stage2_16[18]}
   );
   gpc606_5 gpc2167 (
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[15],stage2_18[17],stage2_17[19],stage2_16[19]}
   );
   gpc606_5 gpc2168 (
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[16],stage2_18[18],stage2_17[20],stage2_16[20]}
   );
   gpc606_5 gpc2169 (
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[5],stage2_19[17],stage2_18[19],stage2_17[21]}
   );
   gpc606_5 gpc2170 (
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[6],stage2_19[18],stage2_18[20],stage2_17[22]}
   );
   gpc606_5 gpc2171 (
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[7],stage2_19[19],stage2_18[21],stage2_17[23]}
   );
   gpc615_5 gpc2172 (
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94]},
      {stage1_18[30]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[8],stage2_19[20],stage2_18[22],stage2_17[24]}
   );
   gpc615_5 gpc2173 (
      {stage1_17[95], stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99]},
      {stage1_18[31]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[9],stage2_19[21],stage2_18[23],stage2_17[25]}
   );
   gpc615_5 gpc2174 (
      {stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35], stage1_18[36]},
      {stage1_19[30]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[5],stage2_20[10],stage2_19[22],stage2_18[24]}
   );
   gpc615_5 gpc2175 (
      {stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage1_19[31]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[6],stage2_20[11],stage2_19[23],stage2_18[25]}
   );
   gpc615_5 gpc2176 (
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46]},
      {stage1_19[32]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[7],stage2_20[12],stage2_19[24],stage2_18[26]}
   );
   gpc615_5 gpc2177 (
      {stage1_19[33], stage1_19[34], stage1_19[35], stage1_19[36], stage1_19[37]},
      {stage1_20[18]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[3],stage2_21[8],stage2_20[13],stage2_19[25]}
   );
   gpc615_5 gpc2178 (
      {stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41], stage1_19[42]},
      {stage1_20[19]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[4],stage2_21[9],stage2_20[14],stage2_19[26]}
   );
   gpc615_5 gpc2179 (
      {stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage1_20[20]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[5],stage2_21[10],stage2_20[15],stage2_19[27]}
   );
   gpc606_5 gpc2180 (
      {stage1_20[21], stage1_20[22], stage1_20[23], stage1_20[24], stage1_20[25], stage1_20[26]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[3],stage2_22[6],stage2_21[11],stage2_20[16]}
   );
   gpc606_5 gpc2181 (
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[1],stage2_23[4],stage2_22[7],stage2_21[12]}
   );
   gpc606_5 gpc2182 (
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[2],stage2_23[5],stage2_22[8],stage2_21[13]}
   );
   gpc606_5 gpc2183 (
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[3],stage2_23[6],stage2_22[9],stage2_21[14]}
   );
   gpc606_5 gpc2184 (
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[4],stage2_23[7],stage2_22[10],stage2_21[15]}
   );
   gpc606_5 gpc2185 (
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[5],stage2_23[8],stage2_22[11],stage2_21[16]}
   );
   gpc1163_5 gpc2186 (
      {stage1_22[6], stage1_22[7], stage1_22[8]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage1_24[0]},
      {stage1_25[0]},
      {stage2_26[0],stage2_25[5],stage2_24[6],stage2_23[9],stage2_22[12]}
   );
   gpc1163_5 gpc2187 (
      {stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage1_24[1]},
      {stage1_25[1]},
      {stage2_26[1],stage2_25[6],stage2_24[7],stage2_23[10],stage2_22[13]}
   );
   gpc1163_5 gpc2188 (
      {stage1_22[12], stage1_22[13], stage1_22[14]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage1_24[2]},
      {stage1_25[2]},
      {stage2_26[2],stage2_25[7],stage2_24[8],stage2_23[11],stage2_22[14]}
   );
   gpc1163_5 gpc2189 (
      {stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage1_24[3]},
      {stage1_25[3]},
      {stage2_26[3],stage2_25[8],stage2_24[9],stage2_23[12],stage2_22[15]}
   );
   gpc1163_5 gpc2190 (
      {stage1_22[18], stage1_22[19], stage1_22[20]},
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage1_24[4]},
      {stage1_25[4]},
      {stage2_26[4],stage2_25[9],stage2_24[10],stage2_23[13],stage2_22[16]}
   );
   gpc1163_5 gpc2191 (
      {stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage1_24[5]},
      {stage1_25[5]},
      {stage2_26[5],stage2_25[10],stage2_24[11],stage2_23[14],stage2_22[17]}
   );
   gpc1163_5 gpc2192 (
      {stage1_22[24], stage1_22[25], stage1_22[26]},
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage1_24[6]},
      {stage1_25[6]},
      {stage2_26[6],stage2_25[11],stage2_24[12],stage2_23[15],stage2_22[18]}
   );
   gpc615_5 gpc2193 (
      {stage1_22[27], stage1_22[28], stage1_22[29], stage1_22[30], stage1_22[31]},
      {stage1_23[72]},
      {stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12]},
      {stage2_26[7],stage2_25[12],stage2_24[13],stage2_23[16],stage2_22[19]}
   );
   gpc615_5 gpc2194 (
      {stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35], stage1_22[36]},
      {stage1_23[73]},
      {stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18]},
      {stage2_26[8],stage2_25[13],stage2_24[14],stage2_23[17],stage2_22[20]}
   );
   gpc615_5 gpc2195 (
      {stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage1_23[74]},
      {stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23], stage1_24[24]},
      {stage2_26[9],stage2_25[14],stage2_24[15],stage2_23[18],stage2_22[21]}
   );
   gpc615_5 gpc2196 (
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46]},
      {stage1_23[75]},
      {stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29], stage1_24[30]},
      {stage2_26[10],stage2_25[15],stage2_24[16],stage2_23[19],stage2_22[22]}
   );
   gpc615_5 gpc2197 (
      {stage1_22[47], stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51]},
      {stage1_23[76]},
      {stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35], stage1_24[36]},
      {stage2_26[11],stage2_25[16],stage2_24[17],stage2_23[20],stage2_22[23]}
   );
   gpc615_5 gpc2198 (
      {stage1_22[52], stage1_22[53], stage1_22[54], stage1_22[55], stage1_22[56]},
      {stage1_23[77]},
      {stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41], stage1_24[42]},
      {stage2_26[12],stage2_25[17],stage2_24[18],stage2_23[21],stage2_22[24]}
   );
   gpc615_5 gpc2199 (
      {stage1_22[57], stage1_22[58], stage1_22[59], stage1_22[60], stage1_22[61]},
      {stage1_23[78]},
      {stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47], stage1_24[48]},
      {stage2_26[13],stage2_25[18],stage2_24[19],stage2_23[22],stage2_22[25]}
   );
   gpc606_5 gpc2200 (
      {stage1_23[79], stage1_23[80], stage1_23[81], stage1_23[82], stage1_23[83], stage1_23[84]},
      {stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12]},
      {stage2_27[0],stage2_26[14],stage2_25[19],stage2_24[20],stage2_23[23]}
   );
   gpc606_5 gpc2201 (
      {stage1_23[85], stage1_23[86], stage1_23[87], stage1_23[88], stage1_23[89], stage1_23[90]},
      {stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17], stage1_25[18]},
      {stage2_27[1],stage2_26[15],stage2_25[20],stage2_24[21],stage2_23[24]}
   );
   gpc606_5 gpc2202 (
      {stage1_23[91], stage1_23[92], stage1_23[93], stage1_23[94], stage1_23[95], stage1_23[96]},
      {stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23], stage1_25[24]},
      {stage2_27[2],stage2_26[16],stage2_25[21],stage2_24[22],stage2_23[25]}
   );
   gpc606_5 gpc2203 (
      {stage1_23[97], stage1_23[98], stage1_23[99], stage1_23[100], stage1_23[101], stage1_23[102]},
      {stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29], stage1_25[30]},
      {stage2_27[3],stage2_26[17],stage2_25[22],stage2_24[23],stage2_23[26]}
   );
   gpc606_5 gpc2204 (
      {stage1_23[103], stage1_23[104], stage1_23[105], stage1_23[106], stage1_23[107], stage1_23[108]},
      {stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35], stage1_25[36]},
      {stage2_27[4],stage2_26[18],stage2_25[23],stage2_24[24],stage2_23[27]}
   );
   gpc606_5 gpc2205 (
      {stage1_23[109], stage1_23[110], stage1_23[111], stage1_23[112], stage1_23[113], stage1_23[114]},
      {stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41], stage1_25[42]},
      {stage2_27[5],stage2_26[19],stage2_25[24],stage2_24[25],stage2_23[28]}
   );
   gpc606_5 gpc2206 (
      {stage1_23[115], stage1_23[116], stage1_23[117], stage1_23[118], stage1_23[119], stage1_23[120]},
      {stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47], stage1_25[48]},
      {stage2_27[6],stage2_26[20],stage2_25[25],stage2_24[26],stage2_23[29]}
   );
   gpc606_5 gpc2207 (
      {stage1_23[121], stage1_23[122], stage1_23[123], stage1_23[124], stage1_23[125], stage1_23[126]},
      {stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53], stage1_25[54]},
      {stage2_27[7],stage2_26[21],stage2_25[26],stage2_24[27],stage2_23[30]}
   );
   gpc615_5 gpc2208 (
      {stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53]},
      {stage1_25[55]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[8],stage2_26[22],stage2_25[27],stage2_24[28]}
   );
   gpc615_5 gpc2209 (
      {stage1_24[54], stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58]},
      {stage1_25[56]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[9],stage2_26[23],stage2_25[28],stage2_24[29]}
   );
   gpc615_5 gpc2210 (
      {stage1_24[59], stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63]},
      {stage1_25[57]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[10],stage2_26[24],stage2_25[29],stage2_24[30]}
   );
   gpc615_5 gpc2211 (
      {stage1_24[64], stage1_24[65], stage1_24[66], stage1_24[67], stage1_24[68]},
      {stage1_25[58]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[11],stage2_26[25],stage2_25[30],stage2_24[31]}
   );
   gpc606_5 gpc2212 (
      {stage1_25[59], stage1_25[60], stage1_25[61], stage1_25[62], stage1_25[63], stage1_25[64]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[4],stage2_27[12],stage2_26[26],stage2_25[31]}
   );
   gpc606_5 gpc2213 (
      {stage1_25[65], stage1_25[66], stage1_25[67], stage1_25[68], stage1_25[69], stage1_25[70]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[5],stage2_27[13],stage2_26[27],stage2_25[32]}
   );
   gpc606_5 gpc2214 (
      {stage1_25[71], stage1_25[72], stage1_25[73], stage1_25[74], stage1_25[75], stage1_25[76]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[6],stage2_27[14],stage2_26[28],stage2_25[33]}
   );
   gpc606_5 gpc2215 (
      {stage1_25[77], stage1_25[78], stage1_25[79], stage1_25[80], stage1_25[81], stage1_25[82]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[7],stage2_27[15],stage2_26[29],stage2_25[34]}
   );
   gpc2116_5 gpc2216 (
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage1_27[24]},
      {stage1_28[0]},
      {stage1_29[0], stage1_29[1]},
      {stage2_30[0],stage2_29[4],stage2_28[8],stage2_27[16],stage2_26[30]}
   );
   gpc2116_5 gpc2217 (
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage1_27[25]},
      {stage1_28[1]},
      {stage1_29[2], stage1_29[3]},
      {stage2_30[1],stage2_29[5],stage2_28[9],stage2_27[17],stage2_26[31]}
   );
   gpc2116_5 gpc2218 (
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage1_27[26]},
      {stage1_28[2]},
      {stage1_29[4], stage1_29[5]},
      {stage2_30[2],stage2_29[6],stage2_28[10],stage2_27[18],stage2_26[32]}
   );
   gpc2116_5 gpc2219 (
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage1_27[27]},
      {stage1_28[3]},
      {stage1_29[6], stage1_29[7]},
      {stage2_30[3],stage2_29[7],stage2_28[11],stage2_27[19],stage2_26[33]}
   );
   gpc2116_5 gpc2220 (
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage1_27[28]},
      {stage1_28[4]},
      {stage1_29[8], stage1_29[9]},
      {stage2_30[4],stage2_29[8],stage2_28[12],stage2_27[20],stage2_26[34]}
   );
   gpc615_5 gpc2221 (
      {stage1_27[29], stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33]},
      {stage1_28[5]},
      {stage1_29[10], stage1_29[11], stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15]},
      {stage2_31[0],stage2_30[5],stage2_29[9],stage2_28[13],stage2_27[21]}
   );
   gpc615_5 gpc2222 (
      {stage1_27[34], stage1_27[35], stage1_27[36], stage1_27[37], stage1_27[38]},
      {stage1_28[6]},
      {stage1_29[16], stage1_29[17], stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21]},
      {stage2_31[1],stage2_30[6],stage2_29[10],stage2_28[14],stage2_27[22]}
   );
   gpc615_5 gpc2223 (
      {stage1_27[39], stage1_27[40], stage1_27[41], stage1_27[42], stage1_27[43]},
      {stage1_28[7]},
      {stage1_29[22], stage1_29[23], stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27]},
      {stage2_31[2],stage2_30[7],stage2_29[11],stage2_28[15],stage2_27[23]}
   );
   gpc615_5 gpc2224 (
      {stage1_27[44], stage1_27[45], stage1_27[46], stage1_27[47], stage1_27[48]},
      {stage1_28[8]},
      {stage1_29[28], stage1_29[29], stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33]},
      {stage2_31[3],stage2_30[8],stage2_29[12],stage2_28[16],stage2_27[24]}
   );
   gpc606_5 gpc2225 (
      {stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12], stage1_28[13], stage1_28[14]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[4],stage2_30[9],stage2_29[13],stage2_28[17]}
   );
   gpc606_5 gpc2226 (
      {stage1_28[15], stage1_28[16], stage1_28[17], stage1_28[18], stage1_28[19], stage1_28[20]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[5],stage2_30[10],stage2_29[14],stage2_28[18]}
   );
   gpc606_5 gpc2227 (
      {stage1_28[21], stage1_28[22], stage1_28[23], stage1_28[24], stage1_28[25], stage1_28[26]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[6],stage2_30[11],stage2_29[15],stage2_28[19]}
   );
   gpc606_5 gpc2228 (
      {stage1_28[27], stage1_28[28], stage1_28[29], stage1_28[30], stage1_28[31], stage1_28[32]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[7],stage2_30[12],stage2_29[16],stage2_28[20]}
   );
   gpc606_5 gpc2229 (
      {stage1_28[33], stage1_28[34], stage1_28[35], stage1_28[36], stage1_28[37], stage1_28[38]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[8],stage2_30[13],stage2_29[17],stage2_28[21]}
   );
   gpc606_5 gpc2230 (
      {stage1_28[39], stage1_28[40], stage1_28[41], stage1_28[42], stage1_28[43], stage1_28[44]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[9],stage2_30[14],stage2_29[18],stage2_28[22]}
   );
   gpc606_5 gpc2231 (
      {stage1_28[45], stage1_28[46], stage1_28[47], stage1_28[48], stage1_28[49], stage1_28[50]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[10],stage2_30[15],stage2_29[19],stage2_28[23]}
   );
   gpc606_5 gpc2232 (
      {stage1_28[51], stage1_28[52], stage1_28[53], stage1_28[54], stage1_28[55], stage1_28[56]},
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage2_32[7],stage2_31[11],stage2_30[16],stage2_29[20],stage2_28[24]}
   );
   gpc606_5 gpc2233 (
      {stage1_28[57], stage1_28[58], stage1_28[59], stage1_28[60], stage1_28[61], stage1_28[62]},
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage2_32[8],stage2_31[12],stage2_30[17],stage2_29[21],stage2_28[25]}
   );
   gpc606_5 gpc2234 (
      {stage1_28[63], stage1_28[64], stage1_28[65], stage1_28[66], stage1_28[67], stage1_28[68]},
      {stage1_30[54], stage1_30[55], stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59]},
      {stage2_32[9],stage2_31[13],stage2_30[18],stage2_29[22],stage2_28[26]}
   );
   gpc606_5 gpc2235 (
      {stage1_29[34], stage1_29[35], stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[10],stage2_31[14],stage2_30[19],stage2_29[23]}
   );
   gpc606_5 gpc2236 (
      {stage1_29[40], stage1_29[41], stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[11],stage2_31[15],stage2_30[20],stage2_29[24]}
   );
   gpc606_5 gpc2237 (
      {stage1_29[46], stage1_29[47], stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[12],stage2_31[16],stage2_30[21],stage2_29[25]}
   );
   gpc606_5 gpc2238 (
      {stage1_29[52], stage1_29[53], stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[13],stage2_31[17],stage2_30[22],stage2_29[26]}
   );
   gpc606_5 gpc2239 (
      {stage1_30[60], stage1_30[61], stage1_30[62], stage1_30[63], stage1_30[64], stage1_30[65]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[4],stage2_32[14],stage2_31[18],stage2_30[23]}
   );
   gpc606_5 gpc2240 (
      {stage1_30[66], stage1_30[67], stage1_30[68], stage1_30[69], stage1_30[70], stage1_30[71]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[5],stage2_32[15],stage2_31[19],stage2_30[24]}
   );
   gpc606_5 gpc2241 (
      {stage1_30[72], stage1_30[73], stage1_30[74], stage1_30[75], stage1_30[76], stage1_30[77]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[6],stage2_32[16],stage2_31[20],stage2_30[25]}
   );
   gpc606_5 gpc2242 (
      {stage1_30[78], stage1_30[79], stage1_30[80], stage1_30[81], stage1_30[82], stage1_30[83]},
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage2_34[3],stage2_33[7],stage2_32[17],stage2_31[21],stage2_30[26]}
   );
   gpc615_5 gpc2243 (
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28]},
      {stage1_32[24]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[4],stage2_33[8],stage2_32[18],stage2_31[22]}
   );
   gpc615_5 gpc2244 (
      {stage1_31[29], stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33]},
      {stage1_32[25]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[5],stage2_33[9],stage2_32[19],stage2_31[23]}
   );
   gpc615_5 gpc2245 (
      {stage1_31[34], stage1_31[35], stage1_31[36], stage1_31[37], stage1_31[38]},
      {stage1_32[26]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[6],stage2_33[10],stage2_32[20],stage2_31[24]}
   );
   gpc615_5 gpc2246 (
      {stage1_31[39], stage1_31[40], stage1_31[41], stage1_31[42], stage1_31[43]},
      {stage1_32[27]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[7],stage2_33[11],stage2_32[21],stage2_31[25]}
   );
   gpc615_5 gpc2247 (
      {stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48]},
      {stage1_32[28]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[8],stage2_33[12],stage2_32[22],stage2_31[26]}
   );
   gpc615_5 gpc2248 (
      {stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53]},
      {stage1_32[29]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage2_35[5],stage2_34[9],stage2_33[13],stage2_32[23],stage2_31[27]}
   );
   gpc615_5 gpc2249 (
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58]},
      {stage1_32[30]},
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41]},
      {stage2_35[6],stage2_34[10],stage2_33[14],stage2_32[24],stage2_31[28]}
   );
   gpc615_5 gpc2250 (
      {stage1_31[59], stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63]},
      {stage1_32[31]},
      {stage1_33[42], stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47]},
      {stage2_35[7],stage2_34[11],stage2_33[15],stage2_32[25],stage2_31[29]}
   );
   gpc615_5 gpc2251 (
      {stage1_31[64], stage1_31[65], stage1_31[66], stage1_31[67], stage1_31[68]},
      {stage1_32[32]},
      {stage1_33[48], stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53]},
      {stage2_35[8],stage2_34[12],stage2_33[16],stage2_32[26],stage2_31[30]}
   );
   gpc615_5 gpc2252 (
      {stage1_31[69], stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73]},
      {stage1_32[33]},
      {stage1_33[54], stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59]},
      {stage2_35[9],stage2_34[13],stage2_33[17],stage2_32[27],stage2_31[31]}
   );
   gpc615_5 gpc2253 (
      {stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78]},
      {stage1_32[34]},
      {stage1_33[60], stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65]},
      {stage2_35[10],stage2_34[14],stage2_33[18],stage2_32[28],stage2_31[32]}
   );
   gpc615_5 gpc2254 (
      {stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage1_32[35]},
      {stage1_33[66], stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71]},
      {stage2_35[11],stage2_34[15],stage2_33[19],stage2_32[29],stage2_31[33]}
   );
   gpc615_5 gpc2255 (
      {stage1_31[84], stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88]},
      {stage1_32[36]},
      {stage1_33[72], stage1_33[73], stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77]},
      {stage2_35[12],stage2_34[16],stage2_33[20],stage2_32[30],stage2_31[34]}
   );
   gpc615_5 gpc2256 (
      {stage1_31[89], stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93]},
      {stage1_32[37]},
      {stage1_33[78], stage1_33[79], stage1_33[80], stage1_33[81], stage1_33[82], stage1_33[83]},
      {stage2_35[13],stage2_34[17],stage2_33[21],stage2_32[31],stage2_31[35]}
   );
   gpc606_5 gpc2257 (
      {stage1_32[38], stage1_32[39], stage1_32[40], stage1_32[41], stage1_32[42], stage1_32[43]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[14],stage2_34[18],stage2_33[22],stage2_32[32]}
   );
   gpc606_5 gpc2258 (
      {stage1_32[44], stage1_32[45], stage1_32[46], stage1_32[47], stage1_32[48], stage1_32[49]},
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11]},
      {stage2_36[1],stage2_35[15],stage2_34[19],stage2_33[23],stage2_32[33]}
   );
   gpc606_5 gpc2259 (
      {stage1_32[50], stage1_32[51], stage1_32[52], stage1_32[53], stage1_32[54], stage1_32[55]},
      {stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17]},
      {stage2_36[2],stage2_35[16],stage2_34[20],stage2_33[24],stage2_32[34]}
   );
   gpc606_5 gpc2260 (
      {stage1_32[56], stage1_32[57], stage1_32[58], stage1_32[59], stage1_32[60], stage1_32[61]},
      {stage1_34[18], stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23]},
      {stage2_36[3],stage2_35[17],stage2_34[21],stage2_33[25],stage2_32[35]}
   );
   gpc606_5 gpc2261 (
      {stage1_32[62], stage1_32[63], stage1_32[64], stage1_32[65], stage1_32[66], stage1_32[67]},
      {stage1_34[24], stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29]},
      {stage2_36[4],stage2_35[18],stage2_34[22],stage2_33[26],stage2_32[36]}
   );
   gpc606_5 gpc2262 (
      {stage1_33[84], stage1_33[85], stage1_33[86], stage1_33[87], stage1_33[88], stage1_33[89]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[5],stage2_35[19],stage2_34[23],stage2_33[27]}
   );
   gpc606_5 gpc2263 (
      {stage1_34[30], stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[1],stage2_36[6],stage2_35[20],stage2_34[24]}
   );
   gpc606_5 gpc2264 (
      {stage1_34[36], stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40], stage1_34[41]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[2],stage2_36[7],stage2_35[21],stage2_34[25]}
   );
   gpc606_5 gpc2265 (
      {stage1_34[42], stage1_34[43], stage1_34[44], stage1_34[45], stage1_34[46], stage1_34[47]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[3],stage2_36[8],stage2_35[22],stage2_34[26]}
   );
   gpc615_5 gpc2266 (
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10]},
      {stage1_36[18]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[3],stage2_37[4],stage2_36[9],stage2_35[23]}
   );
   gpc615_5 gpc2267 (
      {stage1_35[11], stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15]},
      {stage1_36[19]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[4],stage2_37[5],stage2_36[10],stage2_35[24]}
   );
   gpc615_5 gpc2268 (
      {stage1_35[16], stage1_35[17], stage1_35[18], stage1_35[19], stage1_35[20]},
      {stage1_36[20]},
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage2_39[2],stage2_38[5],stage2_37[6],stage2_36[11],stage2_35[25]}
   );
   gpc615_5 gpc2269 (
      {stage1_35[21], stage1_35[22], stage1_35[23], stage1_35[24], stage1_35[25]},
      {stage1_36[21]},
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage2_39[3],stage2_38[6],stage2_37[7],stage2_36[12],stage2_35[26]}
   );
   gpc615_5 gpc2270 (
      {stage1_35[26], stage1_35[27], stage1_35[28], stage1_35[29], stage1_35[30]},
      {stage1_36[22]},
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28], stage1_37[29]},
      {stage2_39[4],stage2_38[7],stage2_37[8],stage2_36[13],stage2_35[27]}
   );
   gpc615_5 gpc2271 (
      {stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35]},
      {stage1_36[23]},
      {stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33], stage1_37[34], stage1_37[35]},
      {stage2_39[5],stage2_38[8],stage2_37[9],stage2_36[14],stage2_35[28]}
   );
   gpc615_5 gpc2272 (
      {stage1_35[36], stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40]},
      {stage1_36[24]},
      {stage1_37[36], stage1_37[37], stage1_37[38], stage1_37[39], stage1_37[40], stage1_37[41]},
      {stage2_39[6],stage2_38[9],stage2_37[10],stage2_36[15],stage2_35[29]}
   );
   gpc615_5 gpc2273 (
      {stage1_35[41], stage1_35[42], stage1_35[43], stage1_35[44], stage1_35[45]},
      {stage1_36[25]},
      {stage1_37[42], stage1_37[43], stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47]},
      {stage2_39[7],stage2_38[10],stage2_37[11],stage2_36[16],stage2_35[30]}
   );
   gpc1343_5 gpc2274 (
      {stage1_36[26], stage1_36[27], stage1_36[28]},
      {stage1_37[48], stage1_37[49], stage1_37[50], stage1_37[51]},
      {stage1_38[0], stage1_38[1], stage1_38[2]},
      {stage1_39[0]},
      {stage2_40[0],stage2_39[8],stage2_38[11],stage2_37[12],stage2_36[17]}
   );
   gpc606_5 gpc2275 (
      {stage1_36[29], stage1_36[30], stage1_36[31], stage1_36[32], stage1_36[33], stage1_36[34]},
      {stage1_38[3], stage1_38[4], stage1_38[5], stage1_38[6], stage1_38[7], stage1_38[8]},
      {stage2_40[1],stage2_39[9],stage2_38[12],stage2_37[13],stage2_36[18]}
   );
   gpc606_5 gpc2276 (
      {stage1_36[35], stage1_36[36], stage1_36[37], stage1_36[38], stage1_36[39], stage1_36[40]},
      {stage1_38[9], stage1_38[10], stage1_38[11], stage1_38[12], stage1_38[13], stage1_38[14]},
      {stage2_40[2],stage2_39[10],stage2_38[13],stage2_37[14],stage2_36[19]}
   );
   gpc606_5 gpc2277 (
      {stage1_36[41], stage1_36[42], stage1_36[43], stage1_36[44], stage1_36[45], stage1_36[46]},
      {stage1_38[15], stage1_38[16], stage1_38[17], stage1_38[18], stage1_38[19], stage1_38[20]},
      {stage2_40[3],stage2_39[11],stage2_38[14],stage2_37[15],stage2_36[20]}
   );
   gpc615_5 gpc2278 (
      {stage1_36[47], stage1_36[48], stage1_36[49], stage1_36[50], stage1_36[51]},
      {stage1_37[52]},
      {stage1_38[21], stage1_38[22], stage1_38[23], stage1_38[24], stage1_38[25], stage1_38[26]},
      {stage2_40[4],stage2_39[12],stage2_38[15],stage2_37[16],stage2_36[21]}
   );
   gpc615_5 gpc2279 (
      {stage1_36[52], stage1_36[53], stage1_36[54], stage1_36[55], stage1_36[56]},
      {stage1_37[53]},
      {stage1_38[27], stage1_38[28], stage1_38[29], stage1_38[30], stage1_38[31], stage1_38[32]},
      {stage2_40[5],stage2_39[13],stage2_38[16],stage2_37[17],stage2_36[22]}
   );
   gpc615_5 gpc2280 (
      {stage1_36[57], stage1_36[58], stage1_36[59], stage1_36[60], stage1_36[61]},
      {stage1_37[54]},
      {stage1_38[33], stage1_38[34], stage1_38[35], stage1_38[36], stage1_38[37], stage1_38[38]},
      {stage2_40[6],stage2_39[14],stage2_38[17],stage2_37[18],stage2_36[23]}
   );
   gpc615_5 gpc2281 (
      {stage1_36[62], stage1_36[63], stage1_36[64], stage1_36[65], stage1_36[66]},
      {stage1_37[55]},
      {stage1_38[39], stage1_38[40], stage1_38[41], stage1_38[42], stage1_38[43], stage1_38[44]},
      {stage2_40[7],stage2_39[15],stage2_38[18],stage2_37[19],stage2_36[24]}
   );
   gpc615_5 gpc2282 (
      {stage1_36[67], stage1_36[68], stage1_36[69], stage1_36[70], stage1_36[71]},
      {stage1_37[56]},
      {stage1_38[45], stage1_38[46], stage1_38[47], stage1_38[48], stage1_38[49], stage1_38[50]},
      {stage2_40[8],stage2_39[16],stage2_38[19],stage2_37[20],stage2_36[25]}
   );
   gpc606_5 gpc2283 (
      {stage1_37[57], stage1_37[58], stage1_37[59], stage1_37[60], stage1_37[61], stage1_37[62]},
      {stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5], stage1_39[6]},
      {stage2_41[0],stage2_40[9],stage2_39[17],stage2_38[20],stage2_37[21]}
   );
   gpc606_5 gpc2284 (
      {stage1_37[63], stage1_37[64], stage1_37[65], stage1_37[66], stage1_37[67], stage1_37[68]},
      {stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11], stage1_39[12]},
      {stage2_41[1],stage2_40[10],stage2_39[18],stage2_38[21],stage2_37[22]}
   );
   gpc606_5 gpc2285 (
      {stage1_37[69], stage1_37[70], stage1_37[71], stage1_37[72], stage1_37[73], stage1_37[74]},
      {stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17], stage1_39[18]},
      {stage2_41[2],stage2_40[11],stage2_39[19],stage2_38[22],stage2_37[23]}
   );
   gpc606_5 gpc2286 (
      {stage1_37[75], stage1_37[76], stage1_37[77], stage1_37[78], stage1_37[79], stage1_37[80]},
      {stage1_39[19], stage1_39[20], stage1_39[21], stage1_39[22], stage1_39[23], stage1_39[24]},
      {stage2_41[3],stage2_40[12],stage2_39[20],stage2_38[23],stage2_37[24]}
   );
   gpc606_5 gpc2287 (
      {stage1_37[81], stage1_37[82], stage1_37[83], stage1_37[84], stage1_37[85], stage1_37[86]},
      {stage1_39[25], stage1_39[26], stage1_39[27], stage1_39[28], stage1_39[29], stage1_39[30]},
      {stage2_41[4],stage2_40[13],stage2_39[21],stage2_38[24],stage2_37[25]}
   );
   gpc606_5 gpc2288 (
      {stage1_37[87], stage1_37[88], stage1_37[89], stage1_37[90], stage1_37[91], stage1_37[92]},
      {stage1_39[31], stage1_39[32], stage1_39[33], stage1_39[34], stage1_39[35], stage1_39[36]},
      {stage2_41[5],stage2_40[14],stage2_39[22],stage2_38[25],stage2_37[26]}
   );
   gpc606_5 gpc2289 (
      {stage1_37[93], stage1_37[94], stage1_37[95], stage1_37[96], stage1_37[97], stage1_37[98]},
      {stage1_39[37], stage1_39[38], stage1_39[39], stage1_39[40], stage1_39[41], stage1_39[42]},
      {stage2_41[6],stage2_40[15],stage2_39[23],stage2_38[26],stage2_37[27]}
   );
   gpc606_5 gpc2290 (
      {stage1_37[99], stage1_37[100], stage1_37[101], stage1_37[102], stage1_37[103], stage1_37[104]},
      {stage1_39[43], stage1_39[44], stage1_39[45], stage1_39[46], stage1_39[47], stage1_39[48]},
      {stage2_41[7],stage2_40[16],stage2_39[24],stage2_38[27],stage2_37[28]}
   );
   gpc606_5 gpc2291 (
      {stage1_37[105], stage1_37[106], stage1_37[107], stage1_37[108], stage1_37[109], stage1_37[110]},
      {stage1_39[49], stage1_39[50], stage1_39[51], stage1_39[52], stage1_39[53], stage1_39[54]},
      {stage2_41[8],stage2_40[17],stage2_39[25],stage2_38[28],stage2_37[29]}
   );
   gpc606_5 gpc2292 (
      {stage1_37[111], stage1_37[112], stage1_37[113], stage1_37[114], stage1_37[115], stage1_37[116]},
      {stage1_39[55], stage1_39[56], stage1_39[57], stage1_39[58], stage1_39[59], stage1_39[60]},
      {stage2_41[9],stage2_40[18],stage2_39[26],stage2_38[29],stage2_37[30]}
   );
   gpc615_5 gpc2293 (
      {stage1_38[51], stage1_38[52], stage1_38[53], stage1_38[54], stage1_38[55]},
      {stage1_39[61]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[10],stage2_40[19],stage2_39[27],stage2_38[30]}
   );
   gpc615_5 gpc2294 (
      {stage1_38[56], stage1_38[57], stage1_38[58], stage1_38[59], stage1_38[60]},
      {stage1_39[62]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[11],stage2_40[20],stage2_39[28],stage2_38[31]}
   );
   gpc615_5 gpc2295 (
      {stage1_38[61], stage1_38[62], stage1_38[63], stage1_38[64], stage1_38[65]},
      {stage1_39[63]},
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage2_42[2],stage2_41[12],stage2_40[21],stage2_39[29],stage2_38[32]}
   );
   gpc606_5 gpc2296 (
      {stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[0],stage2_42[3],stage2_41[13],stage2_40[22]}
   );
   gpc606_5 gpc2297 (
      {stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28], stage1_40[29]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[1],stage2_42[4],stage2_41[14],stage2_40[23]}
   );
   gpc606_5 gpc2298 (
      {stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34], stage1_40[35]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[2],stage2_42[5],stage2_41[15],stage2_40[24]}
   );
   gpc606_5 gpc2299 (
      {stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40], stage1_40[41]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[3],stage2_42[6],stage2_41[16],stage2_40[25]}
   );
   gpc606_5 gpc2300 (
      {stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46], stage1_40[47]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[4],stage2_42[7],stage2_41[17],stage2_40[26]}
   );
   gpc606_5 gpc2301 (
      {stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52], stage1_40[53]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[5],stage2_42[8],stage2_41[18],stage2_40[27]}
   );
   gpc606_5 gpc2302 (
      {stage1_40[54], stage1_40[55], stage1_40[56], stage1_40[57], stage1_40[58], stage1_40[59]},
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage2_44[6],stage2_43[6],stage2_42[9],stage2_41[19],stage2_40[28]}
   );
   gpc606_5 gpc2303 (
      {stage1_40[60], stage1_40[61], stage1_40[62], stage1_40[63], stage1_40[64], stage1_40[65]},
      {stage1_42[42], stage1_42[43], stage1_42[44], stage1_42[45], stage1_42[46], stage1_42[47]},
      {stage2_44[7],stage2_43[7],stage2_42[10],stage2_41[20],stage2_40[29]}
   );
   gpc606_5 gpc2304 (
      {stage1_40[66], stage1_40[67], stage1_40[68], stage1_40[69], stage1_40[70], stage1_40[71]},
      {stage1_42[48], stage1_42[49], stage1_42[50], stage1_42[51], stage1_42[52], stage1_42[53]},
      {stage2_44[8],stage2_43[8],stage2_42[11],stage2_41[21],stage2_40[30]}
   );
   gpc606_5 gpc2305 (
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[9],stage2_43[9],stage2_42[12],stage2_41[22]}
   );
   gpc606_5 gpc2306 (
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[10],stage2_43[10],stage2_42[13],stage2_41[23]}
   );
   gpc606_5 gpc2307 (
      {stage1_41[12], stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[11],stage2_43[11],stage2_42[14],stage2_41[24]}
   );
   gpc606_5 gpc2308 (
      {stage1_41[18], stage1_41[19], stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[12],stage2_43[12],stage2_42[15],stage2_41[25]}
   );
   gpc606_5 gpc2309 (
      {stage1_41[24], stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29]},
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage2_45[4],stage2_44[13],stage2_43[13],stage2_42[16],stage2_41[26]}
   );
   gpc606_5 gpc2310 (
      {stage1_41[30], stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34], stage1_41[35]},
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35]},
      {stage2_45[5],stage2_44[14],stage2_43[14],stage2_42[17],stage2_41[27]}
   );
   gpc606_5 gpc2311 (
      {stage1_41[36], stage1_41[37], stage1_41[38], stage1_41[39], stage1_41[40], stage1_41[41]},
      {stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39], stage1_43[40], stage1_43[41]},
      {stage2_45[6],stage2_44[15],stage2_43[15],stage2_42[18],stage2_41[28]}
   );
   gpc606_5 gpc2312 (
      {stage1_41[42], stage1_41[43], stage1_41[44], stage1_41[45], stage1_41[46], stage1_41[47]},
      {stage1_43[42], stage1_43[43], stage1_43[44], stage1_43[45], stage1_43[46], stage1_43[47]},
      {stage2_45[7],stage2_44[16],stage2_43[16],stage2_42[19],stage2_41[29]}
   );
   gpc606_5 gpc2313 (
      {stage1_43[48], stage1_43[49], stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[0],stage2_45[8],stage2_44[17],stage2_43[17]}
   );
   gpc606_5 gpc2314 (
      {stage1_43[54], stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[1],stage2_45[9],stage2_44[18],stage2_43[18]}
   );
   gpc606_5 gpc2315 (
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64], stage1_43[65]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[2],stage2_45[10],stage2_44[19],stage2_43[19]}
   );
   gpc606_5 gpc2316 (
      {stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69], stage1_43[70], stage1_43[71]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[3],stage2_45[11],stage2_44[20],stage2_43[20]}
   );
   gpc606_5 gpc2317 (
      {stage1_43[72], stage1_43[73], stage1_43[74], stage1_43[75], stage1_43[76], stage1_43[77]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[4],stage2_45[12],stage2_44[21],stage2_43[21]}
   );
   gpc606_5 gpc2318 (
      {stage1_43[78], stage1_43[79], stage1_43[80], stage1_43[81], stage1_43[82], stage1_43[83]},
      {stage1_45[30], stage1_45[31], stage1_45[32], stage1_45[33], stage1_45[34], stage1_45[35]},
      {stage2_47[5],stage2_46[5],stage2_45[13],stage2_44[22],stage2_43[22]}
   );
   gpc606_5 gpc2319 (
      {stage1_43[84], stage1_43[85], stage1_43[86], stage1_43[87], stage1_43[88], stage1_43[89]},
      {stage1_45[36], stage1_45[37], stage1_45[38], stage1_45[39], stage1_45[40], stage1_45[41]},
      {stage2_47[6],stage2_46[6],stage2_45[14],stage2_44[23],stage2_43[23]}
   );
   gpc606_5 gpc2320 (
      {stage1_43[90], stage1_43[91], stage1_43[92], stage1_43[93], stage1_43[94], stage1_43[95]},
      {stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46], stage1_45[47]},
      {stage2_47[7],stage2_46[7],stage2_45[15],stage2_44[24],stage2_43[24]}
   );
   gpc606_5 gpc2321 (
      {stage1_43[96], stage1_43[97], stage1_43[98], stage1_43[99], stage1_43[100], stage1_43[101]},
      {stage1_45[48], stage1_45[49], stage1_45[50], stage1_45[51], stage1_45[52], stage1_45[53]},
      {stage2_47[8],stage2_46[8],stage2_45[16],stage2_44[25],stage2_43[25]}
   );
   gpc606_5 gpc2322 (
      {stage1_43[102], stage1_43[103], stage1_43[104], stage1_43[105], stage1_43[106], stage1_43[107]},
      {stage1_45[54], stage1_45[55], stage1_45[56], stage1_45[57], stage1_45[58], stage1_45[59]},
      {stage2_47[9],stage2_46[9],stage2_45[17],stage2_44[26],stage2_43[26]}
   );
   gpc606_5 gpc2323 (
      {stage1_43[108], stage1_43[109], stage1_43[110], stage1_43[111], stage1_43[112], stage1_43[113]},
      {stage1_45[60], stage1_45[61], stage1_45[62], stage1_45[63], stage1_45[64], stage1_45[65]},
      {stage2_47[10],stage2_46[10],stage2_45[18],stage2_44[27],stage2_43[27]}
   );
   gpc615_5 gpc2324 (
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4]},
      {stage1_45[66]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[11],stage2_46[11],stage2_45[19],stage2_44[28]}
   );
   gpc615_5 gpc2325 (
      {stage1_44[5], stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9]},
      {stage1_45[67]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[12],stage2_46[12],stage2_45[20],stage2_44[29]}
   );
   gpc606_5 gpc2326 (
      {stage1_45[68], stage1_45[69], stage1_45[70], stage1_45[71], stage1_45[72], stage1_45[73]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[2],stage2_47[13],stage2_46[13],stage2_45[21]}
   );
   gpc606_5 gpc2327 (
      {stage1_45[74], stage1_45[75], stage1_45[76], stage1_45[77], stage1_45[78], stage1_45[79]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[3],stage2_47[14],stage2_46[14],stage2_45[22]}
   );
   gpc606_5 gpc2328 (
      {stage1_45[80], stage1_45[81], stage1_45[82], stage1_45[83], stage1_45[84], stage1_45[85]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[4],stage2_47[15],stage2_46[15],stage2_45[23]}
   );
   gpc606_5 gpc2329 (
      {stage1_45[86], stage1_45[87], stage1_45[88], stage1_45[89], stage1_45[90], stage1_45[91]},
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage2_49[3],stage2_48[5],stage2_47[16],stage2_46[16],stage2_45[24]}
   );
   gpc615_5 gpc2330 (
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16]},
      {stage1_47[24]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[4],stage2_48[6],stage2_47[17],stage2_46[17]}
   );
   gpc615_5 gpc2331 (
      {stage1_46[17], stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21]},
      {stage1_47[25]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[5],stage2_48[7],stage2_47[18],stage2_46[18]}
   );
   gpc615_5 gpc2332 (
      {stage1_46[22], stage1_46[23], stage1_46[24], stage1_46[25], stage1_46[26]},
      {stage1_47[26]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[6],stage2_48[8],stage2_47[19],stage2_46[19]}
   );
   gpc615_5 gpc2333 (
      {stage1_46[27], stage1_46[28], stage1_46[29], stage1_46[30], stage1_46[31]},
      {stage1_47[27]},
      {stage1_48[18], stage1_48[19], stage1_48[20], stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage2_50[3],stage2_49[7],stage2_48[9],stage2_47[20],stage2_46[20]}
   );
   gpc615_5 gpc2334 (
      {stage1_46[32], stage1_46[33], stage1_46[34], stage1_46[35], stage1_46[36]},
      {stage1_47[28]},
      {stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27], stage1_48[28], stage1_48[29]},
      {stage2_50[4],stage2_49[8],stage2_48[10],stage2_47[21],stage2_46[21]}
   );
   gpc615_5 gpc2335 (
      {stage1_46[37], stage1_46[38], stage1_46[39], stage1_46[40], stage1_46[41]},
      {stage1_47[29]},
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage2_50[5],stage2_49[9],stage2_48[11],stage2_47[22],stage2_46[22]}
   );
   gpc615_5 gpc2336 (
      {stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45], stage1_46[46]},
      {stage1_47[30]},
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage2_50[6],stage2_49[10],stage2_48[12],stage2_47[23],stage2_46[23]}
   );
   gpc615_5 gpc2337 (
      {stage1_46[47], stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51]},
      {stage1_47[31]},
      {stage1_48[42], stage1_48[43], stage1_48[44], stage1_48[45], stage1_48[46], stage1_48[47]},
      {stage2_50[7],stage2_49[11],stage2_48[13],stage2_47[24],stage2_46[24]}
   );
   gpc615_5 gpc2338 (
      {stage1_46[52], stage1_46[53], stage1_46[54], stage1_46[55], stage1_46[56]},
      {stage1_47[32]},
      {stage1_48[48], stage1_48[49], stage1_48[50], stage1_48[51], stage1_48[52], stage1_48[53]},
      {stage2_50[8],stage2_49[12],stage2_48[14],stage2_47[25],stage2_46[25]}
   );
   gpc606_5 gpc2339 (
      {stage1_47[33], stage1_47[34], stage1_47[35], stage1_47[36], stage1_47[37], stage1_47[38]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[9],stage2_49[13],stage2_48[15],stage2_47[26]}
   );
   gpc606_5 gpc2340 (
      {stage1_48[54], stage1_48[55], stage1_48[56], stage1_48[57], stage1_48[58], stage1_48[59]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[1],stage2_50[10],stage2_49[14],stage2_48[16]}
   );
   gpc606_5 gpc2341 (
      {stage1_48[60], stage1_48[61], stage1_48[62], stage1_48[63], stage1_48[64], stage1_48[65]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[1],stage2_51[2],stage2_50[11],stage2_49[15],stage2_48[17]}
   );
   gpc606_5 gpc2342 (
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[2],stage2_51[3],stage2_50[12],stage2_49[16]}
   );
   gpc606_5 gpc2343 (
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage2_53[1],stage2_52[3],stage2_51[4],stage2_50[13],stage2_49[17]}
   );
   gpc606_5 gpc2344 (
      {stage1_49[18], stage1_49[19], stage1_49[20], stage1_49[21], stage1_49[22], stage1_49[23]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage2_53[2],stage2_52[4],stage2_51[5],stage2_50[14],stage2_49[18]}
   );
   gpc606_5 gpc2345 (
      {stage1_49[24], stage1_49[25], stage1_49[26], stage1_49[27], stage1_49[28], stage1_49[29]},
      {stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21], stage1_51[22], stage1_51[23]},
      {stage2_53[3],stage2_52[5],stage2_51[6],stage2_50[15],stage2_49[19]}
   );
   gpc606_5 gpc2346 (
      {stage1_49[30], stage1_49[31], stage1_49[32], stage1_49[33], stage1_49[34], stage1_49[35]},
      {stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27], stage1_51[28], stage1_51[29]},
      {stage2_53[4],stage2_52[6],stage2_51[7],stage2_50[16],stage2_49[20]}
   );
   gpc606_5 gpc2347 (
      {stage1_49[36], stage1_49[37], stage1_49[38], stage1_49[39], stage1_49[40], stage1_49[41]},
      {stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33], stage1_51[34], stage1_51[35]},
      {stage2_53[5],stage2_52[7],stage2_51[8],stage2_50[17],stage2_49[21]}
   );
   gpc606_5 gpc2348 (
      {stage1_49[42], stage1_49[43], stage1_49[44], stage1_49[45], stage1_49[46], stage1_49[47]},
      {stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39], stage1_51[40], stage1_51[41]},
      {stage2_53[6],stage2_52[8],stage2_51[9],stage2_50[18],stage2_49[22]}
   );
   gpc606_5 gpc2349 (
      {stage1_49[48], stage1_49[49], stage1_49[50], stage1_49[51], stage1_49[52], stage1_49[53]},
      {stage1_51[42], stage1_51[43], stage1_51[44], stage1_51[45], stage1_51[46], stage1_51[47]},
      {stage2_53[7],stage2_52[9],stage2_51[10],stage2_50[19],stage2_49[23]}
   );
   gpc606_5 gpc2350 (
      {stage1_49[54], stage1_49[55], stage1_49[56], stage1_49[57], stage1_49[58], stage1_49[59]},
      {stage1_51[48], stage1_51[49], stage1_51[50], stage1_51[51], stage1_51[52], stage1_51[53]},
      {stage2_53[8],stage2_52[10],stage2_51[11],stage2_50[20],stage2_49[24]}
   );
   gpc606_5 gpc2351 (
      {stage1_49[60], stage1_49[61], stage1_49[62], stage1_49[63], stage1_49[64], stage1_49[65]},
      {stage1_51[54], stage1_51[55], stage1_51[56], stage1_51[57], stage1_51[58], stage1_51[59]},
      {stage2_53[9],stage2_52[11],stage2_51[12],stage2_50[21],stage2_49[25]}
   );
   gpc606_5 gpc2352 (
      {stage1_49[66], stage1_49[67], stage1_49[68], stage1_49[69], stage1_49[70], stage1_49[71]},
      {stage1_51[60], stage1_51[61], stage1_51[62], stage1_51[63], stage1_51[64], stage1_51[65]},
      {stage2_53[10],stage2_52[12],stage2_51[13],stage2_50[22],stage2_49[26]}
   );
   gpc606_5 gpc2353 (
      {stage1_49[72], stage1_49[73], stage1_49[74], stage1_49[75], stage1_49[76], stage1_49[77]},
      {stage1_51[66], stage1_51[67], stage1_51[68], stage1_51[69], stage1_51[70], stage1_51[71]},
      {stage2_53[11],stage2_52[13],stage2_51[14],stage2_50[23],stage2_49[27]}
   );
   gpc117_4 gpc2354 (
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16], stage1_50[17], stage1_50[18]},
      {stage1_51[72]},
      {stage1_52[0]},
      {stage2_53[12],stage2_52[14],stage2_51[15],stage2_50[24]}
   );
   gpc606_5 gpc2355 (
      {stage1_50[19], stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23], stage1_50[24]},
      {stage1_52[1], stage1_52[2], stage1_52[3], stage1_52[4], stage1_52[5], stage1_52[6]},
      {stage2_54[0],stage2_53[13],stage2_52[15],stage2_51[16],stage2_50[25]}
   );
   gpc606_5 gpc2356 (
      {stage1_50[25], stage1_50[26], stage1_50[27], stage1_50[28], stage1_50[29], stage1_50[30]},
      {stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10], stage1_52[11], stage1_52[12]},
      {stage2_54[1],stage2_53[14],stage2_52[16],stage2_51[17],stage2_50[26]}
   );
   gpc606_5 gpc2357 (
      {stage1_50[31], stage1_50[32], stage1_50[33], stage1_50[34], stage1_50[35], stage1_50[36]},
      {stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16], stage1_52[17], stage1_52[18]},
      {stage2_54[2],stage2_53[15],stage2_52[17],stage2_51[18],stage2_50[27]}
   );
   gpc615_5 gpc2358 (
      {stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40], stage1_50[41]},
      {stage1_51[73]},
      {stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22], stage1_52[23], stage1_52[24]},
      {stage2_54[3],stage2_53[16],stage2_52[18],stage2_51[19],stage2_50[28]}
   );
   gpc615_5 gpc2359 (
      {stage1_50[42], stage1_50[43], stage1_50[44], stage1_50[45], stage1_50[46]},
      {stage1_51[74]},
      {stage1_52[25], stage1_52[26], stage1_52[27], stage1_52[28], stage1_52[29], stage1_52[30]},
      {stage2_54[4],stage2_53[17],stage2_52[19],stage2_51[20],stage2_50[29]}
   );
   gpc606_5 gpc2360 (
      {stage1_51[75], stage1_51[76], stage1_51[77], stage1_51[78], stage1_51[79], stage1_51[80]},
      {stage1_53[0], stage1_53[1], stage1_53[2], stage1_53[3], stage1_53[4], stage1_53[5]},
      {stage2_55[0],stage2_54[5],stage2_53[18],stage2_52[20],stage2_51[21]}
   );
   gpc606_5 gpc2361 (
      {stage1_51[81], stage1_51[82], stage1_51[83], stage1_51[84], stage1_51[85], stage1_51[86]},
      {stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9], stage1_53[10], stage1_53[11]},
      {stage2_55[1],stage2_54[6],stage2_53[19],stage2_52[21],stage2_51[22]}
   );
   gpc606_5 gpc2362 (
      {stage1_51[87], stage1_51[88], stage1_51[89], stage1_51[90], stage1_51[91], stage1_51[92]},
      {stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15], stage1_53[16], stage1_53[17]},
      {stage2_55[2],stage2_54[7],stage2_53[20],stage2_52[22],stage2_51[23]}
   );
   gpc606_5 gpc2363 (
      {stage1_52[31], stage1_52[32], stage1_52[33], stage1_52[34], stage1_52[35], stage1_52[36]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[3],stage2_54[8],stage2_53[21],stage2_52[23]}
   );
   gpc606_5 gpc2364 (
      {stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41], stage1_52[42]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[4],stage2_54[9],stage2_53[22],stage2_52[24]}
   );
   gpc606_5 gpc2365 (
      {stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46], stage1_52[47], stage1_52[48]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[5],stage2_54[10],stage2_53[23],stage2_52[25]}
   );
   gpc606_5 gpc2366 (
      {stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52], stage1_52[53], stage1_52[54]},
      {stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21], stage1_54[22], stage1_54[23]},
      {stage2_56[3],stage2_55[6],stage2_54[11],stage2_53[24],stage2_52[26]}
   );
   gpc606_5 gpc2367 (
      {stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58], stage1_52[59], stage1_52[60]},
      {stage1_54[24], stage1_54[25], stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29]},
      {stage2_56[4],stage2_55[7],stage2_54[12],stage2_53[25],stage2_52[27]}
   );
   gpc606_5 gpc2368 (
      {stage1_52[61], stage1_52[62], stage1_52[63], stage1_52[64], stage1_52[65], stage1_52[66]},
      {stage1_54[30], stage1_54[31], stage1_54[32], stage1_54[33], stage1_54[34], stage1_54[35]},
      {stage2_56[5],stage2_55[8],stage2_54[13],stage2_53[26],stage2_52[28]}
   );
   gpc606_5 gpc2369 (
      {stage1_52[67], stage1_52[68], stage1_52[69], stage1_52[70], stage1_52[71], stage1_52[72]},
      {stage1_54[36], stage1_54[37], stage1_54[38], stage1_54[39], stage1_54[40], stage1_54[41]},
      {stage2_56[6],stage2_55[9],stage2_54[14],stage2_53[27],stage2_52[29]}
   );
   gpc606_5 gpc2370 (
      {stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21], stage1_53[22], stage1_53[23]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[7],stage2_55[10],stage2_54[15],stage2_53[28]}
   );
   gpc606_5 gpc2371 (
      {stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28], stage1_53[29]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage2_57[1],stage2_56[8],stage2_55[11],stage2_54[16],stage2_53[29]}
   );
   gpc606_5 gpc2372 (
      {stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34], stage1_53[35]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage2_57[2],stage2_56[9],stage2_55[12],stage2_54[17],stage2_53[30]}
   );
   gpc606_5 gpc2373 (
      {stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39], stage1_53[40], stage1_53[41]},
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22], stage1_55[23]},
      {stage2_57[3],stage2_56[10],stage2_55[13],stage2_54[18],stage2_53[31]}
   );
   gpc606_5 gpc2374 (
      {stage1_53[42], stage1_53[43], stage1_53[44], stage1_53[45], stage1_53[46], stage1_53[47]},
      {stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27], stage1_55[28], stage1_55[29]},
      {stage2_57[4],stage2_56[11],stage2_55[14],stage2_54[19],stage2_53[32]}
   );
   gpc615_5 gpc2375 (
      {stage1_54[42], stage1_54[43], stage1_54[44], stage1_54[45], stage1_54[46]},
      {stage1_55[30]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[5],stage2_56[12],stage2_55[15],stage2_54[20]}
   );
   gpc615_5 gpc2376 (
      {stage1_54[47], stage1_54[48], stage1_54[49], stage1_54[50], stage1_54[51]},
      {stage1_55[31]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[6],stage2_56[13],stage2_55[16],stage2_54[21]}
   );
   gpc606_5 gpc2377 (
      {stage1_55[32], stage1_55[33], stage1_55[34], stage1_55[35], stage1_55[36], stage1_55[37]},
      {stage1_57[0], stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage2_59[0],stage2_58[2],stage2_57[7],stage2_56[14],stage2_55[17]}
   );
   gpc615_5 gpc2378 (
      {stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41], stage1_55[42]},
      {stage1_56[12]},
      {stage1_57[6], stage1_57[7], stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11]},
      {stage2_59[1],stage2_58[3],stage2_57[8],stage2_56[15],stage2_55[18]}
   );
   gpc615_5 gpc2379 (
      {stage1_55[43], stage1_55[44], stage1_55[45], stage1_55[46], stage1_55[47]},
      {stage1_56[13]},
      {stage1_57[12], stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage2_59[2],stage2_58[4],stage2_57[9],stage2_56[16],stage2_55[19]}
   );
   gpc615_5 gpc2380 (
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52]},
      {stage1_56[14]},
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage2_59[3],stage2_58[5],stage2_57[10],stage2_56[17],stage2_55[20]}
   );
   gpc615_5 gpc2381 (
      {stage1_55[53], stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57]},
      {stage1_56[15]},
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage2_59[4],stage2_58[6],stage2_57[11],stage2_56[18],stage2_55[21]}
   );
   gpc615_5 gpc2382 (
      {stage1_55[58], stage1_55[59], stage1_55[60], stage1_55[61], stage1_55[62]},
      {stage1_56[16]},
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage2_59[5],stage2_58[7],stage2_57[12],stage2_56[19],stage2_55[22]}
   );
   gpc615_5 gpc2383 (
      {stage1_55[63], stage1_55[64], stage1_55[65], stage1_55[66], stage1_55[67]},
      {stage1_56[17]},
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage2_59[6],stage2_58[8],stage2_57[13],stage2_56[20],stage2_55[23]}
   );
   gpc615_5 gpc2384 (
      {stage1_55[68], stage1_55[69], stage1_55[70], stage1_55[71], stage1_55[72]},
      {stage1_56[18]},
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage2_59[7],stage2_58[9],stage2_57[14],stage2_56[21],stage2_55[24]}
   );
   gpc615_5 gpc2385 (
      {stage1_55[73], stage1_55[74], stage1_55[75], stage1_55[76], stage1_55[77]},
      {stage1_56[19]},
      {stage1_57[48], stage1_57[49], stage1_57[50], stage1_57[51], stage1_57[52], stage1_57[53]},
      {stage2_59[8],stage2_58[10],stage2_57[15],stage2_56[22],stage2_55[25]}
   );
   gpc615_5 gpc2386 (
      {stage1_55[78], stage1_55[79], stage1_55[80], stage1_55[81], stage1_55[82]},
      {stage1_56[20]},
      {stage1_57[54], stage1_57[55], stage1_57[56], stage1_57[57], stage1_57[58], stage1_57[59]},
      {stage2_59[9],stage2_58[11],stage2_57[16],stage2_56[23],stage2_55[26]}
   );
   gpc615_5 gpc2387 (
      {stage1_55[83], stage1_55[84], stage1_55[85], stage1_55[86], stage1_55[87]},
      {stage1_56[21]},
      {stage1_57[60], stage1_57[61], stage1_57[62], stage1_57[63], stage1_57[64], stage1_57[65]},
      {stage2_59[10],stage2_58[12],stage2_57[17],stage2_56[24],stage2_55[27]}
   );
   gpc606_5 gpc2388 (
      {stage1_56[22], stage1_56[23], stage1_56[24], stage1_56[25], stage1_56[26], stage1_56[27]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[11],stage2_58[13],stage2_57[18],stage2_56[25]}
   );
   gpc606_5 gpc2389 (
      {stage1_56[28], stage1_56[29], stage1_56[30], stage1_56[31], stage1_56[32], stage1_56[33]},
      {stage1_58[6], stage1_58[7], stage1_58[8], stage1_58[9], stage1_58[10], stage1_58[11]},
      {stage2_60[1],stage2_59[12],stage2_58[14],stage2_57[19],stage2_56[26]}
   );
   gpc606_5 gpc2390 (
      {stage1_56[34], stage1_56[35], stage1_56[36], stage1_56[37], stage1_56[38], stage1_56[39]},
      {stage1_58[12], stage1_58[13], stage1_58[14], stage1_58[15], stage1_58[16], stage1_58[17]},
      {stage2_60[2],stage2_59[13],stage2_58[15],stage2_57[20],stage2_56[27]}
   );
   gpc606_5 gpc2391 (
      {stage1_56[40], stage1_56[41], stage1_56[42], stage1_56[43], stage1_56[44], stage1_56[45]},
      {stage1_58[18], stage1_58[19], stage1_58[20], stage1_58[21], stage1_58[22], stage1_58[23]},
      {stage2_60[3],stage2_59[14],stage2_58[16],stage2_57[21],stage2_56[28]}
   );
   gpc606_5 gpc2392 (
      {stage1_56[46], stage1_56[47], stage1_56[48], stage1_56[49], stage1_56[50], stage1_56[51]},
      {stage1_58[24], stage1_58[25], stage1_58[26], stage1_58[27], stage1_58[28], stage1_58[29]},
      {stage2_60[4],stage2_59[15],stage2_58[17],stage2_57[22],stage2_56[29]}
   );
   gpc606_5 gpc2393 (
      {stage1_56[52], stage1_56[53], stage1_56[54], stage1_56[55], stage1_56[56], stage1_56[57]},
      {stage1_58[30], stage1_58[31], stage1_58[32], stage1_58[33], stage1_58[34], stage1_58[35]},
      {stage2_60[5],stage2_59[16],stage2_58[18],stage2_57[23],stage2_56[30]}
   );
   gpc606_5 gpc2394 (
      {stage1_58[36], stage1_58[37], stage1_58[38], stage1_58[39], stage1_58[40], stage1_58[41]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[0],stage2_60[6],stage2_59[17],stage2_58[19]}
   );
   gpc606_5 gpc2395 (
      {stage1_58[42], stage1_58[43], stage1_58[44], stage1_58[45], stage1_58[46], stage1_58[47]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[1],stage2_60[7],stage2_59[18],stage2_58[20]}
   );
   gpc606_5 gpc2396 (
      {stage1_58[48], stage1_58[49], stage1_58[50], stage1_58[51], stage1_58[52], stage1_58[53]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[2],stage2_60[8],stage2_59[19],stage2_58[21]}
   );
   gpc606_5 gpc2397 (
      {stage1_58[54], stage1_58[55], stage1_58[56], stage1_58[57], stage1_58[58], stage1_58[59]},
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22], stage1_60[23]},
      {stage2_62[3],stage2_61[3],stage2_60[9],stage2_59[20],stage2_58[22]}
   );
   gpc615_5 gpc2398 (
      {stage1_58[60], stage1_58[61], stage1_58[62], stage1_58[63], stage1_58[64]},
      {stage1_59[0]},
      {stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27], stage1_60[28], stage1_60[29]},
      {stage2_62[4],stage2_61[4],stage2_60[10],stage2_59[21],stage2_58[23]}
   );
   gpc606_5 gpc2399 (
      {stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5], stage1_59[6]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[5],stage2_61[5],stage2_60[11],stage2_59[22]}
   );
   gpc606_5 gpc2400 (
      {stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11], stage1_59[12]},
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage2_63[1],stage2_62[6],stage2_61[6],stage2_60[12],stage2_59[23]}
   );
   gpc606_5 gpc2401 (
      {stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17], stage1_59[18]},
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage2_63[2],stage2_62[7],stage2_61[7],stage2_60[13],stage2_59[24]}
   );
   gpc606_5 gpc2402 (
      {stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23], stage1_59[24]},
      {stage1_61[18], stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23]},
      {stage2_63[3],stage2_62[8],stage2_61[8],stage2_60[14],stage2_59[25]}
   );
   gpc606_5 gpc2403 (
      {stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33], stage1_60[34], stage1_60[35]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage2_64[0],stage2_63[4],stage2_62[9],stage2_61[9],stage2_60[15]}
   );
   gpc606_5 gpc2404 (
      {stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39], stage1_60[40], stage1_60[41]},
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage2_64[1],stage2_63[5],stage2_62[10],stage2_61[10],stage2_60[16]}
   );
   gpc606_5 gpc2405 (
      {stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45], stage1_60[46], stage1_60[47]},
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage2_64[2],stage2_63[6],stage2_62[11],stage2_61[11],stage2_60[17]}
   );
   gpc606_5 gpc2406 (
      {stage1_60[48], stage1_60[49], stage1_60[50], stage1_60[51], stage1_60[52], stage1_60[53]},
      {stage1_62[18], stage1_62[19], stage1_62[20], stage1_62[21], stage1_62[22], stage1_62[23]},
      {stage2_64[3],stage2_63[7],stage2_62[12],stage2_61[12],stage2_60[18]}
   );
   gpc606_5 gpc2407 (
      {stage1_60[54], stage1_60[55], stage1_60[56], stage1_60[57], stage1_60[58], stage1_60[59]},
      {stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29]},
      {stage2_64[4],stage2_63[8],stage2_62[13],stage2_61[13],stage2_60[19]}
   );
   gpc606_5 gpc2408 (
      {stage1_60[60], stage1_60[61], stage1_60[62], stage1_60[63], stage1_60[64], stage1_60[65]},
      {stage1_62[30], stage1_62[31], stage1_62[32], stage1_62[33], stage1_62[34], stage1_62[35]},
      {stage2_64[5],stage2_63[9],stage2_62[14],stage2_61[14],stage2_60[20]}
   );
   gpc606_5 gpc2409 (
      {stage1_61[24], stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[6],stage2_63[10],stage2_62[15],stage2_61[15]}
   );
   gpc606_5 gpc2410 (
      {stage1_61[30], stage1_61[31], stage1_61[32], stage1_61[33], stage1_61[34], stage1_61[35]},
      {stage1_63[6], stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11]},
      {stage2_65[1],stage2_64[7],stage2_63[11],stage2_62[16],stage2_61[16]}
   );
   gpc606_5 gpc2411 (
      {stage1_61[36], stage1_61[37], stage1_61[38], stage1_61[39], stage1_61[40], stage1_61[41]},
      {stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17]},
      {stage2_65[2],stage2_64[8],stage2_63[12],stage2_62[17],stage2_61[17]}
   );
   gpc2135_5 gpc2412 (
      {stage1_62[36], stage1_62[37], stage1_62[38], stage1_62[39], stage1_62[40]},
      {stage1_63[18], stage1_63[19], stage1_63[20]},
      {stage1_64[0]},
      {stage1_65[0], stage1_65[1]},
      {stage2_66[0],stage2_65[3],stage2_64[9],stage2_63[13],stage2_62[18]}
   );
   gpc2135_5 gpc2413 (
      {stage1_62[41], stage1_62[42], stage1_62[43], stage1_62[44], stage1_62[45]},
      {stage1_63[21], stage1_63[22], stage1_63[23]},
      {stage1_64[1]},
      {stage1_65[2], stage1_65[3]},
      {stage2_66[1],stage2_65[4],stage2_64[10],stage2_63[14],stage2_62[19]}
   );
   gpc2135_5 gpc2414 (
      {stage1_62[46], stage1_62[47], stage1_62[48], stage1_62[49], stage1_62[50]},
      {stage1_63[24], stage1_63[25], stage1_63[26]},
      {stage1_64[2]},
      {stage1_65[4], stage1_65[5]},
      {stage2_66[2],stage2_65[5],stage2_64[11],stage2_63[15],stage2_62[20]}
   );
   gpc2135_5 gpc2415 (
      {stage1_62[51], stage1_62[52], stage1_62[53], stage1_62[54], stage1_62[55]},
      {stage1_63[27], stage1_63[28], stage1_63[29]},
      {stage1_64[3]},
      {stage1_65[6], stage1_65[7]},
      {stage2_66[3],stage2_65[6],stage2_64[12],stage2_63[16],stage2_62[21]}
   );
   gpc2135_5 gpc2416 (
      {stage1_62[56], stage1_62[57], stage1_62[58], stage1_62[59], stage1_62[60]},
      {stage1_63[30], stage1_63[31], stage1_63[32]},
      {stage1_64[4]},
      {stage1_65[8], stage1_65[9]},
      {stage2_66[4],stage2_65[7],stage2_64[13],stage2_63[17],stage2_62[22]}
   );
   gpc2135_5 gpc2417 (
      {stage1_62[61], stage1_62[62], stage1_62[63], stage1_62[64], stage1_62[65]},
      {stage1_63[33], stage1_63[34], stage1_63[35]},
      {stage1_64[5]},
      {stage1_65[10], stage1_65[11]},
      {stage2_66[5],stage2_65[8],stage2_64[14],stage2_63[18],stage2_62[23]}
   );
   gpc606_5 gpc2418 (
      {stage1_62[66], stage1_62[67], stage1_62[68], stage1_62[69], stage1_62[70], stage1_62[71]},
      {stage1_64[6], stage1_64[7], stage1_64[8], stage1_64[9], stage1_64[10], stage1_64[11]},
      {stage2_66[6],stage2_65[9],stage2_64[15],stage2_63[19],stage2_62[24]}
   );
   gpc606_5 gpc2419 (
      {stage1_62[72], stage1_62[73], stage1_62[74], stage1_62[75], stage1_62[76], stage1_62[77]},
      {stage1_64[12], stage1_64[13], stage1_64[14], stage1_64[15], stage1_64[16], stage1_64[17]},
      {stage2_66[7],stage2_65[10],stage2_64[16],stage2_63[20],stage2_62[25]}
   );
   gpc606_5 gpc2420 (
      {stage1_63[36], stage1_63[37], stage1_63[38], stage1_63[39], stage1_63[40], stage1_63[41]},
      {stage1_65[12], stage1_65[13], stage1_65[14], stage1_65[15], stage1_65[16], stage1_65[17]},
      {stage2_67[0],stage2_66[8],stage2_65[11],stage2_64[17],stage2_63[21]}
   );
   gpc606_5 gpc2421 (
      {stage1_63[42], stage1_63[43], stage1_63[44], stage1_63[45], stage1_63[46], stage1_63[47]},
      {stage1_65[18], stage1_65[19], stage1_65[20], stage1_65[21], stage1_65[22], stage1_65[23]},
      {stage2_67[1],stage2_66[9],stage2_65[12],stage2_64[18],stage2_63[22]}
   );
   gpc1_1 gpc2422 (
      {stage1_0[31]},
      {stage2_0[7]}
   );
   gpc1_1 gpc2423 (
      {stage1_0[32]},
      {stage2_0[8]}
   );
   gpc1_1 gpc2424 (
      {stage1_0[33]},
      {stage2_0[9]}
   );
   gpc1_1 gpc2425 (
      {stage1_1[38]},
      {stage2_1[10]}
   );
   gpc1_1 gpc2426 (
      {stage1_1[39]},
      {stage2_1[11]}
   );
   gpc1_1 gpc2427 (
      {stage1_1[40]},
      {stage2_1[12]}
   );
   gpc1_1 gpc2428 (
      {stage1_1[41]},
      {stage2_1[13]}
   );
   gpc1_1 gpc2429 (
      {stage1_1[42]},
      {stage2_1[14]}
   );
   gpc1_1 gpc2430 (
      {stage1_1[43]},
      {stage2_1[15]}
   );
   gpc1_1 gpc2431 (
      {stage1_1[44]},
      {stage2_1[16]}
   );
   gpc1_1 gpc2432 (
      {stage1_1[45]},
      {stage2_1[17]}
   );
   gpc1_1 gpc2433 (
      {stage1_1[46]},
      {stage2_1[18]}
   );
   gpc1_1 gpc2434 (
      {stage1_2[27]},
      {stage2_2[10]}
   );
   gpc1_1 gpc2435 (
      {stage1_2[28]},
      {stage2_2[11]}
   );
   gpc1_1 gpc2436 (
      {stage1_2[29]},
      {stage2_2[12]}
   );
   gpc1_1 gpc2437 (
      {stage1_2[30]},
      {stage2_2[13]}
   );
   gpc1_1 gpc2438 (
      {stage1_2[31]},
      {stage2_2[14]}
   );
   gpc1_1 gpc2439 (
      {stage1_2[32]},
      {stage2_2[15]}
   );
   gpc1_1 gpc2440 (
      {stage1_2[33]},
      {stage2_2[16]}
   );
   gpc1_1 gpc2441 (
      {stage1_2[34]},
      {stage2_2[17]}
   );
   gpc1_1 gpc2442 (
      {stage1_2[35]},
      {stage2_2[18]}
   );
   gpc1_1 gpc2443 (
      {stage1_2[36]},
      {stage2_2[19]}
   );
   gpc1_1 gpc2444 (
      {stage1_2[37]},
      {stage2_2[20]}
   );
   gpc1_1 gpc2445 (
      {stage1_2[38]},
      {stage2_2[21]}
   );
   gpc1_1 gpc2446 (
      {stage1_2[39]},
      {stage2_2[22]}
   );
   gpc1_1 gpc2447 (
      {stage1_2[40]},
      {stage2_2[23]}
   );
   gpc1_1 gpc2448 (
      {stage1_2[41]},
      {stage2_2[24]}
   );
   gpc1_1 gpc2449 (
      {stage1_2[42]},
      {stage2_2[25]}
   );
   gpc1_1 gpc2450 (
      {stage1_2[43]},
      {stage2_2[26]}
   );
   gpc1_1 gpc2451 (
      {stage1_2[44]},
      {stage2_2[27]}
   );
   gpc1_1 gpc2452 (
      {stage1_2[45]},
      {stage2_2[28]}
   );
   gpc1_1 gpc2453 (
      {stage1_2[46]},
      {stage2_2[29]}
   );
   gpc1_1 gpc2454 (
      {stage1_2[47]},
      {stage2_2[30]}
   );
   gpc1_1 gpc2455 (
      {stage1_2[48]},
      {stage2_2[31]}
   );
   gpc1_1 gpc2456 (
      {stage1_2[49]},
      {stage2_2[32]}
   );
   gpc1_1 gpc2457 (
      {stage1_2[50]},
      {stage2_2[33]}
   );
   gpc1_1 gpc2458 (
      {stage1_2[51]},
      {stage2_2[34]}
   );
   gpc1_1 gpc2459 (
      {stage1_2[52]},
      {stage2_2[35]}
   );
   gpc1_1 gpc2460 (
      {stage1_2[53]},
      {stage2_2[36]}
   );
   gpc1_1 gpc2461 (
      {stage1_2[54]},
      {stage2_2[37]}
   );
   gpc1_1 gpc2462 (
      {stage1_4[66]},
      {stage2_4[31]}
   );
   gpc1_1 gpc2463 (
      {stage1_4[67]},
      {stage2_4[32]}
   );
   gpc1_1 gpc2464 (
      {stage1_4[68]},
      {stage2_4[33]}
   );
   gpc1_1 gpc2465 (
      {stage1_4[69]},
      {stage2_4[34]}
   );
   gpc1_1 gpc2466 (
      {stage1_4[70]},
      {stage2_4[35]}
   );
   gpc1_1 gpc2467 (
      {stage1_4[71]},
      {stage2_4[36]}
   );
   gpc1_1 gpc2468 (
      {stage1_4[72]},
      {stage2_4[37]}
   );
   gpc1_1 gpc2469 (
      {stage1_4[73]},
      {stage2_4[38]}
   );
   gpc1_1 gpc2470 (
      {stage1_4[74]},
      {stage2_4[39]}
   );
   gpc1_1 gpc2471 (
      {stage1_4[75]},
      {stage2_4[40]}
   );
   gpc1_1 gpc2472 (
      {stage1_4[76]},
      {stage2_4[41]}
   );
   gpc1_1 gpc2473 (
      {stage1_4[77]},
      {stage2_4[42]}
   );
   gpc1_1 gpc2474 (
      {stage1_4[78]},
      {stage2_4[43]}
   );
   gpc1_1 gpc2475 (
      {stage1_4[79]},
      {stage2_4[44]}
   );
   gpc1_1 gpc2476 (
      {stage1_4[80]},
      {stage2_4[45]}
   );
   gpc1_1 gpc2477 (
      {stage1_4[81]},
      {stage2_4[46]}
   );
   gpc1_1 gpc2478 (
      {stage1_4[82]},
      {stage2_4[47]}
   );
   gpc1_1 gpc2479 (
      {stage1_5[109]},
      {stage2_5[30]}
   );
   gpc1_1 gpc2480 (
      {stage1_5[110]},
      {stage2_5[31]}
   );
   gpc1_1 gpc2481 (
      {stage1_5[111]},
      {stage2_5[32]}
   );
   gpc1_1 gpc2482 (
      {stage1_5[112]},
      {stage2_5[33]}
   );
   gpc1_1 gpc2483 (
      {stage1_5[113]},
      {stage2_5[34]}
   );
   gpc1_1 gpc2484 (
      {stage1_5[114]},
      {stage2_5[35]}
   );
   gpc1_1 gpc2485 (
      {stage1_7[64]},
      {stage2_7[34]}
   );
   gpc1_1 gpc2486 (
      {stage1_7[65]},
      {stage2_7[35]}
   );
   gpc1_1 gpc2487 (
      {stage1_7[66]},
      {stage2_7[36]}
   );
   gpc1_1 gpc2488 (
      {stage1_7[67]},
      {stage2_7[37]}
   );
   gpc1_1 gpc2489 (
      {stage1_7[68]},
      {stage2_7[38]}
   );
   gpc1_1 gpc2490 (
      {stage1_7[69]},
      {stage2_7[39]}
   );
   gpc1_1 gpc2491 (
      {stage1_7[70]},
      {stage2_7[40]}
   );
   gpc1_1 gpc2492 (
      {stage1_8[46]},
      {stage2_8[26]}
   );
   gpc1_1 gpc2493 (
      {stage1_8[47]},
      {stage2_8[27]}
   );
   gpc1_1 gpc2494 (
      {stage1_8[48]},
      {stage2_8[28]}
   );
   gpc1_1 gpc2495 (
      {stage1_8[49]},
      {stage2_8[29]}
   );
   gpc1_1 gpc2496 (
      {stage1_8[50]},
      {stage2_8[30]}
   );
   gpc1_1 gpc2497 (
      {stage1_8[51]},
      {stage2_8[31]}
   );
   gpc1_1 gpc2498 (
      {stage1_8[52]},
      {stage2_8[32]}
   );
   gpc1_1 gpc2499 (
      {stage1_8[53]},
      {stage2_8[33]}
   );
   gpc1_1 gpc2500 (
      {stage1_8[54]},
      {stage2_8[34]}
   );
   gpc1_1 gpc2501 (
      {stage1_8[55]},
      {stage2_8[35]}
   );
   gpc1_1 gpc2502 (
      {stage1_8[56]},
      {stage2_8[36]}
   );
   gpc1_1 gpc2503 (
      {stage1_8[57]},
      {stage2_8[37]}
   );
   gpc1_1 gpc2504 (
      {stage1_8[58]},
      {stage2_8[38]}
   );
   gpc1_1 gpc2505 (
      {stage1_8[59]},
      {stage2_8[39]}
   );
   gpc1_1 gpc2506 (
      {stage1_8[60]},
      {stage2_8[40]}
   );
   gpc1_1 gpc2507 (
      {stage1_8[61]},
      {stage2_8[41]}
   );
   gpc1_1 gpc2508 (
      {stage1_8[62]},
      {stage2_8[42]}
   );
   gpc1_1 gpc2509 (
      {stage1_8[63]},
      {stage2_8[43]}
   );
   gpc1_1 gpc2510 (
      {stage1_8[64]},
      {stage2_8[44]}
   );
   gpc1_1 gpc2511 (
      {stage1_8[65]},
      {stage2_8[45]}
   );
   gpc1_1 gpc2512 (
      {stage1_8[66]},
      {stage2_8[46]}
   );
   gpc1_1 gpc2513 (
      {stage1_8[67]},
      {stage2_8[47]}
   );
   gpc1_1 gpc2514 (
      {stage1_8[68]},
      {stage2_8[48]}
   );
   gpc1_1 gpc2515 (
      {stage1_8[69]},
      {stage2_8[49]}
   );
   gpc1_1 gpc2516 (
      {stage1_8[70]},
      {stage2_8[50]}
   );
   gpc1_1 gpc2517 (
      {stage1_8[71]},
      {stage2_8[51]}
   );
   gpc1_1 gpc2518 (
      {stage1_8[72]},
      {stage2_8[52]}
   );
   gpc1_1 gpc2519 (
      {stage1_8[73]},
      {stage2_8[53]}
   );
   gpc1_1 gpc2520 (
      {stage1_8[74]},
      {stage2_8[54]}
   );
   gpc1_1 gpc2521 (
      {stage1_8[75]},
      {stage2_8[55]}
   );
   gpc1_1 gpc2522 (
      {stage1_8[76]},
      {stage2_8[56]}
   );
   gpc1_1 gpc2523 (
      {stage1_8[77]},
      {stage2_8[57]}
   );
   gpc1_1 gpc2524 (
      {stage1_8[78]},
      {stage2_8[58]}
   );
   gpc1_1 gpc2525 (
      {stage1_8[79]},
      {stage2_8[59]}
   );
   gpc1_1 gpc2526 (
      {stage1_8[80]},
      {stage2_8[60]}
   );
   gpc1_1 gpc2527 (
      {stage1_9[54]},
      {stage2_9[22]}
   );
   gpc1_1 gpc2528 (
      {stage1_9[55]},
      {stage2_9[23]}
   );
   gpc1_1 gpc2529 (
      {stage1_9[56]},
      {stage2_9[24]}
   );
   gpc1_1 gpc2530 (
      {stage1_9[57]},
      {stage2_9[25]}
   );
   gpc1_1 gpc2531 (
      {stage1_10[79]},
      {stage2_10[25]}
   );
   gpc1_1 gpc2532 (
      {stage1_10[80]},
      {stage2_10[26]}
   );
   gpc1_1 gpc2533 (
      {stage1_10[81]},
      {stage2_10[27]}
   );
   gpc1_1 gpc2534 (
      {stage1_10[82]},
      {stage2_10[28]}
   );
   gpc1_1 gpc2535 (
      {stage1_10[83]},
      {stage2_10[29]}
   );
   gpc1_1 gpc2536 (
      {stage1_10[84]},
      {stage2_10[30]}
   );
   gpc1_1 gpc2537 (
      {stage1_10[85]},
      {stage2_10[31]}
   );
   gpc1_1 gpc2538 (
      {stage1_10[86]},
      {stage2_10[32]}
   );
   gpc1_1 gpc2539 (
      {stage1_10[87]},
      {stage2_10[33]}
   );
   gpc1_1 gpc2540 (
      {stage1_10[88]},
      {stage2_10[34]}
   );
   gpc1_1 gpc2541 (
      {stage1_10[89]},
      {stage2_10[35]}
   );
   gpc1_1 gpc2542 (
      {stage1_10[90]},
      {stage2_10[36]}
   );
   gpc1_1 gpc2543 (
      {stage1_10[91]},
      {stage2_10[37]}
   );
   gpc1_1 gpc2544 (
      {stage1_10[92]},
      {stage2_10[38]}
   );
   gpc1_1 gpc2545 (
      {stage1_10[93]},
      {stage2_10[39]}
   );
   gpc1_1 gpc2546 (
      {stage1_10[94]},
      {stage2_10[40]}
   );
   gpc1_1 gpc2547 (
      {stage1_11[74]},
      {stage2_11[32]}
   );
   gpc1_1 gpc2548 (
      {stage1_11[75]},
      {stage2_11[33]}
   );
   gpc1_1 gpc2549 (
      {stage1_11[76]},
      {stage2_11[34]}
   );
   gpc1_1 gpc2550 (
      {stage1_11[77]},
      {stage2_11[35]}
   );
   gpc1_1 gpc2551 (
      {stage1_11[78]},
      {stage2_11[36]}
   );
   gpc1_1 gpc2552 (
      {stage1_11[79]},
      {stage2_11[37]}
   );
   gpc1_1 gpc2553 (
      {stage1_11[80]},
      {stage2_11[38]}
   );
   gpc1_1 gpc2554 (
      {stage1_12[63]},
      {stage2_12[27]}
   );
   gpc1_1 gpc2555 (
      {stage1_12[64]},
      {stage2_12[28]}
   );
   gpc1_1 gpc2556 (
      {stage1_12[65]},
      {stage2_12[29]}
   );
   gpc1_1 gpc2557 (
      {stage1_12[66]},
      {stage2_12[30]}
   );
   gpc1_1 gpc2558 (
      {stage1_13[66]},
      {stage2_13[24]}
   );
   gpc1_1 gpc2559 (
      {stage1_13[67]},
      {stage2_13[25]}
   );
   gpc1_1 gpc2560 (
      {stage1_13[68]},
      {stage2_13[26]}
   );
   gpc1_1 gpc2561 (
      {stage1_13[69]},
      {stage2_13[27]}
   );
   gpc1_1 gpc2562 (
      {stage1_13[70]},
      {stage2_13[28]}
   );
   gpc1_1 gpc2563 (
      {stage1_13[71]},
      {stage2_13[29]}
   );
   gpc1_1 gpc2564 (
      {stage1_13[72]},
      {stage2_13[30]}
   );
   gpc1_1 gpc2565 (
      {stage1_13[73]},
      {stage2_13[31]}
   );
   gpc1_1 gpc2566 (
      {stage1_13[74]},
      {stage2_13[32]}
   );
   gpc1_1 gpc2567 (
      {stage1_13[75]},
      {stage2_13[33]}
   );
   gpc1_1 gpc2568 (
      {stage1_13[76]},
      {stage2_13[34]}
   );
   gpc1_1 gpc2569 (
      {stage1_13[77]},
      {stage2_13[35]}
   );
   gpc1_1 gpc2570 (
      {stage1_13[78]},
      {stage2_13[36]}
   );
   gpc1_1 gpc2571 (
      {stage1_13[79]},
      {stage2_13[37]}
   );
   gpc1_1 gpc2572 (
      {stage1_13[80]},
      {stage2_13[38]}
   );
   gpc1_1 gpc2573 (
      {stage1_13[81]},
      {stage2_13[39]}
   );
   gpc1_1 gpc2574 (
      {stage1_13[82]},
      {stage2_13[40]}
   );
   gpc1_1 gpc2575 (
      {stage1_13[83]},
      {stage2_13[41]}
   );
   gpc1_1 gpc2576 (
      {stage1_13[84]},
      {stage2_13[42]}
   );
   gpc1_1 gpc2577 (
      {stage1_13[85]},
      {stage2_13[43]}
   );
   gpc1_1 gpc2578 (
      {stage1_13[86]},
      {stage2_13[44]}
   );
   gpc1_1 gpc2579 (
      {stage1_14[10]},
      {stage2_14[22]}
   );
   gpc1_1 gpc2580 (
      {stage1_14[11]},
      {stage2_14[23]}
   );
   gpc1_1 gpc2581 (
      {stage1_14[12]},
      {stage2_14[24]}
   );
   gpc1_1 gpc2582 (
      {stage1_14[13]},
      {stage2_14[25]}
   );
   gpc1_1 gpc2583 (
      {stage1_14[14]},
      {stage2_14[26]}
   );
   gpc1_1 gpc2584 (
      {stage1_14[15]},
      {stage2_14[27]}
   );
   gpc1_1 gpc2585 (
      {stage1_14[16]},
      {stage2_14[28]}
   );
   gpc1_1 gpc2586 (
      {stage1_14[17]},
      {stage2_14[29]}
   );
   gpc1_1 gpc2587 (
      {stage1_14[18]},
      {stage2_14[30]}
   );
   gpc1_1 gpc2588 (
      {stage1_14[19]},
      {stage2_14[31]}
   );
   gpc1_1 gpc2589 (
      {stage1_14[20]},
      {stage2_14[32]}
   );
   gpc1_1 gpc2590 (
      {stage1_14[21]},
      {stage2_14[33]}
   );
   gpc1_1 gpc2591 (
      {stage1_14[22]},
      {stage2_14[34]}
   );
   gpc1_1 gpc2592 (
      {stage1_14[23]},
      {stage2_14[35]}
   );
   gpc1_1 gpc2593 (
      {stage1_14[24]},
      {stage2_14[36]}
   );
   gpc1_1 gpc2594 (
      {stage1_14[25]},
      {stage2_14[37]}
   );
   gpc1_1 gpc2595 (
      {stage1_14[26]},
      {stage2_14[38]}
   );
   gpc1_1 gpc2596 (
      {stage1_14[27]},
      {stage2_14[39]}
   );
   gpc1_1 gpc2597 (
      {stage1_14[28]},
      {stage2_14[40]}
   );
   gpc1_1 gpc2598 (
      {stage1_14[29]},
      {stage2_14[41]}
   );
   gpc1_1 gpc2599 (
      {stage1_14[30]},
      {stage2_14[42]}
   );
   gpc1_1 gpc2600 (
      {stage1_14[31]},
      {stage2_14[43]}
   );
   gpc1_1 gpc2601 (
      {stage1_14[32]},
      {stage2_14[44]}
   );
   gpc1_1 gpc2602 (
      {stage1_14[33]},
      {stage2_14[45]}
   );
   gpc1_1 gpc2603 (
      {stage1_14[34]},
      {stage2_14[46]}
   );
   gpc1_1 gpc2604 (
      {stage1_14[35]},
      {stage2_14[47]}
   );
   gpc1_1 gpc2605 (
      {stage1_14[36]},
      {stage2_14[48]}
   );
   gpc1_1 gpc2606 (
      {stage1_14[37]},
      {stage2_14[49]}
   );
   gpc1_1 gpc2607 (
      {stage1_14[38]},
      {stage2_14[50]}
   );
   gpc1_1 gpc2608 (
      {stage1_14[39]},
      {stage2_14[51]}
   );
   gpc1_1 gpc2609 (
      {stage1_14[40]},
      {stage2_14[52]}
   );
   gpc1_1 gpc2610 (
      {stage1_14[41]},
      {stage2_14[53]}
   );
   gpc1_1 gpc2611 (
      {stage1_14[42]},
      {stage2_14[54]}
   );
   gpc1_1 gpc2612 (
      {stage1_14[43]},
      {stage2_14[55]}
   );
   gpc1_1 gpc2613 (
      {stage1_14[44]},
      {stage2_14[56]}
   );
   gpc1_1 gpc2614 (
      {stage1_14[45]},
      {stage2_14[57]}
   );
   gpc1_1 gpc2615 (
      {stage1_14[46]},
      {stage2_14[58]}
   );
   gpc1_1 gpc2616 (
      {stage1_14[47]},
      {stage2_14[59]}
   );
   gpc1_1 gpc2617 (
      {stage1_14[48]},
      {stage2_14[60]}
   );
   gpc1_1 gpc2618 (
      {stage1_14[49]},
      {stage2_14[61]}
   );
   gpc1_1 gpc2619 (
      {stage1_14[50]},
      {stage2_14[62]}
   );
   gpc1_1 gpc2620 (
      {stage1_14[51]},
      {stage2_14[63]}
   );
   gpc1_1 gpc2621 (
      {stage1_14[52]},
      {stage2_14[64]}
   );
   gpc1_1 gpc2622 (
      {stage1_14[53]},
      {stage2_14[65]}
   );
   gpc1_1 gpc2623 (
      {stage1_14[54]},
      {stage2_14[66]}
   );
   gpc1_1 gpc2624 (
      {stage1_14[55]},
      {stage2_14[67]}
   );
   gpc1_1 gpc2625 (
      {stage1_14[56]},
      {stage2_14[68]}
   );
   gpc1_1 gpc2626 (
      {stage1_14[57]},
      {stage2_14[69]}
   );
   gpc1_1 gpc2627 (
      {stage1_14[58]},
      {stage2_14[70]}
   );
   gpc1_1 gpc2628 (
      {stage1_14[59]},
      {stage2_14[71]}
   );
   gpc1_1 gpc2629 (
      {stage1_14[60]},
      {stage2_14[72]}
   );
   gpc1_1 gpc2630 (
      {stage1_14[61]},
      {stage2_14[73]}
   );
   gpc1_1 gpc2631 (
      {stage1_15[86]},
      {stage2_15[25]}
   );
   gpc1_1 gpc2632 (
      {stage1_15[87]},
      {stage2_15[26]}
   );
   gpc1_1 gpc2633 (
      {stage1_15[88]},
      {stage2_15[27]}
   );
   gpc1_1 gpc2634 (
      {stage1_15[89]},
      {stage2_15[28]}
   );
   gpc1_1 gpc2635 (
      {stage1_15[90]},
      {stage2_15[29]}
   );
   gpc1_1 gpc2636 (
      {stage1_15[91]},
      {stage2_15[30]}
   );
   gpc1_1 gpc2637 (
      {stage1_15[92]},
      {stage2_15[31]}
   );
   gpc1_1 gpc2638 (
      {stage1_15[93]},
      {stage2_15[32]}
   );
   gpc1_1 gpc2639 (
      {stage1_15[94]},
      {stage2_15[33]}
   );
   gpc1_1 gpc2640 (
      {stage1_15[95]},
      {stage2_15[34]}
   );
   gpc1_1 gpc2641 (
      {stage1_15[96]},
      {stage2_15[35]}
   );
   gpc1_1 gpc2642 (
      {stage1_15[97]},
      {stage2_15[36]}
   );
   gpc1_1 gpc2643 (
      {stage1_16[42]},
      {stage2_16[21]}
   );
   gpc1_1 gpc2644 (
      {stage1_16[43]},
      {stage2_16[22]}
   );
   gpc1_1 gpc2645 (
      {stage1_16[44]},
      {stage2_16[23]}
   );
   gpc1_1 gpc2646 (
      {stage1_16[45]},
      {stage2_16[24]}
   );
   gpc1_1 gpc2647 (
      {stage1_16[46]},
      {stage2_16[25]}
   );
   gpc1_1 gpc2648 (
      {stage1_16[47]},
      {stage2_16[26]}
   );
   gpc1_1 gpc2649 (
      {stage1_16[48]},
      {stage2_16[27]}
   );
   gpc1_1 gpc2650 (
      {stage1_16[49]},
      {stage2_16[28]}
   );
   gpc1_1 gpc2651 (
      {stage1_16[50]},
      {stage2_16[29]}
   );
   gpc1_1 gpc2652 (
      {stage1_16[51]},
      {stage2_16[30]}
   );
   gpc1_1 gpc2653 (
      {stage1_16[52]},
      {stage2_16[31]}
   );
   gpc1_1 gpc2654 (
      {stage1_16[53]},
      {stage2_16[32]}
   );
   gpc1_1 gpc2655 (
      {stage1_16[54]},
      {stage2_16[33]}
   );
   gpc1_1 gpc2656 (
      {stage1_16[55]},
      {stage2_16[34]}
   );
   gpc1_1 gpc2657 (
      {stage1_16[56]},
      {stage2_16[35]}
   );
   gpc1_1 gpc2658 (
      {stage1_16[57]},
      {stage2_16[36]}
   );
   gpc1_1 gpc2659 (
      {stage1_16[58]},
      {stage2_16[37]}
   );
   gpc1_1 gpc2660 (
      {stage1_16[59]},
      {stage2_16[38]}
   );
   gpc1_1 gpc2661 (
      {stage1_16[60]},
      {stage2_16[39]}
   );
   gpc1_1 gpc2662 (
      {stage1_16[61]},
      {stage2_16[40]}
   );
   gpc1_1 gpc2663 (
      {stage1_16[62]},
      {stage2_16[41]}
   );
   gpc1_1 gpc2664 (
      {stage1_16[63]},
      {stage2_16[42]}
   );
   gpc1_1 gpc2665 (
      {stage1_16[64]},
      {stage2_16[43]}
   );
   gpc1_1 gpc2666 (
      {stage1_16[65]},
      {stage2_16[44]}
   );
   gpc1_1 gpc2667 (
      {stage1_16[66]},
      {stage2_16[45]}
   );
   gpc1_1 gpc2668 (
      {stage1_16[67]},
      {stage2_16[46]}
   );
   gpc1_1 gpc2669 (
      {stage1_17[100]},
      {stage2_17[26]}
   );
   gpc1_1 gpc2670 (
      {stage1_17[101]},
      {stage2_17[27]}
   );
   gpc1_1 gpc2671 (
      {stage1_17[102]},
      {stage2_17[28]}
   );
   gpc1_1 gpc2672 (
      {stage1_17[103]},
      {stage2_17[29]}
   );
   gpc1_1 gpc2673 (
      {stage1_17[104]},
      {stage2_17[30]}
   );
   gpc1_1 gpc2674 (
      {stage1_17[105]},
      {stage2_17[31]}
   );
   gpc1_1 gpc2675 (
      {stage1_17[106]},
      {stage2_17[32]}
   );
   gpc1_1 gpc2676 (
      {stage1_17[107]},
      {stage2_17[33]}
   );
   gpc1_1 gpc2677 (
      {stage1_17[108]},
      {stage2_17[34]}
   );
   gpc1_1 gpc2678 (
      {stage1_17[109]},
      {stage2_17[35]}
   );
   gpc1_1 gpc2679 (
      {stage1_17[110]},
      {stage2_17[36]}
   );
   gpc1_1 gpc2680 (
      {stage1_17[111]},
      {stage2_17[37]}
   );
   gpc1_1 gpc2681 (
      {stage1_17[112]},
      {stage2_17[38]}
   );
   gpc1_1 gpc2682 (
      {stage1_17[113]},
      {stage2_17[39]}
   );
   gpc1_1 gpc2683 (
      {stage1_18[47]},
      {stage2_18[27]}
   );
   gpc1_1 gpc2684 (
      {stage1_18[48]},
      {stage2_18[28]}
   );
   gpc1_1 gpc2685 (
      {stage1_18[49]},
      {stage2_18[29]}
   );
   gpc1_1 gpc2686 (
      {stage1_18[50]},
      {stage2_18[30]}
   );
   gpc1_1 gpc2687 (
      {stage1_18[51]},
      {stage2_18[31]}
   );
   gpc1_1 gpc2688 (
      {stage1_18[52]},
      {stage2_18[32]}
   );
   gpc1_1 gpc2689 (
      {stage1_18[53]},
      {stage2_18[33]}
   );
   gpc1_1 gpc2690 (
      {stage1_18[54]},
      {stage2_18[34]}
   );
   gpc1_1 gpc2691 (
      {stage1_18[55]},
      {stage2_18[35]}
   );
   gpc1_1 gpc2692 (
      {stage1_18[56]},
      {stage2_18[36]}
   );
   gpc1_1 gpc2693 (
      {stage1_18[57]},
      {stage2_18[37]}
   );
   gpc1_1 gpc2694 (
      {stage1_18[58]},
      {stage2_18[38]}
   );
   gpc1_1 gpc2695 (
      {stage1_18[59]},
      {stage2_18[39]}
   );
   gpc1_1 gpc2696 (
      {stage1_18[60]},
      {stage2_18[40]}
   );
   gpc1_1 gpc2697 (
      {stage1_18[61]},
      {stage2_18[41]}
   );
   gpc1_1 gpc2698 (
      {stage1_18[62]},
      {stage2_18[42]}
   );
   gpc1_1 gpc2699 (
      {stage1_19[48]},
      {stage2_19[28]}
   );
   gpc1_1 gpc2700 (
      {stage1_19[49]},
      {stage2_19[29]}
   );
   gpc1_1 gpc2701 (
      {stage1_19[50]},
      {stage2_19[30]}
   );
   gpc1_1 gpc2702 (
      {stage1_19[51]},
      {stage2_19[31]}
   );
   gpc1_1 gpc2703 (
      {stage1_19[52]},
      {stage2_19[32]}
   );
   gpc1_1 gpc2704 (
      {stage1_19[53]},
      {stage2_19[33]}
   );
   gpc1_1 gpc2705 (
      {stage1_19[54]},
      {stage2_19[34]}
   );
   gpc1_1 gpc2706 (
      {stage1_19[55]},
      {stage2_19[35]}
   );
   gpc1_1 gpc2707 (
      {stage1_19[56]},
      {stage2_19[36]}
   );
   gpc1_1 gpc2708 (
      {stage1_19[57]},
      {stage2_19[37]}
   );
   gpc1_1 gpc2709 (
      {stage1_19[58]},
      {stage2_19[38]}
   );
   gpc1_1 gpc2710 (
      {stage1_19[59]},
      {stage2_19[39]}
   );
   gpc1_1 gpc2711 (
      {stage1_19[60]},
      {stage2_19[40]}
   );
   gpc1_1 gpc2712 (
      {stage1_19[61]},
      {stage2_19[41]}
   );
   gpc1_1 gpc2713 (
      {stage1_19[62]},
      {stage2_19[42]}
   );
   gpc1_1 gpc2714 (
      {stage1_19[63]},
      {stage2_19[43]}
   );
   gpc1_1 gpc2715 (
      {stage1_19[64]},
      {stage2_19[44]}
   );
   gpc1_1 gpc2716 (
      {stage1_19[65]},
      {stage2_19[45]}
   );
   gpc1_1 gpc2717 (
      {stage1_19[66]},
      {stage2_19[46]}
   );
   gpc1_1 gpc2718 (
      {stage1_19[67]},
      {stage2_19[47]}
   );
   gpc1_1 gpc2719 (
      {stage1_19[68]},
      {stage2_19[48]}
   );
   gpc1_1 gpc2720 (
      {stage1_19[69]},
      {stage2_19[49]}
   );
   gpc1_1 gpc2721 (
      {stage1_19[70]},
      {stage2_19[50]}
   );
   gpc1_1 gpc2722 (
      {stage1_20[27]},
      {stage2_20[17]}
   );
   gpc1_1 gpc2723 (
      {stage1_20[28]},
      {stage2_20[18]}
   );
   gpc1_1 gpc2724 (
      {stage1_20[29]},
      {stage2_20[19]}
   );
   gpc1_1 gpc2725 (
      {stage1_20[30]},
      {stage2_20[20]}
   );
   gpc1_1 gpc2726 (
      {stage1_20[31]},
      {stage2_20[21]}
   );
   gpc1_1 gpc2727 (
      {stage1_20[32]},
      {stage2_20[22]}
   );
   gpc1_1 gpc2728 (
      {stage1_20[33]},
      {stage2_20[23]}
   );
   gpc1_1 gpc2729 (
      {stage1_20[34]},
      {stage2_20[24]}
   );
   gpc1_1 gpc2730 (
      {stage1_20[35]},
      {stage2_20[25]}
   );
   gpc1_1 gpc2731 (
      {stage1_20[36]},
      {stage2_20[26]}
   );
   gpc1_1 gpc2732 (
      {stage1_20[37]},
      {stage2_20[27]}
   );
   gpc1_1 gpc2733 (
      {stage1_20[38]},
      {stage2_20[28]}
   );
   gpc1_1 gpc2734 (
      {stage1_20[39]},
      {stage2_20[29]}
   );
   gpc1_1 gpc2735 (
      {stage1_20[40]},
      {stage2_20[30]}
   );
   gpc1_1 gpc2736 (
      {stage1_20[41]},
      {stage2_20[31]}
   );
   gpc1_1 gpc2737 (
      {stage1_20[42]},
      {stage2_20[32]}
   );
   gpc1_1 gpc2738 (
      {stage1_20[43]},
      {stage2_20[33]}
   );
   gpc1_1 gpc2739 (
      {stage1_20[44]},
      {stage2_20[34]}
   );
   gpc1_1 gpc2740 (
      {stage1_20[45]},
      {stage2_20[35]}
   );
   gpc1_1 gpc2741 (
      {stage1_20[46]},
      {stage2_20[36]}
   );
   gpc1_1 gpc2742 (
      {stage1_20[47]},
      {stage2_20[37]}
   );
   gpc1_1 gpc2743 (
      {stage1_20[48]},
      {stage2_20[38]}
   );
   gpc1_1 gpc2744 (
      {stage1_20[49]},
      {stage2_20[39]}
   );
   gpc1_1 gpc2745 (
      {stage1_20[50]},
      {stage2_20[40]}
   );
   gpc1_1 gpc2746 (
      {stage1_20[51]},
      {stage2_20[41]}
   );
   gpc1_1 gpc2747 (
      {stage1_20[52]},
      {stage2_20[42]}
   );
   gpc1_1 gpc2748 (
      {stage1_20[53]},
      {stage2_20[43]}
   );
   gpc1_1 gpc2749 (
      {stage1_20[54]},
      {stage2_20[44]}
   );
   gpc1_1 gpc2750 (
      {stage1_20[55]},
      {stage2_20[45]}
   );
   gpc1_1 gpc2751 (
      {stage1_20[56]},
      {stage2_20[46]}
   );
   gpc1_1 gpc2752 (
      {stage1_20[57]},
      {stage2_20[47]}
   );
   gpc1_1 gpc2753 (
      {stage1_20[58]},
      {stage2_20[48]}
   );
   gpc1_1 gpc2754 (
      {stage1_20[59]},
      {stage2_20[49]}
   );
   gpc1_1 gpc2755 (
      {stage1_20[60]},
      {stage2_20[50]}
   );
   gpc1_1 gpc2756 (
      {stage1_20[61]},
      {stage2_20[51]}
   );
   gpc1_1 gpc2757 (
      {stage1_20[62]},
      {stage2_20[52]}
   );
   gpc1_1 gpc2758 (
      {stage1_20[63]},
      {stage2_20[53]}
   );
   gpc1_1 gpc2759 (
      {stage1_20[64]},
      {stage2_20[54]}
   );
   gpc1_1 gpc2760 (
      {stage1_20[65]},
      {stage2_20[55]}
   );
   gpc1_1 gpc2761 (
      {stage1_20[66]},
      {stage2_20[56]}
   );
   gpc1_1 gpc2762 (
      {stage1_20[67]},
      {stage2_20[57]}
   );
   gpc1_1 gpc2763 (
      {stage1_21[48]},
      {stage2_21[17]}
   );
   gpc1_1 gpc2764 (
      {stage1_21[49]},
      {stage2_21[18]}
   );
   gpc1_1 gpc2765 (
      {stage1_21[50]},
      {stage2_21[19]}
   );
   gpc1_1 gpc2766 (
      {stage1_21[51]},
      {stage2_21[20]}
   );
   gpc1_1 gpc2767 (
      {stage1_21[52]},
      {stage2_21[21]}
   );
   gpc1_1 gpc2768 (
      {stage1_21[53]},
      {stage2_21[22]}
   );
   gpc1_1 gpc2769 (
      {stage1_21[54]},
      {stage2_21[23]}
   );
   gpc1_1 gpc2770 (
      {stage1_21[55]},
      {stage2_21[24]}
   );
   gpc1_1 gpc2771 (
      {stage1_21[56]},
      {stage2_21[25]}
   );
   gpc1_1 gpc2772 (
      {stage1_21[57]},
      {stage2_21[26]}
   );
   gpc1_1 gpc2773 (
      {stage1_21[58]},
      {stage2_21[27]}
   );
   gpc1_1 gpc2774 (
      {stage1_21[59]},
      {stage2_21[28]}
   );
   gpc1_1 gpc2775 (
      {stage1_21[60]},
      {stage2_21[29]}
   );
   gpc1_1 gpc2776 (
      {stage1_21[61]},
      {stage2_21[30]}
   );
   gpc1_1 gpc2777 (
      {stage1_21[62]},
      {stage2_21[31]}
   );
   gpc1_1 gpc2778 (
      {stage1_21[63]},
      {stage2_21[32]}
   );
   gpc1_1 gpc2779 (
      {stage1_21[64]},
      {stage2_21[33]}
   );
   gpc1_1 gpc2780 (
      {stage1_21[65]},
      {stage2_21[34]}
   );
   gpc1_1 gpc2781 (
      {stage1_21[66]},
      {stage2_21[35]}
   );
   gpc1_1 gpc2782 (
      {stage1_21[67]},
      {stage2_21[36]}
   );
   gpc1_1 gpc2783 (
      {stage1_21[68]},
      {stage2_21[37]}
   );
   gpc1_1 gpc2784 (
      {stage1_21[69]},
      {stage2_21[38]}
   );
   gpc1_1 gpc2785 (
      {stage1_21[70]},
      {stage2_21[39]}
   );
   gpc1_1 gpc2786 (
      {stage1_22[62]},
      {stage2_22[26]}
   );
   gpc1_1 gpc2787 (
      {stage1_22[63]},
      {stage2_22[27]}
   );
   gpc1_1 gpc2788 (
      {stage1_22[64]},
      {stage2_22[28]}
   );
   gpc1_1 gpc2789 (
      {stage1_22[65]},
      {stage2_22[29]}
   );
   gpc1_1 gpc2790 (
      {stage1_22[66]},
      {stage2_22[30]}
   );
   gpc1_1 gpc2791 (
      {stage1_23[127]},
      {stage2_23[31]}
   );
   gpc1_1 gpc2792 (
      {stage1_23[128]},
      {stage2_23[32]}
   );
   gpc1_1 gpc2793 (
      {stage1_23[129]},
      {stage2_23[33]}
   );
   gpc1_1 gpc2794 (
      {stage1_23[130]},
      {stage2_23[34]}
   );
   gpc1_1 gpc2795 (
      {stage1_23[131]},
      {stage2_23[35]}
   );
   gpc1_1 gpc2796 (
      {stage1_23[132]},
      {stage2_23[36]}
   );
   gpc1_1 gpc2797 (
      {stage1_23[133]},
      {stage2_23[37]}
   );
   gpc1_1 gpc2798 (
      {stage1_23[134]},
      {stage2_23[38]}
   );
   gpc1_1 gpc2799 (
      {stage1_23[135]},
      {stage2_23[39]}
   );
   gpc1_1 gpc2800 (
      {stage1_23[136]},
      {stage2_23[40]}
   );
   gpc1_1 gpc2801 (
      {stage1_23[137]},
      {stage2_23[41]}
   );
   gpc1_1 gpc2802 (
      {stage1_23[138]},
      {stage2_23[42]}
   );
   gpc1_1 gpc2803 (
      {stage1_23[139]},
      {stage2_23[43]}
   );
   gpc1_1 gpc2804 (
      {stage1_23[140]},
      {stage2_23[44]}
   );
   gpc1_1 gpc2805 (
      {stage1_23[141]},
      {stage2_23[45]}
   );
   gpc1_1 gpc2806 (
      {stage1_23[142]},
      {stage2_23[46]}
   );
   gpc1_1 gpc2807 (
      {stage1_24[69]},
      {stage2_24[32]}
   );
   gpc1_1 gpc2808 (
      {stage1_24[70]},
      {stage2_24[33]}
   );
   gpc1_1 gpc2809 (
      {stage1_24[71]},
      {stage2_24[34]}
   );
   gpc1_1 gpc2810 (
      {stage1_24[72]},
      {stage2_24[35]}
   );
   gpc1_1 gpc2811 (
      {stage1_24[73]},
      {stage2_24[36]}
   );
   gpc1_1 gpc2812 (
      {stage1_24[74]},
      {stage2_24[37]}
   );
   gpc1_1 gpc2813 (
      {stage1_24[75]},
      {stage2_24[38]}
   );
   gpc1_1 gpc2814 (
      {stage1_24[76]},
      {stage2_24[39]}
   );
   gpc1_1 gpc2815 (
      {stage1_24[77]},
      {stage2_24[40]}
   );
   gpc1_1 gpc2816 (
      {stage1_24[78]},
      {stage2_24[41]}
   );
   gpc1_1 gpc2817 (
      {stage1_24[79]},
      {stage2_24[42]}
   );
   gpc1_1 gpc2818 (
      {stage1_24[80]},
      {stage2_24[43]}
   );
   gpc1_1 gpc2819 (
      {stage1_24[81]},
      {stage2_24[44]}
   );
   gpc1_1 gpc2820 (
      {stage1_24[82]},
      {stage2_24[45]}
   );
   gpc1_1 gpc2821 (
      {stage1_25[83]},
      {stage2_25[35]}
   );
   gpc1_1 gpc2822 (
      {stage1_25[84]},
      {stage2_25[36]}
   );
   gpc1_1 gpc2823 (
      {stage1_26[54]},
      {stage2_26[35]}
   );
   gpc1_1 gpc2824 (
      {stage1_26[55]},
      {stage2_26[36]}
   );
   gpc1_1 gpc2825 (
      {stage1_26[56]},
      {stage2_26[37]}
   );
   gpc1_1 gpc2826 (
      {stage1_26[57]},
      {stage2_26[38]}
   );
   gpc1_1 gpc2827 (
      {stage1_26[58]},
      {stage2_26[39]}
   );
   gpc1_1 gpc2828 (
      {stage1_26[59]},
      {stage2_26[40]}
   );
   gpc1_1 gpc2829 (
      {stage1_26[60]},
      {stage2_26[41]}
   );
   gpc1_1 gpc2830 (
      {stage1_26[61]},
      {stage2_26[42]}
   );
   gpc1_1 gpc2831 (
      {stage1_26[62]},
      {stage2_26[43]}
   );
   gpc1_1 gpc2832 (
      {stage1_26[63]},
      {stage2_26[44]}
   );
   gpc1_1 gpc2833 (
      {stage1_26[64]},
      {stage2_26[45]}
   );
   gpc1_1 gpc2834 (
      {stage1_26[65]},
      {stage2_26[46]}
   );
   gpc1_1 gpc2835 (
      {stage1_26[66]},
      {stage2_26[47]}
   );
   gpc1_1 gpc2836 (
      {stage1_26[67]},
      {stage2_26[48]}
   );
   gpc1_1 gpc2837 (
      {stage1_26[68]},
      {stage2_26[49]}
   );
   gpc1_1 gpc2838 (
      {stage1_26[69]},
      {stage2_26[50]}
   );
   gpc1_1 gpc2839 (
      {stage1_26[70]},
      {stage2_26[51]}
   );
   gpc1_1 gpc2840 (
      {stage1_26[71]},
      {stage2_26[52]}
   );
   gpc1_1 gpc2841 (
      {stage1_27[49]},
      {stage2_27[25]}
   );
   gpc1_1 gpc2842 (
      {stage1_27[50]},
      {stage2_27[26]}
   );
   gpc1_1 gpc2843 (
      {stage1_27[51]},
      {stage2_27[27]}
   );
   gpc1_1 gpc2844 (
      {stage1_27[52]},
      {stage2_27[28]}
   );
   gpc1_1 gpc2845 (
      {stage1_27[53]},
      {stage2_27[29]}
   );
   gpc1_1 gpc2846 (
      {stage1_27[54]},
      {stage2_27[30]}
   );
   gpc1_1 gpc2847 (
      {stage1_27[55]},
      {stage2_27[31]}
   );
   gpc1_1 gpc2848 (
      {stage1_27[56]},
      {stage2_27[32]}
   );
   gpc1_1 gpc2849 (
      {stage1_27[57]},
      {stage2_27[33]}
   );
   gpc1_1 gpc2850 (
      {stage1_27[58]},
      {stage2_27[34]}
   );
   gpc1_1 gpc2851 (
      {stage1_27[59]},
      {stage2_27[35]}
   );
   gpc1_1 gpc2852 (
      {stage1_27[60]},
      {stage2_27[36]}
   );
   gpc1_1 gpc2853 (
      {stage1_27[61]},
      {stage2_27[37]}
   );
   gpc1_1 gpc2854 (
      {stage1_27[62]},
      {stage2_27[38]}
   );
   gpc1_1 gpc2855 (
      {stage1_27[63]},
      {stage2_27[39]}
   );
   gpc1_1 gpc2856 (
      {stage1_27[64]},
      {stage2_27[40]}
   );
   gpc1_1 gpc2857 (
      {stage1_27[65]},
      {stage2_27[41]}
   );
   gpc1_1 gpc2858 (
      {stage1_27[66]},
      {stage2_27[42]}
   );
   gpc1_1 gpc2859 (
      {stage1_27[67]},
      {stage2_27[43]}
   );
   gpc1_1 gpc2860 (
      {stage1_27[68]},
      {stage2_27[44]}
   );
   gpc1_1 gpc2861 (
      {stage1_27[69]},
      {stage2_27[45]}
   );
   gpc1_1 gpc2862 (
      {stage1_27[70]},
      {stage2_27[46]}
   );
   gpc1_1 gpc2863 (
      {stage1_27[71]},
      {stage2_27[47]}
   );
   gpc1_1 gpc2864 (
      {stage1_27[72]},
      {stage2_27[48]}
   );
   gpc1_1 gpc2865 (
      {stage1_27[73]},
      {stage2_27[49]}
   );
   gpc1_1 gpc2866 (
      {stage1_28[69]},
      {stage2_28[27]}
   );
   gpc1_1 gpc2867 (
      {stage1_28[70]},
      {stage2_28[28]}
   );
   gpc1_1 gpc2868 (
      {stage1_28[71]},
      {stage2_28[29]}
   );
   gpc1_1 gpc2869 (
      {stage1_28[72]},
      {stage2_28[30]}
   );
   gpc1_1 gpc2870 (
      {stage1_28[73]},
      {stage2_28[31]}
   );
   gpc1_1 gpc2871 (
      {stage1_28[74]},
      {stage2_28[32]}
   );
   gpc1_1 gpc2872 (
      {stage1_28[75]},
      {stage2_28[33]}
   );
   gpc1_1 gpc2873 (
      {stage1_28[76]},
      {stage2_28[34]}
   );
   gpc1_1 gpc2874 (
      {stage1_29[58]},
      {stage2_29[27]}
   );
   gpc1_1 gpc2875 (
      {stage1_29[59]},
      {stage2_29[28]}
   );
   gpc1_1 gpc2876 (
      {stage1_29[60]},
      {stage2_29[29]}
   );
   gpc1_1 gpc2877 (
      {stage1_29[61]},
      {stage2_29[30]}
   );
   gpc1_1 gpc2878 (
      {stage1_29[62]},
      {stage2_29[31]}
   );
   gpc1_1 gpc2879 (
      {stage1_29[63]},
      {stage2_29[32]}
   );
   gpc1_1 gpc2880 (
      {stage1_29[64]},
      {stage2_29[33]}
   );
   gpc1_1 gpc2881 (
      {stage1_29[65]},
      {stage2_29[34]}
   );
   gpc1_1 gpc2882 (
      {stage1_29[66]},
      {stage2_29[35]}
   );
   gpc1_1 gpc2883 (
      {stage1_29[67]},
      {stage2_29[36]}
   );
   gpc1_1 gpc2884 (
      {stage1_29[68]},
      {stage2_29[37]}
   );
   gpc1_1 gpc2885 (
      {stage1_29[69]},
      {stage2_29[38]}
   );
   gpc1_1 gpc2886 (
      {stage1_29[70]},
      {stage2_29[39]}
   );
   gpc1_1 gpc2887 (
      {stage1_29[71]},
      {stage2_29[40]}
   );
   gpc1_1 gpc2888 (
      {stage1_29[72]},
      {stage2_29[41]}
   );
   gpc1_1 gpc2889 (
      {stage1_29[73]},
      {stage2_29[42]}
   );
   gpc1_1 gpc2890 (
      {stage1_29[74]},
      {stage2_29[43]}
   );
   gpc1_1 gpc2891 (
      {stage1_29[75]},
      {stage2_29[44]}
   );
   gpc1_1 gpc2892 (
      {stage1_29[76]},
      {stage2_29[45]}
   );
   gpc1_1 gpc2893 (
      {stage1_29[77]},
      {stage2_29[46]}
   );
   gpc1_1 gpc2894 (
      {stage1_29[78]},
      {stage2_29[47]}
   );
   gpc1_1 gpc2895 (
      {stage1_29[79]},
      {stage2_29[48]}
   );
   gpc1_1 gpc2896 (
      {stage1_29[80]},
      {stage2_29[49]}
   );
   gpc1_1 gpc2897 (
      {stage1_30[84]},
      {stage2_30[27]}
   );
   gpc1_1 gpc2898 (
      {stage1_30[85]},
      {stage2_30[28]}
   );
   gpc1_1 gpc2899 (
      {stage1_30[86]},
      {stage2_30[29]}
   );
   gpc1_1 gpc2900 (
      {stage1_30[87]},
      {stage2_30[30]}
   );
   gpc1_1 gpc2901 (
      {stage1_30[88]},
      {stage2_30[31]}
   );
   gpc1_1 gpc2902 (
      {stage1_30[89]},
      {stage2_30[32]}
   );
   gpc1_1 gpc2903 (
      {stage1_30[90]},
      {stage2_30[33]}
   );
   gpc1_1 gpc2904 (
      {stage1_30[91]},
      {stage2_30[34]}
   );
   gpc1_1 gpc2905 (
      {stage1_30[92]},
      {stage2_30[35]}
   );
   gpc1_1 gpc2906 (
      {stage1_30[93]},
      {stage2_30[36]}
   );
   gpc1_1 gpc2907 (
      {stage1_30[94]},
      {stage2_30[37]}
   );
   gpc1_1 gpc2908 (
      {stage1_30[95]},
      {stage2_30[38]}
   );
   gpc1_1 gpc2909 (
      {stage1_30[96]},
      {stage2_30[39]}
   );
   gpc1_1 gpc2910 (
      {stage1_30[97]},
      {stage2_30[40]}
   );
   gpc1_1 gpc2911 (
      {stage1_30[98]},
      {stage2_30[41]}
   );
   gpc1_1 gpc2912 (
      {stage1_30[99]},
      {stage2_30[42]}
   );
   gpc1_1 gpc2913 (
      {stage1_30[100]},
      {stage2_30[43]}
   );
   gpc1_1 gpc2914 (
      {stage1_30[101]},
      {stage2_30[44]}
   );
   gpc1_1 gpc2915 (
      {stage1_30[102]},
      {stage2_30[45]}
   );
   gpc1_1 gpc2916 (
      {stage1_30[103]},
      {stage2_30[46]}
   );
   gpc1_1 gpc2917 (
      {stage1_30[104]},
      {stage2_30[47]}
   );
   gpc1_1 gpc2918 (
      {stage1_30[105]},
      {stage2_30[48]}
   );
   gpc1_1 gpc2919 (
      {stage1_30[106]},
      {stage2_30[49]}
   );
   gpc1_1 gpc2920 (
      {stage1_31[94]},
      {stage2_31[36]}
   );
   gpc1_1 gpc2921 (
      {stage1_31[95]},
      {stage2_31[37]}
   );
   gpc1_1 gpc2922 (
      {stage1_31[96]},
      {stage2_31[38]}
   );
   gpc1_1 gpc2923 (
      {stage1_32[68]},
      {stage2_32[37]}
   );
   gpc1_1 gpc2924 (
      {stage1_32[69]},
      {stage2_32[38]}
   );
   gpc1_1 gpc2925 (
      {stage1_32[70]},
      {stage2_32[39]}
   );
   gpc1_1 gpc2926 (
      {stage1_32[71]},
      {stage2_32[40]}
   );
   gpc1_1 gpc2927 (
      {stage1_32[72]},
      {stage2_32[41]}
   );
   gpc1_1 gpc2928 (
      {stage1_32[73]},
      {stage2_32[42]}
   );
   gpc1_1 gpc2929 (
      {stage1_32[74]},
      {stage2_32[43]}
   );
   gpc1_1 gpc2930 (
      {stage1_32[75]},
      {stage2_32[44]}
   );
   gpc1_1 gpc2931 (
      {stage1_32[76]},
      {stage2_32[45]}
   );
   gpc1_1 gpc2932 (
      {stage1_32[77]},
      {stage2_32[46]}
   );
   gpc1_1 gpc2933 (
      {stage1_32[78]},
      {stage2_32[47]}
   );
   gpc1_1 gpc2934 (
      {stage1_32[79]},
      {stage2_32[48]}
   );
   gpc1_1 gpc2935 (
      {stage1_32[80]},
      {stage2_32[49]}
   );
   gpc1_1 gpc2936 (
      {stage1_32[81]},
      {stage2_32[50]}
   );
   gpc1_1 gpc2937 (
      {stage1_32[82]},
      {stage2_32[51]}
   );
   gpc1_1 gpc2938 (
      {stage1_32[83]},
      {stage2_32[52]}
   );
   gpc1_1 gpc2939 (
      {stage1_32[84]},
      {stage2_32[53]}
   );
   gpc1_1 gpc2940 (
      {stage1_32[85]},
      {stage2_32[54]}
   );
   gpc1_1 gpc2941 (
      {stage1_32[86]},
      {stage2_32[55]}
   );
   gpc1_1 gpc2942 (
      {stage1_34[48]},
      {stage2_34[27]}
   );
   gpc1_1 gpc2943 (
      {stage1_34[49]},
      {stage2_34[28]}
   );
   gpc1_1 gpc2944 (
      {stage1_34[50]},
      {stage2_34[29]}
   );
   gpc1_1 gpc2945 (
      {stage1_34[51]},
      {stage2_34[30]}
   );
   gpc1_1 gpc2946 (
      {stage1_34[52]},
      {stage2_34[31]}
   );
   gpc1_1 gpc2947 (
      {stage1_34[53]},
      {stage2_34[32]}
   );
   gpc1_1 gpc2948 (
      {stage1_34[54]},
      {stage2_34[33]}
   );
   gpc1_1 gpc2949 (
      {stage1_34[55]},
      {stage2_34[34]}
   );
   gpc1_1 gpc2950 (
      {stage1_35[46]},
      {stage2_35[31]}
   );
   gpc1_1 gpc2951 (
      {stage1_35[47]},
      {stage2_35[32]}
   );
   gpc1_1 gpc2952 (
      {stage1_35[48]},
      {stage2_35[33]}
   );
   gpc1_1 gpc2953 (
      {stage1_35[49]},
      {stage2_35[34]}
   );
   gpc1_1 gpc2954 (
      {stage1_35[50]},
      {stage2_35[35]}
   );
   gpc1_1 gpc2955 (
      {stage1_35[51]},
      {stage2_35[36]}
   );
   gpc1_1 gpc2956 (
      {stage1_35[52]},
      {stage2_35[37]}
   );
   gpc1_1 gpc2957 (
      {stage1_35[53]},
      {stage2_35[38]}
   );
   gpc1_1 gpc2958 (
      {stage1_35[54]},
      {stage2_35[39]}
   );
   gpc1_1 gpc2959 (
      {stage1_35[55]},
      {stage2_35[40]}
   );
   gpc1_1 gpc2960 (
      {stage1_35[56]},
      {stage2_35[41]}
   );
   gpc1_1 gpc2961 (
      {stage1_35[57]},
      {stage2_35[42]}
   );
   gpc1_1 gpc2962 (
      {stage1_35[58]},
      {stage2_35[43]}
   );
   gpc1_1 gpc2963 (
      {stage1_35[59]},
      {stage2_35[44]}
   );
   gpc1_1 gpc2964 (
      {stage1_36[72]},
      {stage2_36[26]}
   );
   gpc1_1 gpc2965 (
      {stage1_36[73]},
      {stage2_36[27]}
   );
   gpc1_1 gpc2966 (
      {stage1_36[74]},
      {stage2_36[28]}
   );
   gpc1_1 gpc2967 (
      {stage1_36[75]},
      {stage2_36[29]}
   );
   gpc1_1 gpc2968 (
      {stage1_36[76]},
      {stage2_36[30]}
   );
   gpc1_1 gpc2969 (
      {stage1_36[77]},
      {stage2_36[31]}
   );
   gpc1_1 gpc2970 (
      {stage1_36[78]},
      {stage2_36[32]}
   );
   gpc1_1 gpc2971 (
      {stage1_36[79]},
      {stage2_36[33]}
   );
   gpc1_1 gpc2972 (
      {stage1_36[80]},
      {stage2_36[34]}
   );
   gpc1_1 gpc2973 (
      {stage1_36[81]},
      {stage2_36[35]}
   );
   gpc1_1 gpc2974 (
      {stage1_36[82]},
      {stage2_36[36]}
   );
   gpc1_1 gpc2975 (
      {stage1_37[117]},
      {stage2_37[31]}
   );
   gpc1_1 gpc2976 (
      {stage1_37[118]},
      {stage2_37[32]}
   );
   gpc1_1 gpc2977 (
      {stage1_37[119]},
      {stage2_37[33]}
   );
   gpc1_1 gpc2978 (
      {stage1_37[120]},
      {stage2_37[34]}
   );
   gpc1_1 gpc2979 (
      {stage1_37[121]},
      {stage2_37[35]}
   );
   gpc1_1 gpc2980 (
      {stage1_37[122]},
      {stage2_37[36]}
   );
   gpc1_1 gpc2981 (
      {stage1_37[123]},
      {stage2_37[37]}
   );
   gpc1_1 gpc2982 (
      {stage1_37[124]},
      {stage2_37[38]}
   );
   gpc1_1 gpc2983 (
      {stage1_37[125]},
      {stage2_37[39]}
   );
   gpc1_1 gpc2984 (
      {stage1_37[126]},
      {stage2_37[40]}
   );
   gpc1_1 gpc2985 (
      {stage1_37[127]},
      {stage2_37[41]}
   );
   gpc1_1 gpc2986 (
      {stage1_39[64]},
      {stage2_39[30]}
   );
   gpc1_1 gpc2987 (
      {stage1_39[65]},
      {stage2_39[31]}
   );
   gpc1_1 gpc2988 (
      {stage1_39[66]},
      {stage2_39[32]}
   );
   gpc1_1 gpc2989 (
      {stage1_39[67]},
      {stage2_39[33]}
   );
   gpc1_1 gpc2990 (
      {stage1_40[72]},
      {stage2_40[31]}
   );
   gpc1_1 gpc2991 (
      {stage1_40[73]},
      {stage2_40[32]}
   );
   gpc1_1 gpc2992 (
      {stage1_40[74]},
      {stage2_40[33]}
   );
   gpc1_1 gpc2993 (
      {stage1_40[75]},
      {stage2_40[34]}
   );
   gpc1_1 gpc2994 (
      {stage1_40[76]},
      {stage2_40[35]}
   );
   gpc1_1 gpc2995 (
      {stage1_40[77]},
      {stage2_40[36]}
   );
   gpc1_1 gpc2996 (
      {stage1_40[78]},
      {stage2_40[37]}
   );
   gpc1_1 gpc2997 (
      {stage1_40[79]},
      {stage2_40[38]}
   );
   gpc1_1 gpc2998 (
      {stage1_40[80]},
      {stage2_40[39]}
   );
   gpc1_1 gpc2999 (
      {stage1_40[81]},
      {stage2_40[40]}
   );
   gpc1_1 gpc3000 (
      {stage1_41[48]},
      {stage2_41[30]}
   );
   gpc1_1 gpc3001 (
      {stage1_41[49]},
      {stage2_41[31]}
   );
   gpc1_1 gpc3002 (
      {stage1_41[50]},
      {stage2_41[32]}
   );
   gpc1_1 gpc3003 (
      {stage1_41[51]},
      {stage2_41[33]}
   );
   gpc1_1 gpc3004 (
      {stage1_41[52]},
      {stage2_41[34]}
   );
   gpc1_1 gpc3005 (
      {stage1_41[53]},
      {stage2_41[35]}
   );
   gpc1_1 gpc3006 (
      {stage1_41[54]},
      {stage2_41[36]}
   );
   gpc1_1 gpc3007 (
      {stage1_41[55]},
      {stage2_41[37]}
   );
   gpc1_1 gpc3008 (
      {stage1_41[56]},
      {stage2_41[38]}
   );
   gpc1_1 gpc3009 (
      {stage1_41[57]},
      {stage2_41[39]}
   );
   gpc1_1 gpc3010 (
      {stage1_41[58]},
      {stage2_41[40]}
   );
   gpc1_1 gpc3011 (
      {stage1_41[59]},
      {stage2_41[41]}
   );
   gpc1_1 gpc3012 (
      {stage1_41[60]},
      {stage2_41[42]}
   );
   gpc1_1 gpc3013 (
      {stage1_41[61]},
      {stage2_41[43]}
   );
   gpc1_1 gpc3014 (
      {stage1_41[62]},
      {stage2_41[44]}
   );
   gpc1_1 gpc3015 (
      {stage1_41[63]},
      {stage2_41[45]}
   );
   gpc1_1 gpc3016 (
      {stage1_41[64]},
      {stage2_41[46]}
   );
   gpc1_1 gpc3017 (
      {stage1_41[65]},
      {stage2_41[47]}
   );
   gpc1_1 gpc3018 (
      {stage1_41[66]},
      {stage2_41[48]}
   );
   gpc1_1 gpc3019 (
      {stage1_41[67]},
      {stage2_41[49]}
   );
   gpc1_1 gpc3020 (
      {stage1_41[68]},
      {stage2_41[50]}
   );
   gpc1_1 gpc3021 (
      {stage1_41[69]},
      {stage2_41[51]}
   );
   gpc1_1 gpc3022 (
      {stage1_41[70]},
      {stage2_41[52]}
   );
   gpc1_1 gpc3023 (
      {stage1_41[71]},
      {stage2_41[53]}
   );
   gpc1_1 gpc3024 (
      {stage1_41[72]},
      {stage2_41[54]}
   );
   gpc1_1 gpc3025 (
      {stage1_41[73]},
      {stage2_41[55]}
   );
   gpc1_1 gpc3026 (
      {stage1_42[54]},
      {stage2_42[20]}
   );
   gpc1_1 gpc3027 (
      {stage1_42[55]},
      {stage2_42[21]}
   );
   gpc1_1 gpc3028 (
      {stage1_42[56]},
      {stage2_42[22]}
   );
   gpc1_1 gpc3029 (
      {stage1_42[57]},
      {stage2_42[23]}
   );
   gpc1_1 gpc3030 (
      {stage1_42[58]},
      {stage2_42[24]}
   );
   gpc1_1 gpc3031 (
      {stage1_42[59]},
      {stage2_42[25]}
   );
   gpc1_1 gpc3032 (
      {stage1_42[60]},
      {stage2_42[26]}
   );
   gpc1_1 gpc3033 (
      {stage1_42[61]},
      {stage2_42[27]}
   );
   gpc1_1 gpc3034 (
      {stage1_42[62]},
      {stage2_42[28]}
   );
   gpc1_1 gpc3035 (
      {stage1_42[63]},
      {stage2_42[29]}
   );
   gpc1_1 gpc3036 (
      {stage1_42[64]},
      {stage2_42[30]}
   );
   gpc1_1 gpc3037 (
      {stage1_42[65]},
      {stage2_42[31]}
   );
   gpc1_1 gpc3038 (
      {stage1_42[66]},
      {stage2_42[32]}
   );
   gpc1_1 gpc3039 (
      {stage1_42[67]},
      {stage2_42[33]}
   );
   gpc1_1 gpc3040 (
      {stage1_42[68]},
      {stage2_42[34]}
   );
   gpc1_1 gpc3041 (
      {stage1_42[69]},
      {stage2_42[35]}
   );
   gpc1_1 gpc3042 (
      {stage1_42[70]},
      {stage2_42[36]}
   );
   gpc1_1 gpc3043 (
      {stage1_42[71]},
      {stage2_42[37]}
   );
   gpc1_1 gpc3044 (
      {stage1_42[72]},
      {stage2_42[38]}
   );
   gpc1_1 gpc3045 (
      {stage1_42[73]},
      {stage2_42[39]}
   );
   gpc1_1 gpc3046 (
      {stage1_42[74]},
      {stage2_42[40]}
   );
   gpc1_1 gpc3047 (
      {stage1_42[75]},
      {stage2_42[41]}
   );
   gpc1_1 gpc3048 (
      {stage1_42[76]},
      {stage2_42[42]}
   );
   gpc1_1 gpc3049 (
      {stage1_42[77]},
      {stage2_42[43]}
   );
   gpc1_1 gpc3050 (
      {stage1_42[78]},
      {stage2_42[44]}
   );
   gpc1_1 gpc3051 (
      {stage1_42[79]},
      {stage2_42[45]}
   );
   gpc1_1 gpc3052 (
      {stage1_42[80]},
      {stage2_42[46]}
   );
   gpc1_1 gpc3053 (
      {stage1_42[81]},
      {stage2_42[47]}
   );
   gpc1_1 gpc3054 (
      {stage1_42[82]},
      {stage2_42[48]}
   );
   gpc1_1 gpc3055 (
      {stage1_42[83]},
      {stage2_42[49]}
   );
   gpc1_1 gpc3056 (
      {stage1_42[84]},
      {stage2_42[50]}
   );
   gpc1_1 gpc3057 (
      {stage1_42[85]},
      {stage2_42[51]}
   );
   gpc1_1 gpc3058 (
      {stage1_42[86]},
      {stage2_42[52]}
   );
   gpc1_1 gpc3059 (
      {stage1_42[87]},
      {stage2_42[53]}
   );
   gpc1_1 gpc3060 (
      {stage1_42[88]},
      {stage2_42[54]}
   );
   gpc1_1 gpc3061 (
      {stage1_42[89]},
      {stage2_42[55]}
   );
   gpc1_1 gpc3062 (
      {stage1_42[90]},
      {stage2_42[56]}
   );
   gpc1_1 gpc3063 (
      {stage1_42[91]},
      {stage2_42[57]}
   );
   gpc1_1 gpc3064 (
      {stage1_42[92]},
      {stage2_42[58]}
   );
   gpc1_1 gpc3065 (
      {stage1_42[93]},
      {stage2_42[59]}
   );
   gpc1_1 gpc3066 (
      {stage1_42[94]},
      {stage2_42[60]}
   );
   gpc1_1 gpc3067 (
      {stage1_42[95]},
      {stage2_42[61]}
   );
   gpc1_1 gpc3068 (
      {stage1_43[114]},
      {stage2_43[28]}
   );
   gpc1_1 gpc3069 (
      {stage1_43[115]},
      {stage2_43[29]}
   );
   gpc1_1 gpc3070 (
      {stage1_43[116]},
      {stage2_43[30]}
   );
   gpc1_1 gpc3071 (
      {stage1_43[117]},
      {stage2_43[31]}
   );
   gpc1_1 gpc3072 (
      {stage1_43[118]},
      {stage2_43[32]}
   );
   gpc1_1 gpc3073 (
      {stage1_43[119]},
      {stage2_43[33]}
   );
   gpc1_1 gpc3074 (
      {stage1_43[120]},
      {stage2_43[34]}
   );
   gpc1_1 gpc3075 (
      {stage1_43[121]},
      {stage2_43[35]}
   );
   gpc1_1 gpc3076 (
      {stage1_43[122]},
      {stage2_43[36]}
   );
   gpc1_1 gpc3077 (
      {stage1_43[123]},
      {stage2_43[37]}
   );
   gpc1_1 gpc3078 (
      {stage1_43[124]},
      {stage2_43[38]}
   );
   gpc1_1 gpc3079 (
      {stage1_43[125]},
      {stage2_43[39]}
   );
   gpc1_1 gpc3080 (
      {stage1_43[126]},
      {stage2_43[40]}
   );
   gpc1_1 gpc3081 (
      {stage1_43[127]},
      {stage2_43[41]}
   );
   gpc1_1 gpc3082 (
      {stage1_43[128]},
      {stage2_43[42]}
   );
   gpc1_1 gpc3083 (
      {stage1_43[129]},
      {stage2_43[43]}
   );
   gpc1_1 gpc3084 (
      {stage1_43[130]},
      {stage2_43[44]}
   );
   gpc1_1 gpc3085 (
      {stage1_43[131]},
      {stage2_43[45]}
   );
   gpc1_1 gpc3086 (
      {stage1_43[132]},
      {stage2_43[46]}
   );
   gpc1_1 gpc3087 (
      {stage1_43[133]},
      {stage2_43[47]}
   );
   gpc1_1 gpc3088 (
      {stage1_43[134]},
      {stage2_43[48]}
   );
   gpc1_1 gpc3089 (
      {stage1_43[135]},
      {stage2_43[49]}
   );
   gpc1_1 gpc3090 (
      {stage1_43[136]},
      {stage2_43[50]}
   );
   gpc1_1 gpc3091 (
      {stage1_43[137]},
      {stage2_43[51]}
   );
   gpc1_1 gpc3092 (
      {stage1_44[10]},
      {stage2_44[30]}
   );
   gpc1_1 gpc3093 (
      {stage1_44[11]},
      {stage2_44[31]}
   );
   gpc1_1 gpc3094 (
      {stage1_44[12]},
      {stage2_44[32]}
   );
   gpc1_1 gpc3095 (
      {stage1_44[13]},
      {stage2_44[33]}
   );
   gpc1_1 gpc3096 (
      {stage1_44[14]},
      {stage2_44[34]}
   );
   gpc1_1 gpc3097 (
      {stage1_44[15]},
      {stage2_44[35]}
   );
   gpc1_1 gpc3098 (
      {stage1_44[16]},
      {stage2_44[36]}
   );
   gpc1_1 gpc3099 (
      {stage1_44[17]},
      {stage2_44[37]}
   );
   gpc1_1 gpc3100 (
      {stage1_44[18]},
      {stage2_44[38]}
   );
   gpc1_1 gpc3101 (
      {stage1_44[19]},
      {stage2_44[39]}
   );
   gpc1_1 gpc3102 (
      {stage1_44[20]},
      {stage2_44[40]}
   );
   gpc1_1 gpc3103 (
      {stage1_44[21]},
      {stage2_44[41]}
   );
   gpc1_1 gpc3104 (
      {stage1_44[22]},
      {stage2_44[42]}
   );
   gpc1_1 gpc3105 (
      {stage1_44[23]},
      {stage2_44[43]}
   );
   gpc1_1 gpc3106 (
      {stage1_44[24]},
      {stage2_44[44]}
   );
   gpc1_1 gpc3107 (
      {stage1_44[25]},
      {stage2_44[45]}
   );
   gpc1_1 gpc3108 (
      {stage1_44[26]},
      {stage2_44[46]}
   );
   gpc1_1 gpc3109 (
      {stage1_44[27]},
      {stage2_44[47]}
   );
   gpc1_1 gpc3110 (
      {stage1_44[28]},
      {stage2_44[48]}
   );
   gpc1_1 gpc3111 (
      {stage1_44[29]},
      {stage2_44[49]}
   );
   gpc1_1 gpc3112 (
      {stage1_44[30]},
      {stage2_44[50]}
   );
   gpc1_1 gpc3113 (
      {stage1_44[31]},
      {stage2_44[51]}
   );
   gpc1_1 gpc3114 (
      {stage1_44[32]},
      {stage2_44[52]}
   );
   gpc1_1 gpc3115 (
      {stage1_44[33]},
      {stage2_44[53]}
   );
   gpc1_1 gpc3116 (
      {stage1_44[34]},
      {stage2_44[54]}
   );
   gpc1_1 gpc3117 (
      {stage1_44[35]},
      {stage2_44[55]}
   );
   gpc1_1 gpc3118 (
      {stage1_44[36]},
      {stage2_44[56]}
   );
   gpc1_1 gpc3119 (
      {stage1_44[37]},
      {stage2_44[57]}
   );
   gpc1_1 gpc3120 (
      {stage1_44[38]},
      {stage2_44[58]}
   );
   gpc1_1 gpc3121 (
      {stage1_44[39]},
      {stage2_44[59]}
   );
   gpc1_1 gpc3122 (
      {stage1_44[40]},
      {stage2_44[60]}
   );
   gpc1_1 gpc3123 (
      {stage1_44[41]},
      {stage2_44[61]}
   );
   gpc1_1 gpc3124 (
      {stage1_44[42]},
      {stage2_44[62]}
   );
   gpc1_1 gpc3125 (
      {stage1_44[43]},
      {stage2_44[63]}
   );
   gpc1_1 gpc3126 (
      {stage1_44[44]},
      {stage2_44[64]}
   );
   gpc1_1 gpc3127 (
      {stage1_44[45]},
      {stage2_44[65]}
   );
   gpc1_1 gpc3128 (
      {stage1_45[92]},
      {stage2_45[25]}
   );
   gpc1_1 gpc3129 (
      {stage1_46[57]},
      {stage2_46[26]}
   );
   gpc1_1 gpc3130 (
      {stage1_46[58]},
      {stage2_46[27]}
   );
   gpc1_1 gpc3131 (
      {stage1_46[59]},
      {stage2_46[28]}
   );
   gpc1_1 gpc3132 (
      {stage1_46[60]},
      {stage2_46[29]}
   );
   gpc1_1 gpc3133 (
      {stage1_46[61]},
      {stage2_46[30]}
   );
   gpc1_1 gpc3134 (
      {stage1_46[62]},
      {stage2_46[31]}
   );
   gpc1_1 gpc3135 (
      {stage1_46[63]},
      {stage2_46[32]}
   );
   gpc1_1 gpc3136 (
      {stage1_47[39]},
      {stage2_47[27]}
   );
   gpc1_1 gpc3137 (
      {stage1_47[40]},
      {stage2_47[28]}
   );
   gpc1_1 gpc3138 (
      {stage1_47[41]},
      {stage2_47[29]}
   );
   gpc1_1 gpc3139 (
      {stage1_47[42]},
      {stage2_47[30]}
   );
   gpc1_1 gpc3140 (
      {stage1_47[43]},
      {stage2_47[31]}
   );
   gpc1_1 gpc3141 (
      {stage1_47[44]},
      {stage2_47[32]}
   );
   gpc1_1 gpc3142 (
      {stage1_47[45]},
      {stage2_47[33]}
   );
   gpc1_1 gpc3143 (
      {stage1_47[46]},
      {stage2_47[34]}
   );
   gpc1_1 gpc3144 (
      {stage1_47[47]},
      {stage2_47[35]}
   );
   gpc1_1 gpc3145 (
      {stage1_47[48]},
      {stage2_47[36]}
   );
   gpc1_1 gpc3146 (
      {stage1_47[49]},
      {stage2_47[37]}
   );
   gpc1_1 gpc3147 (
      {stage1_47[50]},
      {stage2_47[38]}
   );
   gpc1_1 gpc3148 (
      {stage1_47[51]},
      {stage2_47[39]}
   );
   gpc1_1 gpc3149 (
      {stage1_47[52]},
      {stage2_47[40]}
   );
   gpc1_1 gpc3150 (
      {stage1_47[53]},
      {stage2_47[41]}
   );
   gpc1_1 gpc3151 (
      {stage1_47[54]},
      {stage2_47[42]}
   );
   gpc1_1 gpc3152 (
      {stage1_47[55]},
      {stage2_47[43]}
   );
   gpc1_1 gpc3153 (
      {stage1_47[56]},
      {stage2_47[44]}
   );
   gpc1_1 gpc3154 (
      {stage1_47[57]},
      {stage2_47[45]}
   );
   gpc1_1 gpc3155 (
      {stage1_48[66]},
      {stage2_48[18]}
   );
   gpc1_1 gpc3156 (
      {stage1_48[67]},
      {stage2_48[19]}
   );
   gpc1_1 gpc3157 (
      {stage1_48[68]},
      {stage2_48[20]}
   );
   gpc1_1 gpc3158 (
      {stage1_48[69]},
      {stage2_48[21]}
   );
   gpc1_1 gpc3159 (
      {stage1_48[70]},
      {stage2_48[22]}
   );
   gpc1_1 gpc3160 (
      {stage1_48[71]},
      {stage2_48[23]}
   );
   gpc1_1 gpc3161 (
      {stage1_49[78]},
      {stage2_49[28]}
   );
   gpc1_1 gpc3162 (
      {stage1_49[79]},
      {stage2_49[29]}
   );
   gpc1_1 gpc3163 (
      {stage1_49[80]},
      {stage2_49[30]}
   );
   gpc1_1 gpc3164 (
      {stage1_49[81]},
      {stage2_49[31]}
   );
   gpc1_1 gpc3165 (
      {stage1_49[82]},
      {stage2_49[32]}
   );
   gpc1_1 gpc3166 (
      {stage1_49[83]},
      {stage2_49[33]}
   );
   gpc1_1 gpc3167 (
      {stage1_49[84]},
      {stage2_49[34]}
   );
   gpc1_1 gpc3168 (
      {stage1_49[85]},
      {stage2_49[35]}
   );
   gpc1_1 gpc3169 (
      {stage1_49[86]},
      {stage2_49[36]}
   );
   gpc1_1 gpc3170 (
      {stage1_50[47]},
      {stage2_50[30]}
   );
   gpc1_1 gpc3171 (
      {stage1_50[48]},
      {stage2_50[31]}
   );
   gpc1_1 gpc3172 (
      {stage1_50[49]},
      {stage2_50[32]}
   );
   gpc1_1 gpc3173 (
      {stage1_50[50]},
      {stage2_50[33]}
   );
   gpc1_1 gpc3174 (
      {stage1_50[51]},
      {stage2_50[34]}
   );
   gpc1_1 gpc3175 (
      {stage1_50[52]},
      {stage2_50[35]}
   );
   gpc1_1 gpc3176 (
      {stage1_50[53]},
      {stage2_50[36]}
   );
   gpc1_1 gpc3177 (
      {stage1_50[54]},
      {stage2_50[37]}
   );
   gpc1_1 gpc3178 (
      {stage1_50[55]},
      {stage2_50[38]}
   );
   gpc1_1 gpc3179 (
      {stage1_50[56]},
      {stage2_50[39]}
   );
   gpc1_1 gpc3180 (
      {stage1_50[57]},
      {stage2_50[40]}
   );
   gpc1_1 gpc3181 (
      {stage1_51[93]},
      {stage2_51[24]}
   );
   gpc1_1 gpc3182 (
      {stage1_52[73]},
      {stage2_52[30]}
   );
   gpc1_1 gpc3183 (
      {stage1_52[74]},
      {stage2_52[31]}
   );
   gpc1_1 gpc3184 (
      {stage1_52[75]},
      {stage2_52[32]}
   );
   gpc1_1 gpc3185 (
      {stage1_52[76]},
      {stage2_52[33]}
   );
   gpc1_1 gpc3186 (
      {stage1_53[48]},
      {stage2_53[33]}
   );
   gpc1_1 gpc3187 (
      {stage1_53[49]},
      {stage2_53[34]}
   );
   gpc1_1 gpc3188 (
      {stage1_53[50]},
      {stage2_53[35]}
   );
   gpc1_1 gpc3189 (
      {stage1_53[51]},
      {stage2_53[36]}
   );
   gpc1_1 gpc3190 (
      {stage1_53[52]},
      {stage2_53[37]}
   );
   gpc1_1 gpc3191 (
      {stage1_53[53]},
      {stage2_53[38]}
   );
   gpc1_1 gpc3192 (
      {stage1_53[54]},
      {stage2_53[39]}
   );
   gpc1_1 gpc3193 (
      {stage1_53[55]},
      {stage2_53[40]}
   );
   gpc1_1 gpc3194 (
      {stage1_53[56]},
      {stage2_53[41]}
   );
   gpc1_1 gpc3195 (
      {stage1_53[57]},
      {stage2_53[42]}
   );
   gpc1_1 gpc3196 (
      {stage1_53[58]},
      {stage2_53[43]}
   );
   gpc1_1 gpc3197 (
      {stage1_53[59]},
      {stage2_53[44]}
   );
   gpc1_1 gpc3198 (
      {stage1_53[60]},
      {stage2_53[45]}
   );
   gpc1_1 gpc3199 (
      {stage1_53[61]},
      {stage2_53[46]}
   );
   gpc1_1 gpc3200 (
      {stage1_53[62]},
      {stage2_53[47]}
   );
   gpc1_1 gpc3201 (
      {stage1_53[63]},
      {stage2_53[48]}
   );
   gpc1_1 gpc3202 (
      {stage1_53[64]},
      {stage2_53[49]}
   );
   gpc1_1 gpc3203 (
      {stage1_53[65]},
      {stage2_53[50]}
   );
   gpc1_1 gpc3204 (
      {stage1_54[52]},
      {stage2_54[22]}
   );
   gpc1_1 gpc3205 (
      {stage1_54[53]},
      {stage2_54[23]}
   );
   gpc1_1 gpc3206 (
      {stage1_54[54]},
      {stage2_54[24]}
   );
   gpc1_1 gpc3207 (
      {stage1_54[55]},
      {stage2_54[25]}
   );
   gpc1_1 gpc3208 (
      {stage1_54[56]},
      {stage2_54[26]}
   );
   gpc1_1 gpc3209 (
      {stage1_54[57]},
      {stage2_54[27]}
   );
   gpc1_1 gpc3210 (
      {stage1_55[88]},
      {stage2_55[28]}
   );
   gpc1_1 gpc3211 (
      {stage1_55[89]},
      {stage2_55[29]}
   );
   gpc1_1 gpc3212 (
      {stage1_55[90]},
      {stage2_55[30]}
   );
   gpc1_1 gpc3213 (
      {stage1_55[91]},
      {stage2_55[31]}
   );
   gpc1_1 gpc3214 (
      {stage1_55[92]},
      {stage2_55[32]}
   );
   gpc1_1 gpc3215 (
      {stage1_55[93]},
      {stage2_55[33]}
   );
   gpc1_1 gpc3216 (
      {stage1_55[94]},
      {stage2_55[34]}
   );
   gpc1_1 gpc3217 (
      {stage1_55[95]},
      {stage2_55[35]}
   );
   gpc1_1 gpc3218 (
      {stage1_55[96]},
      {stage2_55[36]}
   );
   gpc1_1 gpc3219 (
      {stage1_55[97]},
      {stage2_55[37]}
   );
   gpc1_1 gpc3220 (
      {stage1_56[58]},
      {stage2_56[31]}
   );
   gpc1_1 gpc3221 (
      {stage1_56[59]},
      {stage2_56[32]}
   );
   gpc1_1 gpc3222 (
      {stage1_56[60]},
      {stage2_56[33]}
   );
   gpc1_1 gpc3223 (
      {stage1_56[61]},
      {stage2_56[34]}
   );
   gpc1_1 gpc3224 (
      {stage1_56[62]},
      {stage2_56[35]}
   );
   gpc1_1 gpc3225 (
      {stage1_56[63]},
      {stage2_56[36]}
   );
   gpc1_1 gpc3226 (
      {stage1_56[64]},
      {stage2_56[37]}
   );
   gpc1_1 gpc3227 (
      {stage1_56[65]},
      {stage2_56[38]}
   );
   gpc1_1 gpc3228 (
      {stage1_56[66]},
      {stage2_56[39]}
   );
   gpc1_1 gpc3229 (
      {stage1_56[67]},
      {stage2_56[40]}
   );
   gpc1_1 gpc3230 (
      {stage1_56[68]},
      {stage2_56[41]}
   );
   gpc1_1 gpc3231 (
      {stage1_56[69]},
      {stage2_56[42]}
   );
   gpc1_1 gpc3232 (
      {stage1_56[70]},
      {stage2_56[43]}
   );
   gpc1_1 gpc3233 (
      {stage1_56[71]},
      {stage2_56[44]}
   );
   gpc1_1 gpc3234 (
      {stage1_56[72]},
      {stage2_56[45]}
   );
   gpc1_1 gpc3235 (
      {stage1_56[73]},
      {stage2_56[46]}
   );
   gpc1_1 gpc3236 (
      {stage1_56[74]},
      {stage2_56[47]}
   );
   gpc1_1 gpc3237 (
      {stage1_56[75]},
      {stage2_56[48]}
   );
   gpc1_1 gpc3238 (
      {stage1_56[76]},
      {stage2_56[49]}
   );
   gpc1_1 gpc3239 (
      {stage1_56[77]},
      {stage2_56[50]}
   );
   gpc1_1 gpc3240 (
      {stage1_56[78]},
      {stage2_56[51]}
   );
   gpc1_1 gpc3241 (
      {stage1_56[79]},
      {stage2_56[52]}
   );
   gpc1_1 gpc3242 (
      {stage1_57[66]},
      {stage2_57[24]}
   );
   gpc1_1 gpc3243 (
      {stage1_57[67]},
      {stage2_57[25]}
   );
   gpc1_1 gpc3244 (
      {stage1_57[68]},
      {stage2_57[26]}
   );
   gpc1_1 gpc3245 (
      {stage1_57[69]},
      {stage2_57[27]}
   );
   gpc1_1 gpc3246 (
      {stage1_57[70]},
      {stage2_57[28]}
   );
   gpc1_1 gpc3247 (
      {stage1_57[71]},
      {stage2_57[29]}
   );
   gpc1_1 gpc3248 (
      {stage1_58[65]},
      {stage2_58[24]}
   );
   gpc1_1 gpc3249 (
      {stage1_58[66]},
      {stage2_58[25]}
   );
   gpc1_1 gpc3250 (
      {stage1_58[67]},
      {stage2_58[26]}
   );
   gpc1_1 gpc3251 (
      {stage1_58[68]},
      {stage2_58[27]}
   );
   gpc1_1 gpc3252 (
      {stage1_58[69]},
      {stage2_58[28]}
   );
   gpc1_1 gpc3253 (
      {stage1_58[70]},
      {stage2_58[29]}
   );
   gpc1_1 gpc3254 (
      {stage1_58[71]},
      {stage2_58[30]}
   );
   gpc1_1 gpc3255 (
      {stage1_58[72]},
      {stage2_58[31]}
   );
   gpc1_1 gpc3256 (
      {stage1_58[73]},
      {stage2_58[32]}
   );
   gpc1_1 gpc3257 (
      {stage1_59[25]},
      {stage2_59[26]}
   );
   gpc1_1 gpc3258 (
      {stage1_59[26]},
      {stage2_59[27]}
   );
   gpc1_1 gpc3259 (
      {stage1_59[27]},
      {stage2_59[28]}
   );
   gpc1_1 gpc3260 (
      {stage1_59[28]},
      {stage2_59[29]}
   );
   gpc1_1 gpc3261 (
      {stage1_59[29]},
      {stage2_59[30]}
   );
   gpc1_1 gpc3262 (
      {stage1_59[30]},
      {stage2_59[31]}
   );
   gpc1_1 gpc3263 (
      {stage1_59[31]},
      {stage2_59[32]}
   );
   gpc1_1 gpc3264 (
      {stage1_59[32]},
      {stage2_59[33]}
   );
   gpc1_1 gpc3265 (
      {stage1_59[33]},
      {stage2_59[34]}
   );
   gpc1_1 gpc3266 (
      {stage1_59[34]},
      {stage2_59[35]}
   );
   gpc1_1 gpc3267 (
      {stage1_59[35]},
      {stage2_59[36]}
   );
   gpc1_1 gpc3268 (
      {stage1_59[36]},
      {stage2_59[37]}
   );
   gpc1_1 gpc3269 (
      {stage1_59[37]},
      {stage2_59[38]}
   );
   gpc1_1 gpc3270 (
      {stage1_59[38]},
      {stage2_59[39]}
   );
   gpc1_1 gpc3271 (
      {stage1_59[39]},
      {stage2_59[40]}
   );
   gpc1_1 gpc3272 (
      {stage1_59[40]},
      {stage2_59[41]}
   );
   gpc1_1 gpc3273 (
      {stage1_59[41]},
      {stage2_59[42]}
   );
   gpc1_1 gpc3274 (
      {stage1_59[42]},
      {stage2_59[43]}
   );
   gpc1_1 gpc3275 (
      {stage1_59[43]},
      {stage2_59[44]}
   );
   gpc1_1 gpc3276 (
      {stage1_59[44]},
      {stage2_59[45]}
   );
   gpc1_1 gpc3277 (
      {stage1_59[45]},
      {stage2_59[46]}
   );
   gpc1_1 gpc3278 (
      {stage1_59[46]},
      {stage2_59[47]}
   );
   gpc1_1 gpc3279 (
      {stage1_59[47]},
      {stage2_59[48]}
   );
   gpc1_1 gpc3280 (
      {stage1_59[48]},
      {stage2_59[49]}
   );
   gpc1_1 gpc3281 (
      {stage1_59[49]},
      {stage2_59[50]}
   );
   gpc1_1 gpc3282 (
      {stage1_59[50]},
      {stage2_59[51]}
   );
   gpc1_1 gpc3283 (
      {stage1_59[51]},
      {stage2_59[52]}
   );
   gpc1_1 gpc3284 (
      {stage1_59[52]},
      {stage2_59[53]}
   );
   gpc1_1 gpc3285 (
      {stage1_59[53]},
      {stage2_59[54]}
   );
   gpc1_1 gpc3286 (
      {stage1_59[54]},
      {stage2_59[55]}
   );
   gpc1_1 gpc3287 (
      {stage1_59[55]},
      {stage2_59[56]}
   );
   gpc1_1 gpc3288 (
      {stage1_59[56]},
      {stage2_59[57]}
   );
   gpc1_1 gpc3289 (
      {stage1_59[57]},
      {stage2_59[58]}
   );
   gpc1_1 gpc3290 (
      {stage1_59[58]},
      {stage2_59[59]}
   );
   gpc1_1 gpc3291 (
      {stage1_59[59]},
      {stage2_59[60]}
   );
   gpc1_1 gpc3292 (
      {stage1_59[60]},
      {stage2_59[61]}
   );
   gpc1_1 gpc3293 (
      {stage1_59[61]},
      {stage2_59[62]}
   );
   gpc1_1 gpc3294 (
      {stage1_59[62]},
      {stage2_59[63]}
   );
   gpc1_1 gpc3295 (
      {stage1_59[63]},
      {stage2_59[64]}
   );
   gpc1_1 gpc3296 (
      {stage1_59[64]},
      {stage2_59[65]}
   );
   gpc1_1 gpc3297 (
      {stage1_59[65]},
      {stage2_59[66]}
   );
   gpc1_1 gpc3298 (
      {stage1_59[66]},
      {stage2_59[67]}
   );
   gpc1_1 gpc3299 (
      {stage1_59[67]},
      {stage2_59[68]}
   );
   gpc1_1 gpc3300 (
      {stage1_59[68]},
      {stage2_59[69]}
   );
   gpc1_1 gpc3301 (
      {stage1_59[69]},
      {stage2_59[70]}
   );
   gpc1_1 gpc3302 (
      {stage1_59[70]},
      {stage2_59[71]}
   );
   gpc1_1 gpc3303 (
      {stage1_59[71]},
      {stage2_59[72]}
   );
   gpc1_1 gpc3304 (
      {stage1_59[72]},
      {stage2_59[73]}
   );
   gpc1_1 gpc3305 (
      {stage1_59[73]},
      {stage2_59[74]}
   );
   gpc1_1 gpc3306 (
      {stage1_59[74]},
      {stage2_59[75]}
   );
   gpc1_1 gpc3307 (
      {stage1_59[75]},
      {stage2_59[76]}
   );
   gpc1_1 gpc3308 (
      {stage1_59[76]},
      {stage2_59[77]}
   );
   gpc1_1 gpc3309 (
      {stage1_59[77]},
      {stage2_59[78]}
   );
   gpc1_1 gpc3310 (
      {stage1_59[78]},
      {stage2_59[79]}
   );
   gpc1_1 gpc3311 (
      {stage1_59[79]},
      {stage2_59[80]}
   );
   gpc1_1 gpc3312 (
      {stage1_60[66]},
      {stage2_60[21]}
   );
   gpc1_1 gpc3313 (
      {stage1_61[42]},
      {stage2_61[18]}
   );
   gpc1_1 gpc3314 (
      {stage1_61[43]},
      {stage2_61[19]}
   );
   gpc1_1 gpc3315 (
      {stage1_61[44]},
      {stage2_61[20]}
   );
   gpc1_1 gpc3316 (
      {stage1_61[45]},
      {stage2_61[21]}
   );
   gpc1_1 gpc3317 (
      {stage1_61[46]},
      {stage2_61[22]}
   );
   gpc1_1 gpc3318 (
      {stage1_61[47]},
      {stage2_61[23]}
   );
   gpc1_1 gpc3319 (
      {stage1_61[48]},
      {stage2_61[24]}
   );
   gpc1_1 gpc3320 (
      {stage1_61[49]},
      {stage2_61[25]}
   );
   gpc1_1 gpc3321 (
      {stage1_61[50]},
      {stage2_61[26]}
   );
   gpc1_1 gpc3322 (
      {stage1_61[51]},
      {stage2_61[27]}
   );
   gpc1_1 gpc3323 (
      {stage1_61[52]},
      {stage2_61[28]}
   );
   gpc1_1 gpc3324 (
      {stage1_61[53]},
      {stage2_61[29]}
   );
   gpc1_1 gpc3325 (
      {stage1_61[54]},
      {stage2_61[30]}
   );
   gpc1_1 gpc3326 (
      {stage1_61[55]},
      {stage2_61[31]}
   );
   gpc1_1 gpc3327 (
      {stage1_61[56]},
      {stage2_61[32]}
   );
   gpc1_1 gpc3328 (
      {stage1_61[57]},
      {stage2_61[33]}
   );
   gpc1_1 gpc3329 (
      {stage1_61[58]},
      {stage2_61[34]}
   );
   gpc1_1 gpc3330 (
      {stage1_61[59]},
      {stage2_61[35]}
   );
   gpc1_1 gpc3331 (
      {stage1_61[60]},
      {stage2_61[36]}
   );
   gpc1_1 gpc3332 (
      {stage1_61[61]},
      {stage2_61[37]}
   );
   gpc1_1 gpc3333 (
      {stage1_61[62]},
      {stage2_61[38]}
   );
   gpc1_1 gpc3334 (
      {stage1_61[63]},
      {stage2_61[39]}
   );
   gpc1_1 gpc3335 (
      {stage1_61[64]},
      {stage2_61[40]}
   );
   gpc1_1 gpc3336 (
      {stage1_61[65]},
      {stage2_61[41]}
   );
   gpc1_1 gpc3337 (
      {stage1_61[66]},
      {stage2_61[42]}
   );
   gpc1_1 gpc3338 (
      {stage1_61[67]},
      {stage2_61[43]}
   );
   gpc1_1 gpc3339 (
      {stage1_61[68]},
      {stage2_61[44]}
   );
   gpc1_1 gpc3340 (
      {stage1_61[69]},
      {stage2_61[45]}
   );
   gpc1_1 gpc3341 (
      {stage1_61[70]},
      {stage2_61[46]}
   );
   gpc1_1 gpc3342 (
      {stage1_61[71]},
      {stage2_61[47]}
   );
   gpc1_1 gpc3343 (
      {stage1_61[72]},
      {stage2_61[48]}
   );
   gpc1_1 gpc3344 (
      {stage1_61[73]},
      {stage2_61[49]}
   );
   gpc1_1 gpc3345 (
      {stage1_61[74]},
      {stage2_61[50]}
   );
   gpc1_1 gpc3346 (
      {stage1_61[75]},
      {stage2_61[51]}
   );
   gpc1_1 gpc3347 (
      {stage1_61[76]},
      {stage2_61[52]}
   );
   gpc1_1 gpc3348 (
      {stage1_61[77]},
      {stage2_61[53]}
   );
   gpc1_1 gpc3349 (
      {stage1_61[78]},
      {stage2_61[54]}
   );
   gpc1_1 gpc3350 (
      {stage1_61[79]},
      {stage2_61[55]}
   );
   gpc1_1 gpc3351 (
      {stage1_61[80]},
      {stage2_61[56]}
   );
   gpc1_1 gpc3352 (
      {stage1_61[81]},
      {stage2_61[57]}
   );
   gpc1_1 gpc3353 (
      {stage1_61[82]},
      {stage2_61[58]}
   );
   gpc1_1 gpc3354 (
      {stage1_61[83]},
      {stage2_61[59]}
   );
   gpc1_1 gpc3355 (
      {stage1_61[84]},
      {stage2_61[60]}
   );
   gpc1_1 gpc3356 (
      {stage1_61[85]},
      {stage2_61[61]}
   );
   gpc1_1 gpc3357 (
      {stage1_61[86]},
      {stage2_61[62]}
   );
   gpc1_1 gpc3358 (
      {stage1_61[87]},
      {stage2_61[63]}
   );
   gpc1_1 gpc3359 (
      {stage1_61[88]},
      {stage2_61[64]}
   );
   gpc1_1 gpc3360 (
      {stage1_61[89]},
      {stage2_61[65]}
   );
   gpc1_1 gpc3361 (
      {stage1_61[90]},
      {stage2_61[66]}
   );
   gpc1_1 gpc3362 (
      {stage1_62[78]},
      {stage2_62[26]}
   );
   gpc1_1 gpc3363 (
      {stage1_62[79]},
      {stage2_62[27]}
   );
   gpc1_1 gpc3364 (
      {stage1_62[80]},
      {stage2_62[28]}
   );
   gpc1_1 gpc3365 (
      {stage1_62[81]},
      {stage2_62[29]}
   );
   gpc1_1 gpc3366 (
      {stage1_62[82]},
      {stage2_62[30]}
   );
   gpc1_1 gpc3367 (
      {stage1_62[83]},
      {stage2_62[31]}
   );
   gpc1_1 gpc3368 (
      {stage1_62[84]},
      {stage2_62[32]}
   );
   gpc1_1 gpc3369 (
      {stage1_62[85]},
      {stage2_62[33]}
   );
   gpc1_1 gpc3370 (
      {stage1_62[86]},
      {stage2_62[34]}
   );
   gpc1_1 gpc3371 (
      {stage1_63[48]},
      {stage2_63[23]}
   );
   gpc1_1 gpc3372 (
      {stage1_63[49]},
      {stage2_63[24]}
   );
   gpc1_1 gpc3373 (
      {stage1_63[50]},
      {stage2_63[25]}
   );
   gpc1_1 gpc3374 (
      {stage1_63[51]},
      {stage2_63[26]}
   );
   gpc1_1 gpc3375 (
      {stage1_63[52]},
      {stage2_63[27]}
   );
   gpc1_1 gpc3376 (
      {stage1_63[53]},
      {stage2_63[28]}
   );
   gpc1_1 gpc3377 (
      {stage1_63[54]},
      {stage2_63[29]}
   );
   gpc1_1 gpc3378 (
      {stage1_63[55]},
      {stage2_63[30]}
   );
   gpc1_1 gpc3379 (
      {stage1_63[56]},
      {stage2_63[31]}
   );
   gpc1_1 gpc3380 (
      {stage1_63[57]},
      {stage2_63[32]}
   );
   gpc1_1 gpc3381 (
      {stage1_63[58]},
      {stage2_63[33]}
   );
   gpc1_1 gpc3382 (
      {stage1_63[59]},
      {stage2_63[34]}
   );
   gpc1_1 gpc3383 (
      {stage1_63[60]},
      {stage2_63[35]}
   );
   gpc1_1 gpc3384 (
      {stage1_63[61]},
      {stage2_63[36]}
   );
   gpc1_1 gpc3385 (
      {stage1_63[62]},
      {stage2_63[37]}
   );
   gpc1_1 gpc3386 (
      {stage1_64[18]},
      {stage2_64[19]}
   );
   gpc1_1 gpc3387 (
      {stage1_64[19]},
      {stage2_64[20]}
   );
   gpc1_1 gpc3388 (
      {stage1_64[20]},
      {stage2_64[21]}
   );
   gpc1_1 gpc3389 (
      {stage1_64[21]},
      {stage2_64[22]}
   );
   gpc1_1 gpc3390 (
      {stage1_64[22]},
      {stage2_64[23]}
   );
   gpc1_1 gpc3391 (
      {stage1_64[23]},
      {stage2_64[24]}
   );
   gpc1_1 gpc3392 (
      {stage1_64[24]},
      {stage2_64[25]}
   );
   gpc1_1 gpc3393 (
      {stage1_64[25]},
      {stage2_64[26]}
   );
   gpc1_1 gpc3394 (
      {stage1_64[26]},
      {stage2_64[27]}
   );
   gpc1_1 gpc3395 (
      {stage1_64[27]},
      {stage2_64[28]}
   );
   gpc1_1 gpc3396 (
      {stage1_64[28]},
      {stage2_64[29]}
   );
   gpc1_1 gpc3397 (
      {stage1_64[29]},
      {stage2_64[30]}
   );
   gpc1_1 gpc3398 (
      {stage1_64[30]},
      {stage2_64[31]}
   );
   gpc1_1 gpc3399 (
      {stage1_64[31]},
      {stage2_64[32]}
   );
   gpc1_1 gpc3400 (
      {stage1_64[32]},
      {stage2_64[33]}
   );
   gpc1_1 gpc3401 (
      {stage1_64[33]},
      {stage2_64[34]}
   );
   gpc1_1 gpc3402 (
      {stage1_64[34]},
      {stage2_64[35]}
   );
   gpc1_1 gpc3403 (
      {stage1_64[35]},
      {stage2_64[36]}
   );
   gpc1_1 gpc3404 (
      {stage1_64[36]},
      {stage2_64[37]}
   );
   gpc1_1 gpc3405 (
      {stage1_64[37]},
      {stage2_64[38]}
   );
   gpc1_1 gpc3406 (
      {stage1_64[38]},
      {stage2_64[39]}
   );
   gpc1_1 gpc3407 (
      {stage1_64[39]},
      {stage2_64[40]}
   );
   gpc1_1 gpc3408 (
      {stage1_64[40]},
      {stage2_64[41]}
   );
   gpc1_1 gpc3409 (
      {stage1_64[41]},
      {stage2_64[42]}
   );
   gpc1_1 gpc3410 (
      {stage1_64[42]},
      {stage2_64[43]}
   );
   gpc1_1 gpc3411 (
      {stage1_64[43]},
      {stage2_64[44]}
   );
   gpc1_1 gpc3412 (
      {stage1_64[44]},
      {stage2_64[45]}
   );
   gpc1163_5 gpc3413 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc3414 (
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc606_5 gpc3415 (
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[1],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc606_5 gpc3416 (
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[2],stage3_4[3],stage3_3[3],stage3_2[3]}
   );
   gpc615_5 gpc3417 (
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage2_3[1]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[3],stage3_4[4],stage3_3[4],stage3_2[4]}
   );
   gpc615_5 gpc3418 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28]},
      {stage2_3[2]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[4],stage3_4[5],stage3_3[5],stage3_2[5]}
   );
   gpc615_5 gpc3419 (
      {stage2_2[29], stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33]},
      {stage2_3[3]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[5],stage3_4[6],stage3_3[6],stage3_2[6]}
   );
   gpc615_5 gpc3420 (
      {stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7], stage2_3[8]},
      {stage2_4[36]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[6],stage3_5[6],stage3_4[7],stage3_3[7]}
   );
   gpc615_5 gpc3421 (
      {stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage2_4[37]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[7],stage3_5[7],stage3_4[8],stage3_3[8]}
   );
   gpc615_5 gpc3422 (
      {stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage2_4[38]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[8],stage3_5[8],stage3_4[9],stage3_3[9]}
   );
   gpc606_5 gpc3423 (
      {stage2_4[39], stage2_4[40], stage2_4[41], stage2_4[42], stage2_4[43], stage2_4[44]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[9],stage3_5[9],stage3_4[10]}
   );
   gpc606_5 gpc3424 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[1],stage3_7[4],stage3_6[10],stage3_5[10]}
   );
   gpc606_5 gpc3425 (
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[2],stage3_7[5],stage3_6[11],stage3_5[11]}
   );
   gpc606_5 gpc3426 (
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[2],stage3_8[3],stage3_7[6],stage3_6[12]}
   );
   gpc606_5 gpc3427 (
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[3],stage3_8[4],stage3_7[7],stage3_6[13]}
   );
   gpc606_5 gpc3428 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[4],stage3_8[5],stage3_7[8],stage3_6[14]}
   );
   gpc207_4 gpc3429 (
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18]},
      {stage2_9[0], stage2_9[1]},
      {stage3_10[3],stage3_9[5],stage3_8[6],stage3_7[9]}
   );
   gpc207_4 gpc3430 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23], stage2_7[24], stage2_7[25]},
      {stage2_9[2], stage2_9[3]},
      {stage3_10[4],stage3_9[6],stage3_8[7],stage3_7[10]}
   );
   gpc606_5 gpc3431 (
      {stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31]},
      {stage2_9[4], stage2_9[5], stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9]},
      {stage3_11[0],stage3_10[5],stage3_9[7],stage3_8[8],stage3_7[11]}
   );
   gpc615_5 gpc3432 (
      {stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_8[18]},
      {stage2_9[10], stage2_9[11], stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15]},
      {stage3_11[1],stage3_10[6],stage3_9[8],stage3_8[9],stage3_7[12]}
   );
   gpc606_5 gpc3433 (
      {stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[7],stage3_9[9],stage3_8[10]}
   );
   gpc606_5 gpc3434 (
      {stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[3],stage3_10[8],stage3_9[10],stage3_8[11]}
   );
   gpc606_5 gpc3435 (
      {stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35], stage2_8[36]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[4],stage3_10[9],stage3_9[11],stage3_8[12]}
   );
   gpc606_5 gpc3436 (
      {stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41], stage2_8[42]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[5],stage3_10[10],stage3_9[12],stage3_8[13]}
   );
   gpc606_5 gpc3437 (
      {stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47], stage2_8[48]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[6],stage3_10[11],stage3_9[13],stage3_8[14]}
   );
   gpc606_5 gpc3438 (
      {stage2_8[49], stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53], stage2_8[54]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[7],stage3_10[12],stage3_9[14],stage3_8[15]}
   );
   gpc606_5 gpc3439 (
      {stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59], stage2_8[60]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], 1'b0},
      {stage3_12[6],stage3_11[8],stage3_10[13],stage3_9[15],stage3_8[16]}
   );
   gpc606_5 gpc3440 (
      {stage2_9[16], stage2_9[17], stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[7],stage3_11[9],stage3_10[14],stage3_9[16]}
   );
   gpc606_5 gpc3441 (
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[1],stage3_12[8],stage3_11[10]}
   );
   gpc606_5 gpc3442 (
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[2],stage3_12[9],stage3_11[11]}
   );
   gpc606_5 gpc3443 (
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[2],stage3_13[3],stage3_12[10],stage3_11[12]}
   );
   gpc606_5 gpc3444 (
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[3],stage3_13[4],stage3_12[11],stage3_11[13]}
   );
   gpc606_5 gpc3445 (
      {stage2_11[30], stage2_11[31], stage2_11[32], stage2_11[33], stage2_11[34], stage2_11[35]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[4],stage3_13[5],stage3_12[12],stage3_11[14]}
   );
   gpc606_5 gpc3446 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[5],stage3_14[5],stage3_13[6],stage3_12[13]}
   );
   gpc606_5 gpc3447 (
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[6],stage3_14[6],stage3_13[7],stage3_12[14]}
   );
   gpc606_5 gpc3448 (
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[7],stage3_14[7],stage3_13[8],stage3_12[15]}
   );
   gpc606_5 gpc3449 (
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[8],stage3_14[8],stage3_13[9],stage3_12[16]}
   );
   gpc606_5 gpc3450 (
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[9],stage3_14[9],stage3_13[10]}
   );
   gpc615_5 gpc3451 (
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28]},
      {stage2_15[6]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[1],stage3_16[5],stage3_15[10],stage3_14[10]}
   );
   gpc615_5 gpc3452 (
      {stage2_14[29], stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33]},
      {stage2_15[7]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[2],stage3_16[6],stage3_15[11],stage3_14[11]}
   );
   gpc615_5 gpc3453 (
      {stage2_14[34], stage2_14[35], stage2_14[36], stage2_14[37], stage2_14[38]},
      {stage2_15[8]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[3],stage3_16[7],stage3_15[12],stage3_14[12]}
   );
   gpc615_5 gpc3454 (
      {stage2_14[39], stage2_14[40], stage2_14[41], stage2_14[42], stage2_14[43]},
      {stage2_15[9]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[4],stage3_16[8],stage3_15[13],stage3_14[13]}
   );
   gpc615_5 gpc3455 (
      {stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47], stage2_14[48]},
      {stage2_15[10]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[5],stage3_16[9],stage3_15[14],stage3_14[14]}
   );
   gpc615_5 gpc3456 (
      {stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage2_15[11]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[6],stage3_16[10],stage3_15[15],stage3_14[15]}
   );
   gpc615_5 gpc3457 (
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16]},
      {stage2_16[36]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[6],stage3_17[7],stage3_16[11],stage3_15[16]}
   );
   gpc606_5 gpc3458 (
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[1],stage3_18[7],stage3_17[8]}
   );
   gpc606_5 gpc3459 (
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[1],stage3_19[2],stage3_18[8],stage3_17[9]}
   );
   gpc606_5 gpc3460 (
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage3_21[2],stage3_20[2],stage3_19[3],stage3_18[9],stage3_17[10]}
   );
   gpc606_5 gpc3461 (
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage2_19[18], stage2_19[19], stage2_19[20], stage2_19[21], stage2_19[22], stage2_19[23]},
      {stage3_21[3],stage3_20[3],stage3_19[4],stage3_18[10],stage3_17[11]}
   );
   gpc606_5 gpc3462 (
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage2_19[24], stage2_19[25], stage2_19[26], stage2_19[27], stage2_19[28], stage2_19[29]},
      {stage3_21[4],stage3_20[4],stage3_19[5],stage3_18[11],stage3_17[12]}
   );
   gpc615_5 gpc3463 (
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4]},
      {stage2_19[30]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[5],stage3_20[5],stage3_19[6],stage3_18[12]}
   );
   gpc615_5 gpc3464 (
      {stage2_18[5], stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9]},
      {stage2_19[31]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[6],stage3_20[6],stage3_19[7],stage3_18[13]}
   );
   gpc615_5 gpc3465 (
      {stage2_18[10], stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14]},
      {stage2_19[32]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[7],stage3_20[7],stage3_19[8],stage3_18[14]}
   );
   gpc615_5 gpc3466 (
      {stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18], stage2_18[19]},
      {stage2_19[33]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[8],stage3_20[8],stage3_19[9],stage3_18[15]}
   );
   gpc615_5 gpc3467 (
      {stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24]},
      {stage2_19[34]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[9],stage3_20[9],stage3_19[10],stage3_18[16]}
   );
   gpc615_5 gpc3468 (
      {stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29]},
      {stage2_19[35]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[10],stage3_20[10],stage3_19[11],stage3_18[17]}
   );
   gpc615_5 gpc3469 (
      {stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34]},
      {stage2_19[36]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[11],stage3_20[11],stage3_19[12],stage3_18[18]}
   );
   gpc615_5 gpc3470 (
      {stage2_18[35], stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39]},
      {stage2_19[37]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[7],stage3_21[12],stage3_20[12],stage3_19[13],stage3_18[19]}
   );
   gpc615_5 gpc3471 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4]},
      {stage2_22[0]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[8],stage3_21[13]}
   );
   gpc615_5 gpc3472 (
      {stage2_21[5], stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9]},
      {stage2_22[1]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[9],stage3_21[14]}
   );
   gpc615_5 gpc3473 (
      {stage2_21[10], stage2_21[11], stage2_21[12], stage2_21[13], stage2_21[14]},
      {stage2_22[2]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[10],stage3_21[15]}
   );
   gpc615_5 gpc3474 (
      {stage2_21[15], stage2_21[16], stage2_21[17], stage2_21[18], stage2_21[19]},
      {stage2_22[3]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[11],stage3_21[16]}
   );
   gpc615_5 gpc3475 (
      {stage2_21[20], stage2_21[21], stage2_21[22], stage2_21[23], stage2_21[24]},
      {stage2_22[4]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[4],stage3_24[4],stage3_23[4],stage3_22[12],stage3_21[17]}
   );
   gpc615_5 gpc3476 (
      {stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28], stage2_21[29]},
      {stage2_22[5]},
      {stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35]},
      {stage3_25[5],stage3_24[5],stage3_23[5],stage3_22[13],stage3_21[18]}
   );
   gpc615_5 gpc3477 (
      {stage2_21[30], stage2_21[31], stage2_21[32], stage2_21[33], stage2_21[34]},
      {stage2_22[6]},
      {stage2_23[36], stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40], stage2_23[41]},
      {stage3_25[6],stage3_24[6],stage3_23[6],stage3_22[14],stage3_21[19]}
   );
   gpc615_5 gpc3478 (
      {stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage2_23[42]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[7],stage3_24[7],stage3_23[7],stage3_22[15]}
   );
   gpc615_5 gpc3479 (
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16]},
      {stage2_23[43]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[8],stage3_24[8],stage3_23[8],stage3_22[16]}
   );
   gpc615_5 gpc3480 (
      {stage2_22[17], stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21]},
      {stage2_23[44]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[9],stage3_24[9],stage3_23[9],stage3_22[17]}
   );
   gpc615_5 gpc3481 (
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22]},
      {stage2_25[0]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[0],stage3_26[3],stage3_25[10],stage3_24[10]}
   );
   gpc615_5 gpc3482 (
      {stage2_24[23], stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27]},
      {stage2_25[1]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[1],stage3_26[4],stage3_25[11],stage3_24[11]}
   );
   gpc615_5 gpc3483 (
      {stage2_24[28], stage2_24[29], stage2_24[30], stage2_24[31], stage2_24[32]},
      {stage2_25[2]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[2],stage3_26[5],stage3_25[12],stage3_24[12]}
   );
   gpc606_5 gpc3484 (
      {stage2_25[3], stage2_25[4], stage2_25[5], stage2_25[6], stage2_25[7], stage2_25[8]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[3],stage3_27[3],stage3_26[6],stage3_25[13]}
   );
   gpc606_5 gpc3485 (
      {stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12], stage2_25[13], stage2_25[14]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[4],stage3_27[4],stage3_26[7],stage3_25[14]}
   );
   gpc606_5 gpc3486 (
      {stage2_25[15], stage2_25[16], stage2_25[17], stage2_25[18], stage2_25[19], stage2_25[20]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[5],stage3_27[5],stage3_26[8],stage3_25[15]}
   );
   gpc606_5 gpc3487 (
      {stage2_25[21], stage2_25[22], stage2_25[23], stage2_25[24], stage2_25[25], stage2_25[26]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[6],stage3_27[6],stage3_26[9],stage3_25[16]}
   );
   gpc606_5 gpc3488 (
      {stage2_25[27], stage2_25[28], stage2_25[29], stage2_25[30], stage2_25[31], stage2_25[32]},
      {stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29]},
      {stage3_29[4],stage3_28[7],stage3_27[7],stage3_26[10],stage3_25[17]}
   );
   gpc207_4 gpc3489 (
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23], stage2_26[24]},
      {stage2_28[0], stage2_28[1]},
      {stage3_29[5],stage3_28[8],stage3_27[8],stage3_26[11]}
   );
   gpc207_4 gpc3490 (
      {stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29], stage2_26[30], stage2_26[31]},
      {stage2_28[2], stage2_28[3]},
      {stage3_29[6],stage3_28[9],stage3_27[9],stage3_26[12]}
   );
   gpc207_4 gpc3491 (
      {stage2_26[32], stage2_26[33], stage2_26[34], stage2_26[35], stage2_26[36], stage2_26[37], stage2_26[38]},
      {stage2_28[4], stage2_28[5]},
      {stage3_29[7],stage3_28[10],stage3_27[10],stage3_26[13]}
   );
   gpc207_4 gpc3492 (
      {stage2_26[39], stage2_26[40], stage2_26[41], stage2_26[42], stage2_26[43], stage2_26[44], stage2_26[45]},
      {stage2_28[6], stage2_28[7]},
      {stage3_29[8],stage3_28[11],stage3_27[11],stage3_26[14]}
   );
   gpc207_4 gpc3493 (
      {stage2_26[46], stage2_26[47], stage2_26[48], stage2_26[49], stage2_26[50], stage2_26[51], stage2_26[52]},
      {stage2_28[8], stage2_28[9]},
      {stage3_29[9],stage3_28[12],stage3_27[12],stage3_26[15]}
   );
   gpc606_5 gpc3494 (
      {stage2_27[30], stage2_27[31], stage2_27[32], stage2_27[33], stage2_27[34], stage2_27[35]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[0],stage3_29[10],stage3_28[13],stage3_27[13]}
   );
   gpc606_5 gpc3495 (
      {stage2_27[36], stage2_27[37], stage2_27[38], stage2_27[39], stage2_27[40], stage2_27[41]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[1],stage3_29[11],stage3_28[14],stage3_27[14]}
   );
   gpc615_5 gpc3496 (
      {stage2_27[42], stage2_27[43], stage2_27[44], stage2_27[45], stage2_27[46]},
      {stage2_28[10]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[2],stage3_29[12],stage3_28[15],stage3_27[15]}
   );
   gpc606_5 gpc3497 (
      {stage2_28[11], stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[3],stage3_30[3],stage3_29[13],stage3_28[16]}
   );
   gpc606_5 gpc3498 (
      {stage2_28[17], stage2_28[18], stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[4],stage3_30[4],stage3_29[14],stage3_28[17]}
   );
   gpc606_5 gpc3499 (
      {stage2_28[23], stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[5],stage3_30[5],stage3_29[15],stage3_28[18]}
   );
   gpc606_5 gpc3500 (
      {stage2_28[29], stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[6],stage3_30[6],stage3_29[16],stage3_28[19]}
   );
   gpc606_5 gpc3501 (
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[4],stage3_31[7],stage3_30[7],stage3_29[17]}
   );
   gpc606_5 gpc3502 (
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[5],stage3_31[8],stage3_30[8],stage3_29[18]}
   );
   gpc606_5 gpc3503 (
      {stage2_29[30], stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[2],stage3_32[6],stage3_31[9],stage3_30[9],stage3_29[19]}
   );
   gpc606_5 gpc3504 (
      {stage2_29[36], stage2_29[37], stage2_29[38], stage2_29[39], stage2_29[40], stage2_29[41]},
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage3_33[3],stage3_32[7],stage3_31[10],stage3_30[10],stage3_29[20]}
   );
   gpc606_5 gpc3505 (
      {stage2_29[42], stage2_29[43], stage2_29[44], stage2_29[45], stage2_29[46], stage2_29[47]},
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage3_33[4],stage3_32[8],stage3_31[11],stage3_30[11],stage3_29[21]}
   );
   gpc615_5 gpc3506 (
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28]},
      {stage2_31[30]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[5],stage3_32[9],stage3_31[12],stage3_30[12]}
   );
   gpc615_5 gpc3507 (
      {stage2_30[29], stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33]},
      {stage2_31[31]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[6],stage3_32[10],stage3_31[13],stage3_30[13]}
   );
   gpc615_5 gpc3508 (
      {stage2_30[34], stage2_30[35], stage2_30[36], stage2_30[37], stage2_30[38]},
      {stage2_31[32]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[7],stage3_32[11],stage3_31[14],stage3_30[14]}
   );
   gpc606_5 gpc3509 (
      {stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[0],stage3_34[3],stage3_33[8],stage3_32[12]}
   );
   gpc606_5 gpc3510 (
      {stage2_32[24], stage2_32[25], stage2_32[26], stage2_32[27], stage2_32[28], stage2_32[29]},
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage3_36[1],stage3_35[1],stage3_34[4],stage3_33[9],stage3_32[13]}
   );
   gpc606_5 gpc3511 (
      {stage2_32[30], stage2_32[31], stage2_32[32], stage2_32[33], stage2_32[34], stage2_32[35]},
      {stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17]},
      {stage3_36[2],stage3_35[2],stage3_34[5],stage3_33[10],stage3_32[14]}
   );
   gpc7_3 gpc3512 (
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5], stage2_33[6]},
      {stage3_35[3],stage3_34[6],stage3_33[11]}
   );
   gpc7_3 gpc3513 (
      {stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11], stage2_33[12], stage2_33[13]},
      {stage3_35[4],stage3_34[7],stage3_33[12]}
   );
   gpc7_3 gpc3514 (
      {stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17], stage2_33[18], stage2_33[19], stage2_33[20]},
      {stage3_35[5],stage3_34[8],stage3_33[13]}
   );
   gpc7_3 gpc3515 (
      {stage2_33[21], stage2_33[22], stage2_33[23], stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27]},
      {stage3_35[6],stage3_34[9],stage3_33[14]}
   );
   gpc615_5 gpc3516 (
      {stage2_34[18], stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22]},
      {stage2_35[0]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[0],stage3_36[3],stage3_35[7],stage3_34[10]}
   );
   gpc606_5 gpc3517 (
      {stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5], stage2_35[6]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[1],stage3_37[1],stage3_36[4],stage3_35[8]}
   );
   gpc606_5 gpc3518 (
      {stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11], stage2_35[12]},
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage3_39[1],stage3_38[2],stage3_37[2],stage3_36[5],stage3_35[9]}
   );
   gpc615_5 gpc3519 (
      {stage2_35[13], stage2_35[14], stage2_35[15], stage2_35[16], stage2_35[17]},
      {stage2_36[6]},
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage3_39[2],stage3_38[3],stage3_37[3],stage3_36[6],stage3_35[10]}
   );
   gpc615_5 gpc3520 (
      {stage2_35[18], stage2_35[19], stage2_35[20], stage2_35[21], stage2_35[22]},
      {stage2_36[7]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage3_39[3],stage3_38[4],stage3_37[4],stage3_36[7],stage3_35[11]}
   );
   gpc615_5 gpc3521 (
      {stage2_35[23], stage2_35[24], stage2_35[25], stage2_35[26], stage2_35[27]},
      {stage2_36[8]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage3_39[4],stage3_38[5],stage3_37[5],stage3_36[8],stage3_35[12]}
   );
   gpc615_5 gpc3522 (
      {stage2_35[28], stage2_35[29], stage2_35[30], stage2_35[31], stage2_35[32]},
      {stage2_36[9]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage3_39[5],stage3_38[6],stage3_37[6],stage3_36[9],stage3_35[13]}
   );
   gpc606_5 gpc3523 (
      {stage2_36[10], stage2_36[11], stage2_36[12], stage2_36[13], stage2_36[14], stage2_36[15]},
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage3_40[0],stage3_39[6],stage3_38[7],stage3_37[7],stage3_36[10]}
   );
   gpc606_5 gpc3524 (
      {stage2_36[16], stage2_36[17], stage2_36[18], stage2_36[19], stage2_36[20], stage2_36[21]},
      {stage2_38[6], stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11]},
      {stage3_40[1],stage3_39[7],stage3_38[8],stage3_37[8],stage3_36[11]}
   );
   gpc606_5 gpc3525 (
      {stage2_36[22], stage2_36[23], stage2_36[24], stage2_36[25], stage2_36[26], stage2_36[27]},
      {stage2_38[12], stage2_38[13], stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17]},
      {stage3_40[2],stage3_39[8],stage3_38[9],stage3_37[9],stage3_36[12]}
   );
   gpc606_5 gpc3526 (
      {stage2_36[28], stage2_36[29], stage2_36[30], stage2_36[31], stage2_36[32], stage2_36[33]},
      {stage2_38[18], stage2_38[19], stage2_38[20], stage2_38[21], stage2_38[22], stage2_38[23]},
      {stage3_40[3],stage3_39[9],stage3_38[10],stage3_37[10],stage3_36[13]}
   );
   gpc606_5 gpc3527 (
      {stage2_37[36], stage2_37[37], stage2_37[38], stage2_37[39], stage2_37[40], stage2_37[41]},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5]},
      {stage3_41[0],stage3_40[4],stage3_39[10],stage3_38[11],stage3_37[11]}
   );
   gpc615_5 gpc3528 (
      {stage2_38[24], stage2_38[25], stage2_38[26], stage2_38[27], stage2_38[28]},
      {stage2_39[6]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[1],stage3_40[5],stage3_39[11],stage3_38[12]}
   );
   gpc615_5 gpc3529 (
      {stage2_38[29], stage2_38[30], stage2_38[31], stage2_38[32], 1'b0},
      {stage2_39[7]},
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage3_42[1],stage3_41[2],stage3_40[6],stage3_39[12],stage3_38[13]}
   );
   gpc606_5 gpc3530 (
      {stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11], stage2_39[12], stage2_39[13]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[2],stage3_41[3],stage3_40[7],stage3_39[13]}
   );
   gpc606_5 gpc3531 (
      {stage2_39[14], stage2_39[15], stage2_39[16], stage2_39[17], stage2_39[18], stage2_39[19]},
      {stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11]},
      {stage3_43[1],stage3_42[3],stage3_41[4],stage3_40[8],stage3_39[14]}
   );
   gpc606_5 gpc3532 (
      {stage2_39[20], stage2_39[21], stage2_39[22], stage2_39[23], stage2_39[24], stage2_39[25]},
      {stage2_41[12], stage2_41[13], stage2_41[14], stage2_41[15], stage2_41[16], stage2_41[17]},
      {stage3_43[2],stage3_42[4],stage3_41[5],stage3_40[9],stage3_39[15]}
   );
   gpc606_5 gpc3533 (
      {stage2_40[12], stage2_40[13], stage2_40[14], stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[3],stage3_42[5],stage3_41[6],stage3_40[10]}
   );
   gpc606_5 gpc3534 (
      {stage2_40[18], stage2_40[19], stage2_40[20], stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage3_44[1],stage3_43[4],stage3_42[6],stage3_41[7],stage3_40[11]}
   );
   gpc606_5 gpc3535 (
      {stage2_40[24], stage2_40[25], stage2_40[26], stage2_40[27], stage2_40[28], stage2_40[29]},
      {stage2_42[12], stage2_42[13], stage2_42[14], stage2_42[15], stage2_42[16], stage2_42[17]},
      {stage3_44[2],stage3_43[5],stage3_42[7],stage3_41[8],stage3_40[12]}
   );
   gpc606_5 gpc3536 (
      {stage2_41[18], stage2_41[19], stage2_41[20], stage2_41[21], stage2_41[22], stage2_41[23]},
      {stage2_43[0], stage2_43[1], stage2_43[2], stage2_43[3], stage2_43[4], stage2_43[5]},
      {stage3_45[0],stage3_44[3],stage3_43[6],stage3_42[8],stage3_41[9]}
   );
   gpc606_5 gpc3537 (
      {stage2_41[24], stage2_41[25], stage2_41[26], stage2_41[27], stage2_41[28], stage2_41[29]},
      {stage2_43[6], stage2_43[7], stage2_43[8], stage2_43[9], stage2_43[10], stage2_43[11]},
      {stage3_45[1],stage3_44[4],stage3_43[7],stage3_42[9],stage3_41[10]}
   );
   gpc615_5 gpc3538 (
      {stage2_41[30], stage2_41[31], stage2_41[32], stage2_41[33], stage2_41[34]},
      {stage2_42[18]},
      {stage2_43[12], stage2_43[13], stage2_43[14], stage2_43[15], stage2_43[16], stage2_43[17]},
      {stage3_45[2],stage3_44[5],stage3_43[8],stage3_42[10],stage3_41[11]}
   );
   gpc615_5 gpc3539 (
      {stage2_41[35], stage2_41[36], stage2_41[37], stage2_41[38], stage2_41[39]},
      {stage2_42[19]},
      {stage2_43[18], stage2_43[19], stage2_43[20], stage2_43[21], stage2_43[22], stage2_43[23]},
      {stage3_45[3],stage3_44[6],stage3_43[9],stage3_42[11],stage3_41[12]}
   );
   gpc615_5 gpc3540 (
      {stage2_41[40], stage2_41[41], stage2_41[42], stage2_41[43], stage2_41[44]},
      {stage2_42[20]},
      {stage2_43[24], stage2_43[25], stage2_43[26], stage2_43[27], stage2_43[28], stage2_43[29]},
      {stage3_45[4],stage3_44[7],stage3_43[10],stage3_42[12],stage3_41[13]}
   );
   gpc615_5 gpc3541 (
      {stage2_42[21], stage2_42[22], stage2_42[23], stage2_42[24], stage2_42[25]},
      {stage2_43[30]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[5],stage3_44[8],stage3_43[11],stage3_42[13]}
   );
   gpc615_5 gpc3542 (
      {stage2_42[26], stage2_42[27], stage2_42[28], stage2_42[29], stage2_42[30]},
      {stage2_43[31]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[6],stage3_44[9],stage3_43[12],stage3_42[14]}
   );
   gpc615_5 gpc3543 (
      {stage2_42[31], stage2_42[32], stage2_42[33], stage2_42[34], stage2_42[35]},
      {stage2_43[32]},
      {stage2_44[12], stage2_44[13], stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17]},
      {stage3_46[2],stage3_45[7],stage3_44[10],stage3_43[13],stage3_42[15]}
   );
   gpc615_5 gpc3544 (
      {stage2_42[36], stage2_42[37], stage2_42[38], stage2_42[39], stage2_42[40]},
      {stage2_43[33]},
      {stage2_44[18], stage2_44[19], stage2_44[20], stage2_44[21], stage2_44[22], stage2_44[23]},
      {stage3_46[3],stage3_45[8],stage3_44[11],stage3_43[14],stage3_42[16]}
   );
   gpc615_5 gpc3545 (
      {stage2_42[41], stage2_42[42], stage2_42[43], stage2_42[44], stage2_42[45]},
      {stage2_43[34]},
      {stage2_44[24], stage2_44[25], stage2_44[26], stage2_44[27], stage2_44[28], stage2_44[29]},
      {stage3_46[4],stage3_45[9],stage3_44[12],stage3_43[15],stage3_42[17]}
   );
   gpc615_5 gpc3546 (
      {stage2_42[46], stage2_42[47], stage2_42[48], stage2_42[49], stage2_42[50]},
      {stage2_43[35]},
      {stage2_44[30], stage2_44[31], stage2_44[32], stage2_44[33], stage2_44[34], stage2_44[35]},
      {stage3_46[5],stage3_45[10],stage3_44[13],stage3_43[16],stage3_42[18]}
   );
   gpc615_5 gpc3547 (
      {stage2_42[51], stage2_42[52], stage2_42[53], stage2_42[54], stage2_42[55]},
      {stage2_43[36]},
      {stage2_44[36], stage2_44[37], stage2_44[38], stage2_44[39], stage2_44[40], stage2_44[41]},
      {stage3_46[6],stage3_45[11],stage3_44[14],stage3_43[17],stage3_42[19]}
   );
   gpc615_5 gpc3548 (
      {stage2_43[37], stage2_43[38], stage2_43[39], stage2_43[40], stage2_43[41]},
      {stage2_44[42]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[7],stage3_45[12],stage3_44[15],stage3_43[18]}
   );
   gpc615_5 gpc3549 (
      {stage2_43[42], stage2_43[43], stage2_43[44], stage2_43[45], stage2_43[46]},
      {stage2_44[43]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[8],stage3_45[13],stage3_44[16],stage3_43[19]}
   );
   gpc615_5 gpc3550 (
      {stage2_43[47], stage2_43[48], stage2_43[49], stage2_43[50], stage2_43[51]},
      {stage2_44[44]},
      {stage2_45[12], stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage3_47[2],stage3_46[9],stage3_45[14],stage3_44[17],stage3_43[20]}
   );
   gpc615_5 gpc3551 (
      {stage2_44[45], stage2_44[46], stage2_44[47], stage2_44[48], stage2_44[49]},
      {stage2_45[18]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[3],stage3_46[10],stage3_45[15],stage3_44[18]}
   );
   gpc615_5 gpc3552 (
      {stage2_44[50], stage2_44[51], stage2_44[52], stage2_44[53], stage2_44[54]},
      {stage2_45[19]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[4],stage3_46[11],stage3_45[16],stage3_44[19]}
   );
   gpc606_5 gpc3553 (
      {stage2_45[20], stage2_45[21], stage2_45[22], stage2_45[23], stage2_45[24], stage2_45[25]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[2],stage3_47[5],stage3_46[12],stage3_45[17]}
   );
   gpc606_5 gpc3554 (
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage2_48[0], stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage3_50[0],stage3_49[1],stage3_48[3],stage3_47[6],stage3_46[13]}
   );
   gpc1325_5 gpc3555 (
      {stage2_46[18], stage2_46[19], stage2_46[20], stage2_46[21], stage2_46[22]},
      {stage2_47[6], stage2_47[7]},
      {stage2_48[6], stage2_48[7], stage2_48[8]},
      {stage2_49[0]},
      {stage3_50[1],stage3_49[2],stage3_48[4],stage3_47[7],stage3_46[14]}
   );
   gpc1325_5 gpc3556 (
      {stage2_46[23], stage2_46[24], stage2_46[25], stage2_46[26], stage2_46[27]},
      {stage2_47[8], stage2_47[9]},
      {stage2_48[9], stage2_48[10], stage2_48[11]},
      {stage2_49[1]},
      {stage3_50[2],stage3_49[3],stage3_48[5],stage3_47[8],stage3_46[15]}
   );
   gpc1325_5 gpc3557 (
      {stage2_46[28], stage2_46[29], stage2_46[30], stage2_46[31], stage2_46[32]},
      {stage2_47[10], stage2_47[11]},
      {stage2_48[12], stage2_48[13], stage2_48[14]},
      {stage2_49[2]},
      {stage3_50[3],stage3_49[4],stage3_48[6],stage3_47[9],stage3_46[16]}
   );
   gpc615_5 gpc3558 (
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16]},
      {stage2_48[15]},
      {stage2_49[3], stage2_49[4], stage2_49[5], stage2_49[6], stage2_49[7], stage2_49[8]},
      {stage3_51[0],stage3_50[4],stage3_49[5],stage3_48[7],stage3_47[10]}
   );
   gpc615_5 gpc3559 (
      {stage2_47[17], stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21]},
      {stage2_48[16]},
      {stage2_49[9], stage2_49[10], stage2_49[11], stage2_49[12], stage2_49[13], stage2_49[14]},
      {stage3_51[1],stage3_50[5],stage3_49[6],stage3_48[8],stage3_47[11]}
   );
   gpc615_5 gpc3560 (
      {stage2_47[22], stage2_47[23], stage2_47[24], stage2_47[25], stage2_47[26]},
      {stage2_48[17]},
      {stage2_49[15], stage2_49[16], stage2_49[17], stage2_49[18], stage2_49[19], stage2_49[20]},
      {stage3_51[2],stage3_50[6],stage3_49[7],stage3_48[9],stage3_47[12]}
   );
   gpc615_5 gpc3561 (
      {stage2_47[27], stage2_47[28], stage2_47[29], stage2_47[30], stage2_47[31]},
      {stage2_48[18]},
      {stage2_49[21], stage2_49[22], stage2_49[23], stage2_49[24], stage2_49[25], stage2_49[26]},
      {stage3_51[3],stage3_50[7],stage3_49[8],stage3_48[10],stage3_47[13]}
   );
   gpc615_5 gpc3562 (
      {stage2_47[32], stage2_47[33], stage2_47[34], stage2_47[35], stage2_47[36]},
      {stage2_48[19]},
      {stage2_49[27], stage2_49[28], stage2_49[29], stage2_49[30], stage2_49[31], stage2_49[32]},
      {stage3_51[4],stage3_50[8],stage3_49[9],stage3_48[11],stage3_47[14]}
   );
   gpc2116_5 gpc3563 (
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage2_51[0]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1]},
      {stage3_54[0],stage3_53[0],stage3_52[0],stage3_51[5],stage3_50[9]}
   );
   gpc2116_5 gpc3564 (
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage2_51[1]},
      {stage2_52[1]},
      {stage2_53[2], stage2_53[3]},
      {stage3_54[1],stage3_53[1],stage3_52[1],stage3_51[6],stage3_50[10]}
   );
   gpc615_5 gpc3565 (
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16]},
      {stage2_51[2]},
      {stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5], stage2_52[6], stage2_52[7]},
      {stage3_54[2],stage3_53[2],stage3_52[2],stage3_51[7],stage3_50[11]}
   );
   gpc615_5 gpc3566 (
      {stage2_50[17], stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21]},
      {stage2_51[3]},
      {stage2_52[8], stage2_52[9], stage2_52[10], stage2_52[11], stage2_52[12], stage2_52[13]},
      {stage3_54[3],stage3_53[3],stage3_52[3],stage3_51[8],stage3_50[12]}
   );
   gpc615_5 gpc3567 (
      {stage2_51[4], stage2_51[5], stage2_51[6], stage2_51[7], stage2_51[8]},
      {stage2_52[14]},
      {stage2_53[4], stage2_53[5], stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9]},
      {stage3_55[0],stage3_54[4],stage3_53[4],stage3_52[4],stage3_51[9]}
   );
   gpc615_5 gpc3568 (
      {stage2_51[9], stage2_51[10], stage2_51[11], stage2_51[12], stage2_51[13]},
      {stage2_52[15]},
      {stage2_53[10], stage2_53[11], stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15]},
      {stage3_55[1],stage3_54[5],stage3_53[5],stage3_52[5],stage3_51[10]}
   );
   gpc615_5 gpc3569 (
      {stage2_51[14], stage2_51[15], stage2_51[16], stage2_51[17], stage2_51[18]},
      {stage2_52[16]},
      {stage2_53[16], stage2_53[17], stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21]},
      {stage3_55[2],stage3_54[6],stage3_53[6],stage3_52[6],stage3_51[11]}
   );
   gpc615_5 gpc3570 (
      {stage2_51[19], stage2_51[20], stage2_51[21], stage2_51[22], stage2_51[23]},
      {stage2_52[17]},
      {stage2_53[22], stage2_53[23], stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27]},
      {stage3_55[3],stage3_54[7],stage3_53[7],stage3_52[7],stage3_51[12]}
   );
   gpc606_5 gpc3571 (
      {stage2_53[28], stage2_53[29], stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[0],stage3_55[4],stage3_54[8],stage3_53[8]}
   );
   gpc606_5 gpc3572 (
      {stage2_53[34], stage2_53[35], stage2_53[36], stage2_53[37], stage2_53[38], stage2_53[39]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[1],stage3_55[5],stage3_54[9],stage3_53[9]}
   );
   gpc606_5 gpc3573 (
      {stage2_53[40], stage2_53[41], stage2_53[42], stage2_53[43], stage2_53[44], stage2_53[45]},
      {stage2_55[12], stage2_55[13], stage2_55[14], stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage3_57[2],stage3_56[2],stage3_55[6],stage3_54[10],stage3_53[10]}
   );
   gpc606_5 gpc3574 (
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5]},
      {stage3_58[0],stage3_57[3],stage3_56[3],stage3_55[7],stage3_54[11]}
   );
   gpc606_5 gpc3575 (
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9], stage2_56[10], stage2_56[11]},
      {stage3_58[1],stage3_57[4],stage3_56[4],stage3_55[8],stage3_54[12]}
   );
   gpc606_5 gpc3576 (
      {stage2_54[12], stage2_54[13], stage2_54[14], stage2_54[15], stage2_54[16], stage2_54[17]},
      {stage2_56[12], stage2_56[13], stage2_56[14], stage2_56[15], stage2_56[16], stage2_56[17]},
      {stage3_58[2],stage3_57[5],stage3_56[5],stage3_55[9],stage3_54[13]}
   );
   gpc615_5 gpc3577 (
      {stage2_54[18], stage2_54[19], stage2_54[20], stage2_54[21], stage2_54[22]},
      {stage2_55[18]},
      {stage2_56[18], stage2_56[19], stage2_56[20], stage2_56[21], stage2_56[22], stage2_56[23]},
      {stage3_58[3],stage3_57[6],stage3_56[6],stage3_55[10],stage3_54[14]}
   );
   gpc615_5 gpc3578 (
      {stage2_54[23], stage2_54[24], stage2_54[25], stage2_54[26], stage2_54[27]},
      {stage2_55[19]},
      {stage2_56[24], stage2_56[25], stage2_56[26], stage2_56[27], stage2_56[28], stage2_56[29]},
      {stage3_58[4],stage3_57[7],stage3_56[7],stage3_55[11],stage3_54[15]}
   );
   gpc615_5 gpc3579 (
      {stage2_55[20], stage2_55[21], stage2_55[22], stage2_55[23], stage2_55[24]},
      {stage2_56[30]},
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5]},
      {stage3_59[0],stage3_58[5],stage3_57[8],stage3_56[8],stage3_55[12]}
   );
   gpc615_5 gpc3580 (
      {stage2_55[25], stage2_55[26], stage2_55[27], stage2_55[28], stage2_55[29]},
      {stage2_56[31]},
      {stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10], stage2_57[11]},
      {stage3_59[1],stage3_58[6],stage3_57[9],stage3_56[9],stage3_55[13]}
   );
   gpc615_5 gpc3581 (
      {stage2_55[30], stage2_55[31], stage2_55[32], stage2_55[33], stage2_55[34]},
      {stage2_56[32]},
      {stage2_57[12], stage2_57[13], stage2_57[14], stage2_57[15], stage2_57[16], stage2_57[17]},
      {stage3_59[2],stage3_58[7],stage3_57[10],stage3_56[10],stage3_55[14]}
   );
   gpc606_5 gpc3582 (
      {stage2_57[18], stage2_57[19], stage2_57[20], stage2_57[21], stage2_57[22], stage2_57[23]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[0],stage3_59[3],stage3_58[8],stage3_57[11]}
   );
   gpc606_5 gpc3583 (
      {stage2_57[24], stage2_57[25], stage2_57[26], stage2_57[27], stage2_57[28], stage2_57[29]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[1],stage3_59[4],stage3_58[9],stage3_57[12]}
   );
   gpc1163_5 gpc3584 (
      {stage2_58[0], stage2_58[1], stage2_58[2]},
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17]},
      {stage2_60[0]},
      {stage2_61[0]},
      {stage3_62[0],stage3_61[2],stage3_60[2],stage3_59[5],stage3_58[10]}
   );
   gpc615_5 gpc3585 (
      {stage2_58[3], stage2_58[4], stage2_58[5], stage2_58[6], stage2_58[7]},
      {stage2_59[18]},
      {stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5], stage2_60[6]},
      {stage3_62[1],stage3_61[3],stage3_60[3],stage3_59[6],stage3_58[11]}
   );
   gpc615_5 gpc3586 (
      {stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11], stage2_58[12]},
      {stage2_59[19]},
      {stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11], stage2_60[12]},
      {stage3_62[2],stage3_61[4],stage3_60[4],stage3_59[7],stage3_58[12]}
   );
   gpc135_4 gpc3587 (
      {stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23], stage2_59[24]},
      {stage2_60[13], stage2_60[14], stage2_60[15]},
      {stage2_61[1]},
      {stage3_62[3],stage3_61[5],stage3_60[5],stage3_59[8]}
   );
   gpc606_5 gpc3588 (
      {stage2_59[25], stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29], stage2_59[30]},
      {stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5], stage2_61[6], stage2_61[7]},
      {stage3_63[0],stage3_62[4],stage3_61[6],stage3_60[6],stage3_59[9]}
   );
   gpc606_5 gpc3589 (
      {stage2_59[31], stage2_59[32], stage2_59[33], stage2_59[34], stage2_59[35], stage2_59[36]},
      {stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11], stage2_61[12], stage2_61[13]},
      {stage3_63[1],stage3_62[5],stage3_61[7],stage3_60[7],stage3_59[10]}
   );
   gpc606_5 gpc3590 (
      {stage2_59[37], stage2_59[38], stage2_59[39], stage2_59[40], stage2_59[41], stage2_59[42]},
      {stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17], stage2_61[18], stage2_61[19]},
      {stage3_63[2],stage3_62[6],stage3_61[8],stage3_60[8],stage3_59[11]}
   );
   gpc606_5 gpc3591 (
      {stage2_59[43], stage2_59[44], stage2_59[45], stage2_59[46], stage2_59[47], stage2_59[48]},
      {stage2_61[20], stage2_61[21], stage2_61[22], stage2_61[23], stage2_61[24], stage2_61[25]},
      {stage3_63[3],stage3_62[7],stage3_61[9],stage3_60[9],stage3_59[12]}
   );
   gpc606_5 gpc3592 (
      {stage2_59[49], stage2_59[50], stage2_59[51], stage2_59[52], stage2_59[53], stage2_59[54]},
      {stage2_61[26], stage2_61[27], stage2_61[28], stage2_61[29], stage2_61[30], stage2_61[31]},
      {stage3_63[4],stage3_62[8],stage3_61[10],stage3_60[10],stage3_59[13]}
   );
   gpc615_5 gpc3593 (
      {stage2_59[55], stage2_59[56], stage2_59[57], stage2_59[58], stage2_59[59]},
      {stage2_60[16]},
      {stage2_61[32], stage2_61[33], stage2_61[34], stage2_61[35], stage2_61[36], stage2_61[37]},
      {stage3_63[5],stage3_62[9],stage3_61[11],stage3_60[11],stage3_59[14]}
   );
   gpc615_5 gpc3594 (
      {stage2_59[60], stage2_59[61], stage2_59[62], stage2_59[63], stage2_59[64]},
      {stage2_60[17]},
      {stage2_61[38], stage2_61[39], stage2_61[40], stage2_61[41], stage2_61[42], stage2_61[43]},
      {stage3_63[6],stage3_62[10],stage3_61[12],stage3_60[12],stage3_59[15]}
   );
   gpc615_5 gpc3595 (
      {stage2_59[65], stage2_59[66], stage2_59[67], stage2_59[68], stage2_59[69]},
      {stage2_60[18]},
      {stage2_61[44], stage2_61[45], stage2_61[46], stage2_61[47], stage2_61[48], stage2_61[49]},
      {stage3_63[7],stage3_62[11],stage3_61[13],stage3_60[13],stage3_59[16]}
   );
   gpc606_5 gpc3596 (
      {stage2_60[19], stage2_60[20], stage2_60[21], 1'b0, 1'b0, 1'b0},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[8],stage3_62[12],stage3_61[14],stage3_60[14]}
   );
   gpc1163_5 gpc3597 (
      {stage2_61[50], stage2_61[51], stage2_61[52]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage2_63[0]},
      {stage2_64[0]},
      {stage3_65[0],stage3_64[1],stage3_63[9],stage3_62[13],stage3_61[15]}
   );
   gpc606_5 gpc3598 (
      {stage2_61[53], stage2_61[54], stage2_61[55], stage2_61[56], stage2_61[57], stage2_61[58]},
      {stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5], stage2_63[6]},
      {stage3_65[1],stage3_64[2],stage3_63[10],stage3_62[14],stage3_61[16]}
   );
   gpc1163_5 gpc3599 (
      {stage2_62[12], stage2_62[13], stage2_62[14]},
      {stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11], stage2_63[12]},
      {stage2_64[1]},
      {stage2_65[0]},
      {stage3_66[0],stage3_65[2],stage3_64[3],stage3_63[11],stage3_62[15]}
   );
   gpc1163_5 gpc3600 (
      {stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage2_63[13], stage2_63[14], stage2_63[15], stage2_63[16], stage2_63[17], stage2_63[18]},
      {stage2_64[2]},
      {stage2_65[1]},
      {stage3_66[1],stage3_65[3],stage3_64[4],stage3_63[12],stage3_62[16]}
   );
   gpc1163_5 gpc3601 (
      {stage2_62[18], stage2_62[19], stage2_62[20]},
      {stage2_63[19], stage2_63[20], stage2_63[21], stage2_63[22], stage2_63[23], stage2_63[24]},
      {stage2_64[3]},
      {stage2_65[2]},
      {stage3_66[2],stage3_65[4],stage3_64[5],stage3_63[13],stage3_62[17]}
   );
   gpc1163_5 gpc3602 (
      {stage2_62[21], stage2_62[22], stage2_62[23]},
      {stage2_63[25], stage2_63[26], stage2_63[27], stage2_63[28], stage2_63[29], stage2_63[30]},
      {stage2_64[4]},
      {stage2_65[3]},
      {stage3_66[3],stage3_65[5],stage3_64[6],stage3_63[14],stage3_62[18]}
   );
   gpc606_5 gpc3603 (
      {stage2_62[24], stage2_62[25], stage2_62[26], stage2_62[27], stage2_62[28], stage2_62[29]},
      {stage2_64[5], stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9], stage2_64[10]},
      {stage3_66[4],stage3_65[6],stage3_64[7],stage3_63[15],stage3_62[19]}
   );
   gpc615_5 gpc3604 (
      {stage2_62[30], stage2_62[31], stage2_62[32], stage2_62[33], stage2_62[34]},
      {stage2_63[31]},
      {stage2_64[11], stage2_64[12], stage2_64[13], stage2_64[14], stage2_64[15], stage2_64[16]},
      {stage3_66[5],stage3_65[7],stage3_64[8],stage3_63[16],stage3_62[20]}
   );
   gpc606_5 gpc3605 (
      {stage2_63[32], stage2_63[33], stage2_63[34], stage2_63[35], stage2_63[36], stage2_63[37]},
      {stage2_65[4], stage2_65[5], stage2_65[6], stage2_65[7], stage2_65[8], stage2_65[9]},
      {stage3_67[0],stage3_66[6],stage3_65[8],stage3_64[9],stage3_63[17]}
   );
   gpc606_5 gpc3606 (
      {stage2_64[17], stage2_64[18], stage2_64[19], stage2_64[20], stage2_64[21], stage2_64[22]},
      {stage2_66[0], stage2_66[1], stage2_66[2], stage2_66[3], stage2_66[4], stage2_66[5]},
      {stage3_68[0],stage3_67[1],stage3_66[7],stage3_65[9],stage3_64[10]}
   );
   gpc606_5 gpc3607 (
      {stage2_64[23], stage2_64[24], stage2_64[25], stage2_64[26], stage2_64[27], stage2_64[28]},
      {stage2_66[6], stage2_66[7], stage2_66[8], stage2_66[9], 1'b0, 1'b0},
      {stage3_68[1],stage3_67[2],stage3_66[8],stage3_65[10],stage3_64[11]}
   );
   gpc1_1 gpc3608 (
      {stage2_0[3]},
      {stage3_0[1]}
   );
   gpc1_1 gpc3609 (
      {stage2_0[4]},
      {stage3_0[2]}
   );
   gpc1_1 gpc3610 (
      {stage2_0[5]},
      {stage3_0[3]}
   );
   gpc1_1 gpc3611 (
      {stage2_0[6]},
      {stage3_0[4]}
   );
   gpc1_1 gpc3612 (
      {stage2_0[7]},
      {stage3_0[5]}
   );
   gpc1_1 gpc3613 (
      {stage2_0[8]},
      {stage3_0[6]}
   );
   gpc1_1 gpc3614 (
      {stage2_0[9]},
      {stage3_0[7]}
   );
   gpc1_1 gpc3615 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc3616 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc3617 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc3618 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc3619 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc3620 (
      {stage2_1[11]},
      {stage3_1[6]}
   );
   gpc1_1 gpc3621 (
      {stage2_1[12]},
      {stage3_1[7]}
   );
   gpc1_1 gpc3622 (
      {stage2_1[13]},
      {stage3_1[8]}
   );
   gpc1_1 gpc3623 (
      {stage2_1[14]},
      {stage3_1[9]}
   );
   gpc1_1 gpc3624 (
      {stage2_1[15]},
      {stage3_1[10]}
   );
   gpc1_1 gpc3625 (
      {stage2_1[16]},
      {stage3_1[11]}
   );
   gpc1_1 gpc3626 (
      {stage2_1[17]},
      {stage3_1[12]}
   );
   gpc1_1 gpc3627 (
      {stage2_1[18]},
      {stage3_1[13]}
   );
   gpc1_1 gpc3628 (
      {stage2_2[34]},
      {stage3_2[7]}
   );
   gpc1_1 gpc3629 (
      {stage2_2[35]},
      {stage3_2[8]}
   );
   gpc1_1 gpc3630 (
      {stage2_2[36]},
      {stage3_2[9]}
   );
   gpc1_1 gpc3631 (
      {stage2_2[37]},
      {stage3_2[10]}
   );
   gpc1_1 gpc3632 (
      {stage2_3[19]},
      {stage3_3[10]}
   );
   gpc1_1 gpc3633 (
      {stage2_3[20]},
      {stage3_3[11]}
   );
   gpc1_1 gpc3634 (
      {stage2_3[21]},
      {stage3_3[12]}
   );
   gpc1_1 gpc3635 (
      {stage2_3[22]},
      {stage3_3[13]}
   );
   gpc1_1 gpc3636 (
      {stage2_4[45]},
      {stage3_4[11]}
   );
   gpc1_1 gpc3637 (
      {stage2_4[46]},
      {stage3_4[12]}
   );
   gpc1_1 gpc3638 (
      {stage2_4[47]},
      {stage3_4[13]}
   );
   gpc1_1 gpc3639 (
      {stage2_5[30]},
      {stage3_5[12]}
   );
   gpc1_1 gpc3640 (
      {stage2_5[31]},
      {stage3_5[13]}
   );
   gpc1_1 gpc3641 (
      {stage2_5[32]},
      {stage3_5[14]}
   );
   gpc1_1 gpc3642 (
      {stage2_5[33]},
      {stage3_5[15]}
   );
   gpc1_1 gpc3643 (
      {stage2_5[34]},
      {stage3_5[16]}
   );
   gpc1_1 gpc3644 (
      {stage2_5[35]},
      {stage3_5[17]}
   );
   gpc1_1 gpc3645 (
      {stage2_6[24]},
      {stage3_6[15]}
   );
   gpc1_1 gpc3646 (
      {stage2_6[25]},
      {stage3_6[16]}
   );
   gpc1_1 gpc3647 (
      {stage2_6[26]},
      {stage3_6[17]}
   );
   gpc1_1 gpc3648 (
      {stage2_6[27]},
      {stage3_6[18]}
   );
   gpc1_1 gpc3649 (
      {stage2_6[28]},
      {stage3_6[19]}
   );
   gpc1_1 gpc3650 (
      {stage2_7[37]},
      {stage3_7[13]}
   );
   gpc1_1 gpc3651 (
      {stage2_7[38]},
      {stage3_7[14]}
   );
   gpc1_1 gpc3652 (
      {stage2_7[39]},
      {stage3_7[15]}
   );
   gpc1_1 gpc3653 (
      {stage2_7[40]},
      {stage3_7[16]}
   );
   gpc1_1 gpc3654 (
      {stage2_9[22]},
      {stage3_9[17]}
   );
   gpc1_1 gpc3655 (
      {stage2_9[23]},
      {stage3_9[18]}
   );
   gpc1_1 gpc3656 (
      {stage2_9[24]},
      {stage3_9[19]}
   );
   gpc1_1 gpc3657 (
      {stage2_9[25]},
      {stage3_9[20]}
   );
   gpc1_1 gpc3658 (
      {stage2_11[36]},
      {stage3_11[15]}
   );
   gpc1_1 gpc3659 (
      {stage2_11[37]},
      {stage3_11[16]}
   );
   gpc1_1 gpc3660 (
      {stage2_11[38]},
      {stage3_11[17]}
   );
   gpc1_1 gpc3661 (
      {stage2_12[24]},
      {stage3_12[17]}
   );
   gpc1_1 gpc3662 (
      {stage2_12[25]},
      {stage3_12[18]}
   );
   gpc1_1 gpc3663 (
      {stage2_12[26]},
      {stage3_12[19]}
   );
   gpc1_1 gpc3664 (
      {stage2_12[27]},
      {stage3_12[20]}
   );
   gpc1_1 gpc3665 (
      {stage2_12[28]},
      {stage3_12[21]}
   );
   gpc1_1 gpc3666 (
      {stage2_12[29]},
      {stage3_12[22]}
   );
   gpc1_1 gpc3667 (
      {stage2_12[30]},
      {stage3_12[23]}
   );
   gpc1_1 gpc3668 (
      {stage2_13[36]},
      {stage3_13[11]}
   );
   gpc1_1 gpc3669 (
      {stage2_13[37]},
      {stage3_13[12]}
   );
   gpc1_1 gpc3670 (
      {stage2_13[38]},
      {stage3_13[13]}
   );
   gpc1_1 gpc3671 (
      {stage2_13[39]},
      {stage3_13[14]}
   );
   gpc1_1 gpc3672 (
      {stage2_13[40]},
      {stage3_13[15]}
   );
   gpc1_1 gpc3673 (
      {stage2_13[41]},
      {stage3_13[16]}
   );
   gpc1_1 gpc3674 (
      {stage2_13[42]},
      {stage3_13[17]}
   );
   gpc1_1 gpc3675 (
      {stage2_13[43]},
      {stage3_13[18]}
   );
   gpc1_1 gpc3676 (
      {stage2_13[44]},
      {stage3_13[19]}
   );
   gpc1_1 gpc3677 (
      {stage2_14[54]},
      {stage3_14[16]}
   );
   gpc1_1 gpc3678 (
      {stage2_14[55]},
      {stage3_14[17]}
   );
   gpc1_1 gpc3679 (
      {stage2_14[56]},
      {stage3_14[18]}
   );
   gpc1_1 gpc3680 (
      {stage2_14[57]},
      {stage3_14[19]}
   );
   gpc1_1 gpc3681 (
      {stage2_14[58]},
      {stage3_14[20]}
   );
   gpc1_1 gpc3682 (
      {stage2_14[59]},
      {stage3_14[21]}
   );
   gpc1_1 gpc3683 (
      {stage2_14[60]},
      {stage3_14[22]}
   );
   gpc1_1 gpc3684 (
      {stage2_14[61]},
      {stage3_14[23]}
   );
   gpc1_1 gpc3685 (
      {stage2_14[62]},
      {stage3_14[24]}
   );
   gpc1_1 gpc3686 (
      {stage2_14[63]},
      {stage3_14[25]}
   );
   gpc1_1 gpc3687 (
      {stage2_14[64]},
      {stage3_14[26]}
   );
   gpc1_1 gpc3688 (
      {stage2_14[65]},
      {stage3_14[27]}
   );
   gpc1_1 gpc3689 (
      {stage2_14[66]},
      {stage3_14[28]}
   );
   gpc1_1 gpc3690 (
      {stage2_14[67]},
      {stage3_14[29]}
   );
   gpc1_1 gpc3691 (
      {stage2_14[68]},
      {stage3_14[30]}
   );
   gpc1_1 gpc3692 (
      {stage2_14[69]},
      {stage3_14[31]}
   );
   gpc1_1 gpc3693 (
      {stage2_14[70]},
      {stage3_14[32]}
   );
   gpc1_1 gpc3694 (
      {stage2_14[71]},
      {stage3_14[33]}
   );
   gpc1_1 gpc3695 (
      {stage2_14[72]},
      {stage3_14[34]}
   );
   gpc1_1 gpc3696 (
      {stage2_14[73]},
      {stage3_14[35]}
   );
   gpc1_1 gpc3697 (
      {stage2_15[17]},
      {stage3_15[17]}
   );
   gpc1_1 gpc3698 (
      {stage2_15[18]},
      {stage3_15[18]}
   );
   gpc1_1 gpc3699 (
      {stage2_15[19]},
      {stage3_15[19]}
   );
   gpc1_1 gpc3700 (
      {stage2_15[20]},
      {stage3_15[20]}
   );
   gpc1_1 gpc3701 (
      {stage2_15[21]},
      {stage3_15[21]}
   );
   gpc1_1 gpc3702 (
      {stage2_15[22]},
      {stage3_15[22]}
   );
   gpc1_1 gpc3703 (
      {stage2_15[23]},
      {stage3_15[23]}
   );
   gpc1_1 gpc3704 (
      {stage2_15[24]},
      {stage3_15[24]}
   );
   gpc1_1 gpc3705 (
      {stage2_15[25]},
      {stage3_15[25]}
   );
   gpc1_1 gpc3706 (
      {stage2_15[26]},
      {stage3_15[26]}
   );
   gpc1_1 gpc3707 (
      {stage2_15[27]},
      {stage3_15[27]}
   );
   gpc1_1 gpc3708 (
      {stage2_15[28]},
      {stage3_15[28]}
   );
   gpc1_1 gpc3709 (
      {stage2_15[29]},
      {stage3_15[29]}
   );
   gpc1_1 gpc3710 (
      {stage2_15[30]},
      {stage3_15[30]}
   );
   gpc1_1 gpc3711 (
      {stage2_15[31]},
      {stage3_15[31]}
   );
   gpc1_1 gpc3712 (
      {stage2_15[32]},
      {stage3_15[32]}
   );
   gpc1_1 gpc3713 (
      {stage2_15[33]},
      {stage3_15[33]}
   );
   gpc1_1 gpc3714 (
      {stage2_15[34]},
      {stage3_15[34]}
   );
   gpc1_1 gpc3715 (
      {stage2_15[35]},
      {stage3_15[35]}
   );
   gpc1_1 gpc3716 (
      {stage2_15[36]},
      {stage3_15[36]}
   );
   gpc1_1 gpc3717 (
      {stage2_16[37]},
      {stage3_16[12]}
   );
   gpc1_1 gpc3718 (
      {stage2_16[38]},
      {stage3_16[13]}
   );
   gpc1_1 gpc3719 (
      {stage2_16[39]},
      {stage3_16[14]}
   );
   gpc1_1 gpc3720 (
      {stage2_16[40]},
      {stage3_16[15]}
   );
   gpc1_1 gpc3721 (
      {stage2_16[41]},
      {stage3_16[16]}
   );
   gpc1_1 gpc3722 (
      {stage2_16[42]},
      {stage3_16[17]}
   );
   gpc1_1 gpc3723 (
      {stage2_16[43]},
      {stage3_16[18]}
   );
   gpc1_1 gpc3724 (
      {stage2_16[44]},
      {stage3_16[19]}
   );
   gpc1_1 gpc3725 (
      {stage2_16[45]},
      {stage3_16[20]}
   );
   gpc1_1 gpc3726 (
      {stage2_16[46]},
      {stage3_16[21]}
   );
   gpc1_1 gpc3727 (
      {stage2_17[36]},
      {stage3_17[13]}
   );
   gpc1_1 gpc3728 (
      {stage2_17[37]},
      {stage3_17[14]}
   );
   gpc1_1 gpc3729 (
      {stage2_17[38]},
      {stage3_17[15]}
   );
   gpc1_1 gpc3730 (
      {stage2_17[39]},
      {stage3_17[16]}
   );
   gpc1_1 gpc3731 (
      {stage2_18[40]},
      {stage3_18[20]}
   );
   gpc1_1 gpc3732 (
      {stage2_18[41]},
      {stage3_18[21]}
   );
   gpc1_1 gpc3733 (
      {stage2_18[42]},
      {stage3_18[22]}
   );
   gpc1_1 gpc3734 (
      {stage2_19[38]},
      {stage3_19[14]}
   );
   gpc1_1 gpc3735 (
      {stage2_19[39]},
      {stage3_19[15]}
   );
   gpc1_1 gpc3736 (
      {stage2_19[40]},
      {stage3_19[16]}
   );
   gpc1_1 gpc3737 (
      {stage2_19[41]},
      {stage3_19[17]}
   );
   gpc1_1 gpc3738 (
      {stage2_19[42]},
      {stage3_19[18]}
   );
   gpc1_1 gpc3739 (
      {stage2_19[43]},
      {stage3_19[19]}
   );
   gpc1_1 gpc3740 (
      {stage2_19[44]},
      {stage3_19[20]}
   );
   gpc1_1 gpc3741 (
      {stage2_19[45]},
      {stage3_19[21]}
   );
   gpc1_1 gpc3742 (
      {stage2_19[46]},
      {stage3_19[22]}
   );
   gpc1_1 gpc3743 (
      {stage2_19[47]},
      {stage3_19[23]}
   );
   gpc1_1 gpc3744 (
      {stage2_19[48]},
      {stage3_19[24]}
   );
   gpc1_1 gpc3745 (
      {stage2_19[49]},
      {stage3_19[25]}
   );
   gpc1_1 gpc3746 (
      {stage2_19[50]},
      {stage3_19[26]}
   );
   gpc1_1 gpc3747 (
      {stage2_20[48]},
      {stage3_20[13]}
   );
   gpc1_1 gpc3748 (
      {stage2_20[49]},
      {stage3_20[14]}
   );
   gpc1_1 gpc3749 (
      {stage2_20[50]},
      {stage3_20[15]}
   );
   gpc1_1 gpc3750 (
      {stage2_20[51]},
      {stage3_20[16]}
   );
   gpc1_1 gpc3751 (
      {stage2_20[52]},
      {stage3_20[17]}
   );
   gpc1_1 gpc3752 (
      {stage2_20[53]},
      {stage3_20[18]}
   );
   gpc1_1 gpc3753 (
      {stage2_20[54]},
      {stage3_20[19]}
   );
   gpc1_1 gpc3754 (
      {stage2_20[55]},
      {stage3_20[20]}
   );
   gpc1_1 gpc3755 (
      {stage2_20[56]},
      {stage3_20[21]}
   );
   gpc1_1 gpc3756 (
      {stage2_20[57]},
      {stage3_20[22]}
   );
   gpc1_1 gpc3757 (
      {stage2_21[35]},
      {stage3_21[20]}
   );
   gpc1_1 gpc3758 (
      {stage2_21[36]},
      {stage3_21[21]}
   );
   gpc1_1 gpc3759 (
      {stage2_21[37]},
      {stage3_21[22]}
   );
   gpc1_1 gpc3760 (
      {stage2_21[38]},
      {stage3_21[23]}
   );
   gpc1_1 gpc3761 (
      {stage2_21[39]},
      {stage3_21[24]}
   );
   gpc1_1 gpc3762 (
      {stage2_22[22]},
      {stage3_22[18]}
   );
   gpc1_1 gpc3763 (
      {stage2_22[23]},
      {stage3_22[19]}
   );
   gpc1_1 gpc3764 (
      {stage2_22[24]},
      {stage3_22[20]}
   );
   gpc1_1 gpc3765 (
      {stage2_22[25]},
      {stage3_22[21]}
   );
   gpc1_1 gpc3766 (
      {stage2_22[26]},
      {stage3_22[22]}
   );
   gpc1_1 gpc3767 (
      {stage2_22[27]},
      {stage3_22[23]}
   );
   gpc1_1 gpc3768 (
      {stage2_22[28]},
      {stage3_22[24]}
   );
   gpc1_1 gpc3769 (
      {stage2_22[29]},
      {stage3_22[25]}
   );
   gpc1_1 gpc3770 (
      {stage2_22[30]},
      {stage3_22[26]}
   );
   gpc1_1 gpc3771 (
      {stage2_23[45]},
      {stage3_23[10]}
   );
   gpc1_1 gpc3772 (
      {stage2_23[46]},
      {stage3_23[11]}
   );
   gpc1_1 gpc3773 (
      {stage2_24[33]},
      {stage3_24[13]}
   );
   gpc1_1 gpc3774 (
      {stage2_24[34]},
      {stage3_24[14]}
   );
   gpc1_1 gpc3775 (
      {stage2_24[35]},
      {stage3_24[15]}
   );
   gpc1_1 gpc3776 (
      {stage2_24[36]},
      {stage3_24[16]}
   );
   gpc1_1 gpc3777 (
      {stage2_24[37]},
      {stage3_24[17]}
   );
   gpc1_1 gpc3778 (
      {stage2_24[38]},
      {stage3_24[18]}
   );
   gpc1_1 gpc3779 (
      {stage2_24[39]},
      {stage3_24[19]}
   );
   gpc1_1 gpc3780 (
      {stage2_24[40]},
      {stage3_24[20]}
   );
   gpc1_1 gpc3781 (
      {stage2_24[41]},
      {stage3_24[21]}
   );
   gpc1_1 gpc3782 (
      {stage2_24[42]},
      {stage3_24[22]}
   );
   gpc1_1 gpc3783 (
      {stage2_24[43]},
      {stage3_24[23]}
   );
   gpc1_1 gpc3784 (
      {stage2_24[44]},
      {stage3_24[24]}
   );
   gpc1_1 gpc3785 (
      {stage2_24[45]},
      {stage3_24[25]}
   );
   gpc1_1 gpc3786 (
      {stage2_25[33]},
      {stage3_25[18]}
   );
   gpc1_1 gpc3787 (
      {stage2_25[34]},
      {stage3_25[19]}
   );
   gpc1_1 gpc3788 (
      {stage2_25[35]},
      {stage3_25[20]}
   );
   gpc1_1 gpc3789 (
      {stage2_25[36]},
      {stage3_25[21]}
   );
   gpc1_1 gpc3790 (
      {stage2_27[47]},
      {stage3_27[16]}
   );
   gpc1_1 gpc3791 (
      {stage2_27[48]},
      {stage3_27[17]}
   );
   gpc1_1 gpc3792 (
      {stage2_27[49]},
      {stage3_27[18]}
   );
   gpc1_1 gpc3793 (
      {stage2_29[48]},
      {stage3_29[22]}
   );
   gpc1_1 gpc3794 (
      {stage2_29[49]},
      {stage3_29[23]}
   );
   gpc1_1 gpc3795 (
      {stage2_30[39]},
      {stage3_30[15]}
   );
   gpc1_1 gpc3796 (
      {stage2_30[40]},
      {stage3_30[16]}
   );
   gpc1_1 gpc3797 (
      {stage2_30[41]},
      {stage3_30[17]}
   );
   gpc1_1 gpc3798 (
      {stage2_30[42]},
      {stage3_30[18]}
   );
   gpc1_1 gpc3799 (
      {stage2_30[43]},
      {stage3_30[19]}
   );
   gpc1_1 gpc3800 (
      {stage2_30[44]},
      {stage3_30[20]}
   );
   gpc1_1 gpc3801 (
      {stage2_30[45]},
      {stage3_30[21]}
   );
   gpc1_1 gpc3802 (
      {stage2_30[46]},
      {stage3_30[22]}
   );
   gpc1_1 gpc3803 (
      {stage2_30[47]},
      {stage3_30[23]}
   );
   gpc1_1 gpc3804 (
      {stage2_30[48]},
      {stage3_30[24]}
   );
   gpc1_1 gpc3805 (
      {stage2_30[49]},
      {stage3_30[25]}
   );
   gpc1_1 gpc3806 (
      {stage2_31[33]},
      {stage3_31[15]}
   );
   gpc1_1 gpc3807 (
      {stage2_31[34]},
      {stage3_31[16]}
   );
   gpc1_1 gpc3808 (
      {stage2_31[35]},
      {stage3_31[17]}
   );
   gpc1_1 gpc3809 (
      {stage2_31[36]},
      {stage3_31[18]}
   );
   gpc1_1 gpc3810 (
      {stage2_31[37]},
      {stage3_31[19]}
   );
   gpc1_1 gpc3811 (
      {stage2_31[38]},
      {stage3_31[20]}
   );
   gpc1_1 gpc3812 (
      {stage2_32[36]},
      {stage3_32[15]}
   );
   gpc1_1 gpc3813 (
      {stage2_32[37]},
      {stage3_32[16]}
   );
   gpc1_1 gpc3814 (
      {stage2_32[38]},
      {stage3_32[17]}
   );
   gpc1_1 gpc3815 (
      {stage2_32[39]},
      {stage3_32[18]}
   );
   gpc1_1 gpc3816 (
      {stage2_32[40]},
      {stage3_32[19]}
   );
   gpc1_1 gpc3817 (
      {stage2_32[41]},
      {stage3_32[20]}
   );
   gpc1_1 gpc3818 (
      {stage2_32[42]},
      {stage3_32[21]}
   );
   gpc1_1 gpc3819 (
      {stage2_32[43]},
      {stage3_32[22]}
   );
   gpc1_1 gpc3820 (
      {stage2_32[44]},
      {stage3_32[23]}
   );
   gpc1_1 gpc3821 (
      {stage2_32[45]},
      {stage3_32[24]}
   );
   gpc1_1 gpc3822 (
      {stage2_32[46]},
      {stage3_32[25]}
   );
   gpc1_1 gpc3823 (
      {stage2_32[47]},
      {stage3_32[26]}
   );
   gpc1_1 gpc3824 (
      {stage2_32[48]},
      {stage3_32[27]}
   );
   gpc1_1 gpc3825 (
      {stage2_32[49]},
      {stage3_32[28]}
   );
   gpc1_1 gpc3826 (
      {stage2_32[50]},
      {stage3_32[29]}
   );
   gpc1_1 gpc3827 (
      {stage2_32[51]},
      {stage3_32[30]}
   );
   gpc1_1 gpc3828 (
      {stage2_32[52]},
      {stage3_32[31]}
   );
   gpc1_1 gpc3829 (
      {stage2_32[53]},
      {stage3_32[32]}
   );
   gpc1_1 gpc3830 (
      {stage2_32[54]},
      {stage3_32[33]}
   );
   gpc1_1 gpc3831 (
      {stage2_32[55]},
      {stage3_32[34]}
   );
   gpc1_1 gpc3832 (
      {stage2_34[23]},
      {stage3_34[11]}
   );
   gpc1_1 gpc3833 (
      {stage2_34[24]},
      {stage3_34[12]}
   );
   gpc1_1 gpc3834 (
      {stage2_34[25]},
      {stage3_34[13]}
   );
   gpc1_1 gpc3835 (
      {stage2_34[26]},
      {stage3_34[14]}
   );
   gpc1_1 gpc3836 (
      {stage2_34[27]},
      {stage3_34[15]}
   );
   gpc1_1 gpc3837 (
      {stage2_34[28]},
      {stage3_34[16]}
   );
   gpc1_1 gpc3838 (
      {stage2_34[29]},
      {stage3_34[17]}
   );
   gpc1_1 gpc3839 (
      {stage2_34[30]},
      {stage3_34[18]}
   );
   gpc1_1 gpc3840 (
      {stage2_34[31]},
      {stage3_34[19]}
   );
   gpc1_1 gpc3841 (
      {stage2_34[32]},
      {stage3_34[20]}
   );
   gpc1_1 gpc3842 (
      {stage2_34[33]},
      {stage3_34[21]}
   );
   gpc1_1 gpc3843 (
      {stage2_34[34]},
      {stage3_34[22]}
   );
   gpc1_1 gpc3844 (
      {stage2_35[33]},
      {stage3_35[14]}
   );
   gpc1_1 gpc3845 (
      {stage2_35[34]},
      {stage3_35[15]}
   );
   gpc1_1 gpc3846 (
      {stage2_35[35]},
      {stage3_35[16]}
   );
   gpc1_1 gpc3847 (
      {stage2_35[36]},
      {stage3_35[17]}
   );
   gpc1_1 gpc3848 (
      {stage2_35[37]},
      {stage3_35[18]}
   );
   gpc1_1 gpc3849 (
      {stage2_35[38]},
      {stage3_35[19]}
   );
   gpc1_1 gpc3850 (
      {stage2_35[39]},
      {stage3_35[20]}
   );
   gpc1_1 gpc3851 (
      {stage2_35[40]},
      {stage3_35[21]}
   );
   gpc1_1 gpc3852 (
      {stage2_35[41]},
      {stage3_35[22]}
   );
   gpc1_1 gpc3853 (
      {stage2_35[42]},
      {stage3_35[23]}
   );
   gpc1_1 gpc3854 (
      {stage2_35[43]},
      {stage3_35[24]}
   );
   gpc1_1 gpc3855 (
      {stage2_35[44]},
      {stage3_35[25]}
   );
   gpc1_1 gpc3856 (
      {stage2_36[34]},
      {stage3_36[14]}
   );
   gpc1_1 gpc3857 (
      {stage2_36[35]},
      {stage3_36[15]}
   );
   gpc1_1 gpc3858 (
      {stage2_36[36]},
      {stage3_36[16]}
   );
   gpc1_1 gpc3859 (
      {stage2_39[26]},
      {stage3_39[16]}
   );
   gpc1_1 gpc3860 (
      {stage2_39[27]},
      {stage3_39[17]}
   );
   gpc1_1 gpc3861 (
      {stage2_39[28]},
      {stage3_39[18]}
   );
   gpc1_1 gpc3862 (
      {stage2_39[29]},
      {stage3_39[19]}
   );
   gpc1_1 gpc3863 (
      {stage2_39[30]},
      {stage3_39[20]}
   );
   gpc1_1 gpc3864 (
      {stage2_39[31]},
      {stage3_39[21]}
   );
   gpc1_1 gpc3865 (
      {stage2_39[32]},
      {stage3_39[22]}
   );
   gpc1_1 gpc3866 (
      {stage2_39[33]},
      {stage3_39[23]}
   );
   gpc1_1 gpc3867 (
      {stage2_40[30]},
      {stage3_40[13]}
   );
   gpc1_1 gpc3868 (
      {stage2_40[31]},
      {stage3_40[14]}
   );
   gpc1_1 gpc3869 (
      {stage2_40[32]},
      {stage3_40[15]}
   );
   gpc1_1 gpc3870 (
      {stage2_40[33]},
      {stage3_40[16]}
   );
   gpc1_1 gpc3871 (
      {stage2_40[34]},
      {stage3_40[17]}
   );
   gpc1_1 gpc3872 (
      {stage2_40[35]},
      {stage3_40[18]}
   );
   gpc1_1 gpc3873 (
      {stage2_40[36]},
      {stage3_40[19]}
   );
   gpc1_1 gpc3874 (
      {stage2_40[37]},
      {stage3_40[20]}
   );
   gpc1_1 gpc3875 (
      {stage2_40[38]},
      {stage3_40[21]}
   );
   gpc1_1 gpc3876 (
      {stage2_40[39]},
      {stage3_40[22]}
   );
   gpc1_1 gpc3877 (
      {stage2_40[40]},
      {stage3_40[23]}
   );
   gpc1_1 gpc3878 (
      {stage2_41[45]},
      {stage3_41[14]}
   );
   gpc1_1 gpc3879 (
      {stage2_41[46]},
      {stage3_41[15]}
   );
   gpc1_1 gpc3880 (
      {stage2_41[47]},
      {stage3_41[16]}
   );
   gpc1_1 gpc3881 (
      {stage2_41[48]},
      {stage3_41[17]}
   );
   gpc1_1 gpc3882 (
      {stage2_41[49]},
      {stage3_41[18]}
   );
   gpc1_1 gpc3883 (
      {stage2_41[50]},
      {stage3_41[19]}
   );
   gpc1_1 gpc3884 (
      {stage2_41[51]},
      {stage3_41[20]}
   );
   gpc1_1 gpc3885 (
      {stage2_41[52]},
      {stage3_41[21]}
   );
   gpc1_1 gpc3886 (
      {stage2_41[53]},
      {stage3_41[22]}
   );
   gpc1_1 gpc3887 (
      {stage2_41[54]},
      {stage3_41[23]}
   );
   gpc1_1 gpc3888 (
      {stage2_41[55]},
      {stage3_41[24]}
   );
   gpc1_1 gpc3889 (
      {stage2_42[56]},
      {stage3_42[20]}
   );
   gpc1_1 gpc3890 (
      {stage2_42[57]},
      {stage3_42[21]}
   );
   gpc1_1 gpc3891 (
      {stage2_42[58]},
      {stage3_42[22]}
   );
   gpc1_1 gpc3892 (
      {stage2_42[59]},
      {stage3_42[23]}
   );
   gpc1_1 gpc3893 (
      {stage2_42[60]},
      {stage3_42[24]}
   );
   gpc1_1 gpc3894 (
      {stage2_42[61]},
      {stage3_42[25]}
   );
   gpc1_1 gpc3895 (
      {stage2_44[55]},
      {stage3_44[20]}
   );
   gpc1_1 gpc3896 (
      {stage2_44[56]},
      {stage3_44[21]}
   );
   gpc1_1 gpc3897 (
      {stage2_44[57]},
      {stage3_44[22]}
   );
   gpc1_1 gpc3898 (
      {stage2_44[58]},
      {stage3_44[23]}
   );
   gpc1_1 gpc3899 (
      {stage2_44[59]},
      {stage3_44[24]}
   );
   gpc1_1 gpc3900 (
      {stage2_44[60]},
      {stage3_44[25]}
   );
   gpc1_1 gpc3901 (
      {stage2_44[61]},
      {stage3_44[26]}
   );
   gpc1_1 gpc3902 (
      {stage2_44[62]},
      {stage3_44[27]}
   );
   gpc1_1 gpc3903 (
      {stage2_44[63]},
      {stage3_44[28]}
   );
   gpc1_1 gpc3904 (
      {stage2_44[64]},
      {stage3_44[29]}
   );
   gpc1_1 gpc3905 (
      {stage2_44[65]},
      {stage3_44[30]}
   );
   gpc1_1 gpc3906 (
      {stage2_47[37]},
      {stage3_47[15]}
   );
   gpc1_1 gpc3907 (
      {stage2_47[38]},
      {stage3_47[16]}
   );
   gpc1_1 gpc3908 (
      {stage2_47[39]},
      {stage3_47[17]}
   );
   gpc1_1 gpc3909 (
      {stage2_47[40]},
      {stage3_47[18]}
   );
   gpc1_1 gpc3910 (
      {stage2_47[41]},
      {stage3_47[19]}
   );
   gpc1_1 gpc3911 (
      {stage2_47[42]},
      {stage3_47[20]}
   );
   gpc1_1 gpc3912 (
      {stage2_47[43]},
      {stage3_47[21]}
   );
   gpc1_1 gpc3913 (
      {stage2_47[44]},
      {stage3_47[22]}
   );
   gpc1_1 gpc3914 (
      {stage2_47[45]},
      {stage3_47[23]}
   );
   gpc1_1 gpc3915 (
      {stage2_48[20]},
      {stage3_48[12]}
   );
   gpc1_1 gpc3916 (
      {stage2_48[21]},
      {stage3_48[13]}
   );
   gpc1_1 gpc3917 (
      {stage2_48[22]},
      {stage3_48[14]}
   );
   gpc1_1 gpc3918 (
      {stage2_48[23]},
      {stage3_48[15]}
   );
   gpc1_1 gpc3919 (
      {stage2_49[33]},
      {stage3_49[10]}
   );
   gpc1_1 gpc3920 (
      {stage2_49[34]},
      {stage3_49[11]}
   );
   gpc1_1 gpc3921 (
      {stage2_49[35]},
      {stage3_49[12]}
   );
   gpc1_1 gpc3922 (
      {stage2_49[36]},
      {stage3_49[13]}
   );
   gpc1_1 gpc3923 (
      {stage2_50[22]},
      {stage3_50[13]}
   );
   gpc1_1 gpc3924 (
      {stage2_50[23]},
      {stage3_50[14]}
   );
   gpc1_1 gpc3925 (
      {stage2_50[24]},
      {stage3_50[15]}
   );
   gpc1_1 gpc3926 (
      {stage2_50[25]},
      {stage3_50[16]}
   );
   gpc1_1 gpc3927 (
      {stage2_50[26]},
      {stage3_50[17]}
   );
   gpc1_1 gpc3928 (
      {stage2_50[27]},
      {stage3_50[18]}
   );
   gpc1_1 gpc3929 (
      {stage2_50[28]},
      {stage3_50[19]}
   );
   gpc1_1 gpc3930 (
      {stage2_50[29]},
      {stage3_50[20]}
   );
   gpc1_1 gpc3931 (
      {stage2_50[30]},
      {stage3_50[21]}
   );
   gpc1_1 gpc3932 (
      {stage2_50[31]},
      {stage3_50[22]}
   );
   gpc1_1 gpc3933 (
      {stage2_50[32]},
      {stage3_50[23]}
   );
   gpc1_1 gpc3934 (
      {stage2_50[33]},
      {stage3_50[24]}
   );
   gpc1_1 gpc3935 (
      {stage2_50[34]},
      {stage3_50[25]}
   );
   gpc1_1 gpc3936 (
      {stage2_50[35]},
      {stage3_50[26]}
   );
   gpc1_1 gpc3937 (
      {stage2_50[36]},
      {stage3_50[27]}
   );
   gpc1_1 gpc3938 (
      {stage2_50[37]},
      {stage3_50[28]}
   );
   gpc1_1 gpc3939 (
      {stage2_50[38]},
      {stage3_50[29]}
   );
   gpc1_1 gpc3940 (
      {stage2_50[39]},
      {stage3_50[30]}
   );
   gpc1_1 gpc3941 (
      {stage2_50[40]},
      {stage3_50[31]}
   );
   gpc1_1 gpc3942 (
      {stage2_51[24]},
      {stage3_51[13]}
   );
   gpc1_1 gpc3943 (
      {stage2_52[18]},
      {stage3_52[8]}
   );
   gpc1_1 gpc3944 (
      {stage2_52[19]},
      {stage3_52[9]}
   );
   gpc1_1 gpc3945 (
      {stage2_52[20]},
      {stage3_52[10]}
   );
   gpc1_1 gpc3946 (
      {stage2_52[21]},
      {stage3_52[11]}
   );
   gpc1_1 gpc3947 (
      {stage2_52[22]},
      {stage3_52[12]}
   );
   gpc1_1 gpc3948 (
      {stage2_52[23]},
      {stage3_52[13]}
   );
   gpc1_1 gpc3949 (
      {stage2_52[24]},
      {stage3_52[14]}
   );
   gpc1_1 gpc3950 (
      {stage2_52[25]},
      {stage3_52[15]}
   );
   gpc1_1 gpc3951 (
      {stage2_52[26]},
      {stage3_52[16]}
   );
   gpc1_1 gpc3952 (
      {stage2_52[27]},
      {stage3_52[17]}
   );
   gpc1_1 gpc3953 (
      {stage2_52[28]},
      {stage3_52[18]}
   );
   gpc1_1 gpc3954 (
      {stage2_52[29]},
      {stage3_52[19]}
   );
   gpc1_1 gpc3955 (
      {stage2_52[30]},
      {stage3_52[20]}
   );
   gpc1_1 gpc3956 (
      {stage2_52[31]},
      {stage3_52[21]}
   );
   gpc1_1 gpc3957 (
      {stage2_52[32]},
      {stage3_52[22]}
   );
   gpc1_1 gpc3958 (
      {stage2_52[33]},
      {stage3_52[23]}
   );
   gpc1_1 gpc3959 (
      {stage2_53[46]},
      {stage3_53[11]}
   );
   gpc1_1 gpc3960 (
      {stage2_53[47]},
      {stage3_53[12]}
   );
   gpc1_1 gpc3961 (
      {stage2_53[48]},
      {stage3_53[13]}
   );
   gpc1_1 gpc3962 (
      {stage2_53[49]},
      {stage3_53[14]}
   );
   gpc1_1 gpc3963 (
      {stage2_53[50]},
      {stage3_53[15]}
   );
   gpc1_1 gpc3964 (
      {stage2_55[35]},
      {stage3_55[15]}
   );
   gpc1_1 gpc3965 (
      {stage2_55[36]},
      {stage3_55[16]}
   );
   gpc1_1 gpc3966 (
      {stage2_55[37]},
      {stage3_55[17]}
   );
   gpc1_1 gpc3967 (
      {stage2_56[33]},
      {stage3_56[11]}
   );
   gpc1_1 gpc3968 (
      {stage2_56[34]},
      {stage3_56[12]}
   );
   gpc1_1 gpc3969 (
      {stage2_56[35]},
      {stage3_56[13]}
   );
   gpc1_1 gpc3970 (
      {stage2_56[36]},
      {stage3_56[14]}
   );
   gpc1_1 gpc3971 (
      {stage2_56[37]},
      {stage3_56[15]}
   );
   gpc1_1 gpc3972 (
      {stage2_56[38]},
      {stage3_56[16]}
   );
   gpc1_1 gpc3973 (
      {stage2_56[39]},
      {stage3_56[17]}
   );
   gpc1_1 gpc3974 (
      {stage2_56[40]},
      {stage3_56[18]}
   );
   gpc1_1 gpc3975 (
      {stage2_56[41]},
      {stage3_56[19]}
   );
   gpc1_1 gpc3976 (
      {stage2_56[42]},
      {stage3_56[20]}
   );
   gpc1_1 gpc3977 (
      {stage2_56[43]},
      {stage3_56[21]}
   );
   gpc1_1 gpc3978 (
      {stage2_56[44]},
      {stage3_56[22]}
   );
   gpc1_1 gpc3979 (
      {stage2_56[45]},
      {stage3_56[23]}
   );
   gpc1_1 gpc3980 (
      {stage2_56[46]},
      {stage3_56[24]}
   );
   gpc1_1 gpc3981 (
      {stage2_56[47]},
      {stage3_56[25]}
   );
   gpc1_1 gpc3982 (
      {stage2_56[48]},
      {stage3_56[26]}
   );
   gpc1_1 gpc3983 (
      {stage2_56[49]},
      {stage3_56[27]}
   );
   gpc1_1 gpc3984 (
      {stage2_56[50]},
      {stage3_56[28]}
   );
   gpc1_1 gpc3985 (
      {stage2_56[51]},
      {stage3_56[29]}
   );
   gpc1_1 gpc3986 (
      {stage2_56[52]},
      {stage3_56[30]}
   );
   gpc1_1 gpc3987 (
      {stage2_58[13]},
      {stage3_58[13]}
   );
   gpc1_1 gpc3988 (
      {stage2_58[14]},
      {stage3_58[14]}
   );
   gpc1_1 gpc3989 (
      {stage2_58[15]},
      {stage3_58[15]}
   );
   gpc1_1 gpc3990 (
      {stage2_58[16]},
      {stage3_58[16]}
   );
   gpc1_1 gpc3991 (
      {stage2_58[17]},
      {stage3_58[17]}
   );
   gpc1_1 gpc3992 (
      {stage2_58[18]},
      {stage3_58[18]}
   );
   gpc1_1 gpc3993 (
      {stage2_58[19]},
      {stage3_58[19]}
   );
   gpc1_1 gpc3994 (
      {stage2_58[20]},
      {stage3_58[20]}
   );
   gpc1_1 gpc3995 (
      {stage2_58[21]},
      {stage3_58[21]}
   );
   gpc1_1 gpc3996 (
      {stage2_58[22]},
      {stage3_58[22]}
   );
   gpc1_1 gpc3997 (
      {stage2_58[23]},
      {stage3_58[23]}
   );
   gpc1_1 gpc3998 (
      {stage2_58[24]},
      {stage3_58[24]}
   );
   gpc1_1 gpc3999 (
      {stage2_58[25]},
      {stage3_58[25]}
   );
   gpc1_1 gpc4000 (
      {stage2_58[26]},
      {stage3_58[26]}
   );
   gpc1_1 gpc4001 (
      {stage2_58[27]},
      {stage3_58[27]}
   );
   gpc1_1 gpc4002 (
      {stage2_58[28]},
      {stage3_58[28]}
   );
   gpc1_1 gpc4003 (
      {stage2_58[29]},
      {stage3_58[29]}
   );
   gpc1_1 gpc4004 (
      {stage2_58[30]},
      {stage3_58[30]}
   );
   gpc1_1 gpc4005 (
      {stage2_58[31]},
      {stage3_58[31]}
   );
   gpc1_1 gpc4006 (
      {stage2_58[32]},
      {stage3_58[32]}
   );
   gpc1_1 gpc4007 (
      {stage2_59[70]},
      {stage3_59[17]}
   );
   gpc1_1 gpc4008 (
      {stage2_59[71]},
      {stage3_59[18]}
   );
   gpc1_1 gpc4009 (
      {stage2_59[72]},
      {stage3_59[19]}
   );
   gpc1_1 gpc4010 (
      {stage2_59[73]},
      {stage3_59[20]}
   );
   gpc1_1 gpc4011 (
      {stage2_59[74]},
      {stage3_59[21]}
   );
   gpc1_1 gpc4012 (
      {stage2_59[75]},
      {stage3_59[22]}
   );
   gpc1_1 gpc4013 (
      {stage2_59[76]},
      {stage3_59[23]}
   );
   gpc1_1 gpc4014 (
      {stage2_59[77]},
      {stage3_59[24]}
   );
   gpc1_1 gpc4015 (
      {stage2_59[78]},
      {stage3_59[25]}
   );
   gpc1_1 gpc4016 (
      {stage2_59[79]},
      {stage3_59[26]}
   );
   gpc1_1 gpc4017 (
      {stage2_59[80]},
      {stage3_59[27]}
   );
   gpc1_1 gpc4018 (
      {stage2_61[59]},
      {stage3_61[17]}
   );
   gpc1_1 gpc4019 (
      {stage2_61[60]},
      {stage3_61[18]}
   );
   gpc1_1 gpc4020 (
      {stage2_61[61]},
      {stage3_61[19]}
   );
   gpc1_1 gpc4021 (
      {stage2_61[62]},
      {stage3_61[20]}
   );
   gpc1_1 gpc4022 (
      {stage2_61[63]},
      {stage3_61[21]}
   );
   gpc1_1 gpc4023 (
      {stage2_61[64]},
      {stage3_61[22]}
   );
   gpc1_1 gpc4024 (
      {stage2_61[65]},
      {stage3_61[23]}
   );
   gpc1_1 gpc4025 (
      {stage2_61[66]},
      {stage3_61[24]}
   );
   gpc1_1 gpc4026 (
      {stage2_64[29]},
      {stage3_64[12]}
   );
   gpc1_1 gpc4027 (
      {stage2_64[30]},
      {stage3_64[13]}
   );
   gpc1_1 gpc4028 (
      {stage2_64[31]},
      {stage3_64[14]}
   );
   gpc1_1 gpc4029 (
      {stage2_64[32]},
      {stage3_64[15]}
   );
   gpc1_1 gpc4030 (
      {stage2_64[33]},
      {stage3_64[16]}
   );
   gpc1_1 gpc4031 (
      {stage2_64[34]},
      {stage3_64[17]}
   );
   gpc1_1 gpc4032 (
      {stage2_64[35]},
      {stage3_64[18]}
   );
   gpc1_1 gpc4033 (
      {stage2_64[36]},
      {stage3_64[19]}
   );
   gpc1_1 gpc4034 (
      {stage2_64[37]},
      {stage3_64[20]}
   );
   gpc1_1 gpc4035 (
      {stage2_64[38]},
      {stage3_64[21]}
   );
   gpc1_1 gpc4036 (
      {stage2_64[39]},
      {stage3_64[22]}
   );
   gpc1_1 gpc4037 (
      {stage2_64[40]},
      {stage3_64[23]}
   );
   gpc1_1 gpc4038 (
      {stage2_64[41]},
      {stage3_64[24]}
   );
   gpc1_1 gpc4039 (
      {stage2_64[42]},
      {stage3_64[25]}
   );
   gpc1_1 gpc4040 (
      {stage2_64[43]},
      {stage3_64[26]}
   );
   gpc1_1 gpc4041 (
      {stage2_64[44]},
      {stage3_64[27]}
   );
   gpc1_1 gpc4042 (
      {stage2_64[45]},
      {stage3_64[28]}
   );
   gpc1_1 gpc4043 (
      {stage2_65[10]},
      {stage3_65[11]}
   );
   gpc1_1 gpc4044 (
      {stage2_65[11]},
      {stage3_65[12]}
   );
   gpc1_1 gpc4045 (
      {stage2_65[12]},
      {stage3_65[13]}
   );
   gpc1_1 gpc4046 (
      {stage2_67[0]},
      {stage3_67[3]}
   );
   gpc1_1 gpc4047 (
      {stage2_67[1]},
      {stage3_67[4]}
   );
   gpc1163_5 gpc4048 (
      {stage3_0[0], stage3_0[1], stage3_0[2]},
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_2[0]},
      {stage3_3[0]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc1163_5 gpc4049 (
      {stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_2[1]},
      {stage3_3[1]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1],stage4_0[1]}
   );
   gpc615_5 gpc4050 (
      {stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5], stage3_2[6]},
      {stage3_3[2]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[2],stage4_3[2],stage4_2[2]}
   );
   gpc606_5 gpc4051 (
      {stage3_3[3], stage3_3[4], stage3_3[5], stage3_3[6], stage3_3[7], stage3_3[8]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[3],stage4_3[3]}
   );
   gpc606_5 gpc4052 (
      {stage3_3[9], stage3_3[10], stage3_3[11], stage3_3[12], stage3_3[13], 1'b0},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[2],stage4_5[2],stage4_4[4],stage4_3[4]}
   );
   gpc615_5 gpc4053 (
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10]},
      {stage3_5[12]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[2],stage4_6[3],stage4_5[3],stage4_4[5]}
   );
   gpc615_5 gpc4054 (
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[3],stage4_6[4]}
   );
   gpc207_4 gpc4055 (
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage3_9[0], stage3_9[1]},
      {stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[4]}
   );
   gpc207_4 gpc4056 (
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12], stage3_7[13], stage3_7[14]},
      {stage3_9[2], stage3_9[3]},
      {stage4_10[2],stage4_9[2],stage4_8[3],stage4_7[5]}
   );
   gpc606_5 gpc4057 (
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[0],stage4_10[3],stage4_9[3],stage4_8[4]}
   );
   gpc2135_5 gpc4058 (
      {stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7], stage3_9[8]},
      {stage3_10[6], stage3_10[7], stage3_10[8]},
      {stage3_11[0]},
      {stage3_12[0], stage3_12[1]},
      {stage4_13[0],stage4_12[1],stage4_11[1],stage4_10[4],stage4_9[4]}
   );
   gpc606_5 gpc4059 (
      {stage3_9[9], stage3_9[10], stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14]},
      {stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5], stage3_11[6]},
      {stage4_13[1],stage4_12[2],stage4_11[2],stage4_10[5],stage4_9[5]}
   );
   gpc606_5 gpc4060 (
      {stage3_9[15], stage3_9[16], stage3_9[17], stage3_9[18], stage3_9[19], stage3_9[20]},
      {stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11], stage3_11[12]},
      {stage4_13[2],stage4_12[3],stage4_11[3],stage4_10[6],stage4_9[6]}
   );
   gpc2135_5 gpc4061 (
      {stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13]},
      {stage3_11[13], stage3_11[14], stage3_11[15]},
      {stage3_12[2]},
      {stage3_13[0], stage3_13[1]},
      {stage4_14[0],stage4_13[3],stage4_12[4],stage4_11[4],stage4_10[7]}
   );
   gpc207_4 gpc4062 (
      {stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9]},
      {stage3_14[0], stage3_14[1]},
      {stage4_15[0],stage4_14[1],stage4_13[4],stage4_12[5]}
   );
   gpc207_4 gpc4063 (
      {stage3_12[10], stage3_12[11], stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16]},
      {stage3_14[2], stage3_14[3]},
      {stage4_15[1],stage4_14[2],stage4_13[5],stage4_12[6]}
   );
   gpc606_5 gpc4064 (
      {stage3_12[17], stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22]},
      {stage3_14[4], stage3_14[5], stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9]},
      {stage4_16[0],stage4_15[2],stage4_14[3],stage4_13[6],stage4_12[7]}
   );
   gpc606_5 gpc4065 (
      {stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[3],stage4_14[4],stage4_13[7]}
   );
   gpc606_5 gpc4066 (
      {stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[2],stage4_15[4],stage4_14[5],stage4_13[8]}
   );
   gpc606_5 gpc4067 (
      {stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19]},
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17]},
      {stage4_17[2],stage4_16[3],stage4_15[5],stage4_14[6],stage4_13[9]}
   );
   gpc117_4 gpc4068 (
      {stage3_14[10], stage3_14[11], stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16]},
      {stage3_15[18]},
      {stage3_16[0]},
      {stage4_17[3],stage4_16[4],stage4_15[6],stage4_14[7]}
   );
   gpc117_4 gpc4069 (
      {stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage3_15[19]},
      {stage3_16[1]},
      {stage4_17[4],stage4_16[5],stage4_15[7],stage4_14[8]}
   );
   gpc117_4 gpc4070 (
      {stage3_14[24], stage3_14[25], stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29], stage3_14[30]},
      {stage3_15[20]},
      {stage3_16[2]},
      {stage4_17[5],stage4_16[6],stage4_15[8],stage4_14[9]}
   );
   gpc117_4 gpc4071 (
      {stage3_14[31], stage3_14[32], stage3_14[33], stage3_14[34], stage3_14[35], 1'b0, 1'b0},
      {stage3_15[21]},
      {stage3_16[3]},
      {stage4_17[6],stage4_16[7],stage4_15[9],stage4_14[10]}
   );
   gpc615_5 gpc4072 (
      {stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25], stage3_15[26]},
      {stage3_16[4]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[0],stage4_17[7],stage4_16[8],stage4_15[10]}
   );
   gpc615_5 gpc4073 (
      {stage3_15[27], stage3_15[28], stage3_15[29], stage3_15[30], stage3_15[31]},
      {stage3_16[5]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[1],stage4_17[8],stage4_16[9],stage4_15[11]}
   );
   gpc606_5 gpc4074 (
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[2],stage4_18[2],stage4_17[9],stage4_16[10]}
   );
   gpc606_5 gpc4075 (
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[3],stage4_18[3],stage4_17[10],stage4_16[11]}
   );
   gpc606_5 gpc4076 (
      {stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], 1'b0, 1'b0},
      {stage3_18[12], stage3_18[13], stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17]},
      {stage4_20[2],stage4_19[4],stage4_18[4],stage4_17[11],stage4_16[12]}
   );
   gpc615_5 gpc4077 (
      {stage3_18[18], stage3_18[19], stage3_18[20], stage3_18[21], stage3_18[22]},
      {stage3_19[0]},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage4_22[0],stage4_21[0],stage4_20[3],stage4_19[5],stage4_18[5]}
   );
   gpc615_5 gpc4078 (
      {stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage3_20[6]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[1],stage4_21[1],stage4_20[4],stage4_19[6]}
   );
   gpc615_5 gpc4079 (
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10]},
      {stage3_20[7]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[2],stage4_21[2],stage4_20[5],stage4_19[7]}
   );
   gpc615_5 gpc4080 (
      {stage3_19[11], stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15]},
      {stage3_20[8]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[3],stage4_21[3],stage4_20[6],stage4_19[8]}
   );
   gpc615_5 gpc4081 (
      {stage3_19[16], stage3_19[17], stage3_19[18], stage3_19[19], stage3_19[20]},
      {stage3_20[9]},
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage4_23[3],stage4_22[4],stage4_21[4],stage4_20[7],stage4_19[9]}
   );
   gpc606_5 gpc4082 (
      {stage3_20[10], stage3_20[11], stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[4],stage4_22[5],stage4_21[5],stage4_20[8]}
   );
   gpc606_5 gpc4083 (
      {stage3_20[16], stage3_20[17], stage3_20[18], stage3_20[19], stage3_20[20], stage3_20[21]},
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10], stage3_22[11]},
      {stage4_24[1],stage4_23[5],stage4_22[6],stage4_21[6],stage4_20[9]}
   );
   gpc615_5 gpc4084 (
      {stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15], stage3_22[16]},
      {stage3_23[0]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[0],stage4_24[2],stage4_23[6],stage4_22[7]}
   );
   gpc615_5 gpc4085 (
      {stage3_22[17], stage3_22[18], stage3_22[19], stage3_22[20], stage3_22[21]},
      {stage3_23[1]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[1],stage4_24[3],stage4_23[7],stage4_22[8]}
   );
   gpc615_5 gpc4086 (
      {stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5], stage3_23[6]},
      {stage3_24[12]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[2],stage4_25[2],stage4_24[4],stage4_23[8]}
   );
   gpc615_5 gpc4087 (
      {stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage3_24[13]},
      {stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage4_27[1],stage4_26[3],stage4_25[3],stage4_24[5],stage4_23[9]}
   );
   gpc615_5 gpc4088 (
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16]},
      {stage3_26[0]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[2],stage4_26[4],stage4_25[4]}
   );
   gpc615_5 gpc4089 (
      {stage3_25[17], stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21]},
      {stage3_26[1]},
      {stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage4_29[1],stage4_28[1],stage4_27[3],stage4_26[5],stage4_25[5]}
   );
   gpc117_4 gpc4090 (
      {stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5], stage3_26[6], stage3_26[7], stage3_26[8]},
      {stage3_27[12]},
      {stage3_28[0]},
      {stage4_29[2],stage4_28[2],stage4_27[4],stage4_26[6]}
   );
   gpc207_4 gpc4091 (
      {stage3_26[9], stage3_26[10], stage3_26[11], stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15]},
      {stage3_28[1], stage3_28[2]},
      {stage4_29[3],stage4_28[3],stage4_27[5],stage4_26[7]}
   );
   gpc606_5 gpc4092 (
      {stage3_27[13], stage3_27[14], stage3_27[15], stage3_27[16], stage3_27[17], stage3_27[18]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[0],stage4_29[4],stage4_28[4],stage4_27[6]}
   );
   gpc606_5 gpc4093 (
      {stage3_28[3], stage3_28[4], stage3_28[5], stage3_28[6], stage3_28[7], stage3_28[8]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[1],stage4_30[1],stage4_29[5],stage4_28[5]}
   );
   gpc606_5 gpc4094 (
      {stage3_28[9], stage3_28[10], stage3_28[11], stage3_28[12], stage3_28[13], stage3_28[14]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[2],stage4_30[2],stage4_29[6],stage4_28[6]}
   );
   gpc606_5 gpc4095 (
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[2],stage4_31[3],stage4_30[3],stage4_29[7]}
   );
   gpc606_5 gpc4096 (
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11]},
      {stage4_33[1],stage4_32[3],stage4_31[4],stage4_30[4],stage4_29[8]}
   );
   gpc606_5 gpc4097 (
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17]},
      {stage4_33[2],stage4_32[4],stage4_31[5],stage4_30[5],stage4_29[9]}
   );
   gpc615_5 gpc4098 (
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16]},
      {stage3_31[18]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[3],stage4_32[5],stage4_31[6],stage4_30[6]}
   );
   gpc606_5 gpc4099 (
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[0],stage4_34[1],stage4_33[4],stage4_32[6]}
   );
   gpc606_5 gpc4100 (
      {stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15], stage3_32[16], stage3_32[17]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage4_36[1],stage4_35[1],stage4_34[2],stage4_33[5],stage4_32[7]}
   );
   gpc606_5 gpc4101 (
      {stage3_32[18], stage3_32[19], stage3_32[20], stage3_32[21], stage3_32[22], stage3_32[23]},
      {stage3_34[12], stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage4_36[2],stage4_35[2],stage4_34[3],stage4_33[6],stage4_32[8]}
   );
   gpc606_5 gpc4102 (
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[3],stage4_35[3],stage4_34[4],stage4_33[7]}
   );
   gpc606_5 gpc4103 (
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage3_35[6], stage3_35[7], stage3_35[8], stage3_35[9], stage3_35[10], stage3_35[11]},
      {stage4_37[1],stage4_36[4],stage4_35[4],stage4_34[5],stage4_33[8]}
   );
   gpc1343_5 gpc4104 (
      {stage3_35[12], stage3_35[13], stage3_35[14]},
      {stage3_36[0], stage3_36[1], stage3_36[2], stage3_36[3]},
      {stage3_37[0], stage3_37[1], stage3_37[2]},
      {stage3_38[0]},
      {stage4_39[0],stage4_38[0],stage4_37[2],stage4_36[5],stage4_35[5]}
   );
   gpc1343_5 gpc4105 (
      {stage3_35[15], stage3_35[16], stage3_35[17]},
      {stage3_36[4], stage3_36[5], stage3_36[6], stage3_36[7]},
      {stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage3_38[1]},
      {stage4_39[1],stage4_38[1],stage4_37[3],stage4_36[6],stage4_35[6]}
   );
   gpc1343_5 gpc4106 (
      {stage3_35[18], stage3_35[19], stage3_35[20]},
      {stage3_36[8], stage3_36[9], stage3_36[10], stage3_36[11]},
      {stage3_37[6], stage3_37[7], stage3_37[8]},
      {stage3_38[2]},
      {stage4_39[2],stage4_38[2],stage4_37[4],stage4_36[7],stage4_35[7]}
   );
   gpc1343_5 gpc4107 (
      {stage3_35[21], stage3_35[22], stage3_35[23]},
      {stage3_36[12], stage3_36[13], stage3_36[14], stage3_36[15]},
      {stage3_37[9], stage3_37[10], stage3_37[11]},
      {stage3_38[3]},
      {stage4_39[3],stage4_38[3],stage4_37[5],stage4_36[8],stage4_35[8]}
   );
   gpc615_5 gpc4108 (
      {stage3_38[4], stage3_38[5], stage3_38[6], stage3_38[7], stage3_38[8]},
      {stage3_39[0]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[0],stage4_40[0],stage4_39[4],stage4_38[4]}
   );
   gpc615_5 gpc4109 (
      {stage3_38[9], stage3_38[10], stage3_38[11], stage3_38[12], stage3_38[13]},
      {stage3_39[1]},
      {stage3_40[6], stage3_40[7], stage3_40[8], stage3_40[9], stage3_40[10], stage3_40[11]},
      {stage4_42[1],stage4_41[1],stage4_40[1],stage4_39[5],stage4_38[5]}
   );
   gpc117_4 gpc4110 (
      {stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5], stage3_39[6], stage3_39[7], stage3_39[8]},
      {stage3_40[12]},
      {stage3_41[0]},
      {stage4_42[2],stage4_41[2],stage4_40[2],stage4_39[6]}
   );
   gpc117_4 gpc4111 (
      {stage3_39[9], stage3_39[10], stage3_39[11], stage3_39[12], stage3_39[13], stage3_39[14], stage3_39[15]},
      {stage3_40[13]},
      {stage3_41[1]},
      {stage4_42[3],stage4_41[3],stage4_40[3],stage4_39[7]}
   );
   gpc117_4 gpc4112 (
      {stage3_39[16], stage3_39[17], stage3_39[18], stage3_39[19], stage3_39[20], stage3_39[21], stage3_39[22]},
      {stage3_40[14]},
      {stage3_41[2]},
      {stage4_42[4],stage4_41[4],stage4_40[4],stage4_39[8]}
   );
   gpc606_5 gpc4113 (
      {stage3_41[3], stage3_41[4], stage3_41[5], stage3_41[6], stage3_41[7], stage3_41[8]},
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4], stage3_43[5]},
      {stage4_45[0],stage4_44[0],stage4_43[0],stage4_42[5],stage4_41[5]}
   );
   gpc606_5 gpc4114 (
      {stage3_41[9], stage3_41[10], stage3_41[11], stage3_41[12], stage3_41[13], stage3_41[14]},
      {stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9], stage3_43[10], stage3_43[11]},
      {stage4_45[1],stage4_44[1],stage4_43[1],stage4_42[6],stage4_41[6]}
   );
   gpc615_5 gpc4115 (
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4]},
      {stage3_43[12]},
      {stage3_44[0], stage3_44[1], stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5]},
      {stage4_46[0],stage4_45[2],stage4_44[2],stage4_43[2],stage4_42[7]}
   );
   gpc615_5 gpc4116 (
      {stage3_42[5], stage3_42[6], stage3_42[7], stage3_42[8], stage3_42[9]},
      {stage3_43[13]},
      {stage3_44[6], stage3_44[7], stage3_44[8], stage3_44[9], stage3_44[10], stage3_44[11]},
      {stage4_46[1],stage4_45[3],stage4_44[3],stage4_43[3],stage4_42[8]}
   );
   gpc615_5 gpc4117 (
      {stage3_42[10], stage3_42[11], stage3_42[12], stage3_42[13], stage3_42[14]},
      {stage3_43[14]},
      {stage3_44[12], stage3_44[13], stage3_44[14], stage3_44[15], stage3_44[16], stage3_44[17]},
      {stage4_46[2],stage4_45[4],stage4_44[4],stage4_43[4],stage4_42[9]}
   );
   gpc615_5 gpc4118 (
      {stage3_42[15], stage3_42[16], stage3_42[17], stage3_42[18], stage3_42[19]},
      {stage3_43[15]},
      {stage3_44[18], stage3_44[19], stage3_44[20], stage3_44[21], stage3_44[22], stage3_44[23]},
      {stage4_46[3],stage4_45[5],stage4_44[5],stage4_43[5],stage4_42[10]}
   );
   gpc615_5 gpc4119 (
      {stage3_43[16], stage3_43[17], stage3_43[18], stage3_43[19], stage3_43[20]},
      {stage3_44[24]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[4],stage4_45[6],stage4_44[6],stage4_43[6]}
   );
   gpc606_5 gpc4120 (
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9], stage3_45[10], stage3_45[11]},
      {stage3_47[0], stage3_47[1], stage3_47[2], stage3_47[3], stage3_47[4], stage3_47[5]},
      {stage4_49[0],stage4_48[0],stage4_47[1],stage4_46[5],stage4_45[7]}
   );
   gpc606_5 gpc4121 (
      {stage3_45[12], stage3_45[13], stage3_45[14], stage3_45[15], stage3_45[16], stage3_45[17]},
      {stage3_47[6], stage3_47[7], stage3_47[8], stage3_47[9], stage3_47[10], stage3_47[11]},
      {stage4_49[1],stage4_48[1],stage4_47[2],stage4_46[6],stage4_45[8]}
   );
   gpc207_4 gpc4122 (
      {stage3_46[0], stage3_46[1], stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5], stage3_46[6]},
      {stage3_48[0], stage3_48[1]},
      {stage4_49[2],stage4_48[2],stage4_47[3],stage4_46[7]}
   );
   gpc606_5 gpc4123 (
      {stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5], stage3_48[6], stage3_48[7]},
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5]},
      {stage4_52[0],stage4_51[0],stage4_50[0],stage4_49[3],stage4_48[3]}
   );
   gpc606_5 gpc4124 (
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5]},
      {stage3_51[0], stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage4_53[0],stage4_52[1],stage4_51[1],stage4_50[1],stage4_49[4]}
   );
   gpc7_3 gpc4125 (
      {stage3_50[6], stage3_50[7], stage3_50[8], stage3_50[9], stage3_50[10], stage3_50[11], stage3_50[12]},
      {stage4_52[2],stage4_51[2],stage4_50[2]}
   );
   gpc606_5 gpc4126 (
      {stage3_50[13], stage3_50[14], stage3_50[15], stage3_50[16], stage3_50[17], stage3_50[18]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[1],stage4_52[3],stage4_51[3],stage4_50[3]}
   );
   gpc606_5 gpc4127 (
      {stage3_50[19], stage3_50[20], stage3_50[21], stage3_50[22], stage3_50[23], stage3_50[24]},
      {stage3_52[6], stage3_52[7], stage3_52[8], stage3_52[9], stage3_52[10], stage3_52[11]},
      {stage4_54[1],stage4_53[2],stage4_52[4],stage4_51[4],stage4_50[4]}
   );
   gpc606_5 gpc4128 (
      {stage3_50[25], stage3_50[26], stage3_50[27], stage3_50[28], stage3_50[29], stage3_50[30]},
      {stage3_52[12], stage3_52[13], stage3_52[14], stage3_52[15], stage3_52[16], stage3_52[17]},
      {stage4_54[2],stage4_53[3],stage4_52[5],stage4_51[5],stage4_50[5]}
   );
   gpc606_5 gpc4129 (
      {stage3_51[6], stage3_51[7], stage3_51[8], stage3_51[9], stage3_51[10], stage3_51[11]},
      {stage3_53[0], stage3_53[1], stage3_53[2], stage3_53[3], stage3_53[4], stage3_53[5]},
      {stage4_55[0],stage4_54[3],stage4_53[4],stage4_52[6],stage4_51[6]}
   );
   gpc615_5 gpc4130 (
      {stage3_52[18], stage3_52[19], stage3_52[20], stage3_52[21], stage3_52[22]},
      {stage3_53[6]},
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage4_56[0],stage4_55[1],stage4_54[4],stage4_53[5],stage4_52[7]}
   );
   gpc606_5 gpc4131 (
      {stage3_54[6], stage3_54[7], stage3_54[8], stage3_54[9], stage3_54[10], stage3_54[11]},
      {stage3_56[0], stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5]},
      {stage4_58[0],stage4_57[0],stage4_56[1],stage4_55[2],stage4_54[5]}
   );
   gpc615_5 gpc4132 (
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3], stage3_55[4]},
      {stage3_56[6]},
      {stage3_57[0], stage3_57[1], stage3_57[2], stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage4_59[0],stage4_58[1],stage4_57[1],stage4_56[2],stage4_55[3]}
   );
   gpc606_5 gpc4133 (
      {stage3_56[7], stage3_56[8], stage3_56[9], stage3_56[10], stage3_56[11], stage3_56[12]},
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5]},
      {stage4_60[0],stage4_59[1],stage4_58[2],stage4_57[2],stage4_56[3]}
   );
   gpc606_5 gpc4134 (
      {stage3_56[13], stage3_56[14], stage3_56[15], stage3_56[16], stage3_56[17], stage3_56[18]},
      {stage3_58[6], stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10], stage3_58[11]},
      {stage4_60[1],stage4_59[2],stage4_58[3],stage4_57[3],stage4_56[4]}
   );
   gpc615_5 gpc4135 (
      {stage3_56[19], stage3_56[20], stage3_56[21], stage3_56[22], stage3_56[23]},
      {stage3_57[6]},
      {stage3_58[12], stage3_58[13], stage3_58[14], stage3_58[15], stage3_58[16], stage3_58[17]},
      {stage4_60[2],stage4_59[3],stage4_58[4],stage4_57[4],stage4_56[5]}
   );
   gpc606_5 gpc4136 (
      {stage3_57[7], stage3_57[8], stage3_57[9], stage3_57[10], stage3_57[11], stage3_57[12]},
      {stage3_59[0], stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5]},
      {stage4_61[0],stage4_60[3],stage4_59[4],stage4_58[5],stage4_57[5]}
   );
   gpc606_5 gpc4137 (
      {stage3_59[6], stage3_59[7], stage3_59[8], stage3_59[9], stage3_59[10], stage3_59[11]},
      {stage3_61[0], stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5]},
      {stage4_63[0],stage4_62[0],stage4_61[1],stage4_60[4],stage4_59[5]}
   );
   gpc606_5 gpc4138 (
      {stage3_59[12], stage3_59[13], stage3_59[14], stage3_59[15], stage3_59[16], stage3_59[17]},
      {stage3_61[6], stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11]},
      {stage4_63[1],stage4_62[1],stage4_61[2],stage4_60[5],stage4_59[6]}
   );
   gpc606_5 gpc4139 (
      {stage3_60[0], stage3_60[1], stage3_60[2], stage3_60[3], stage3_60[4], stage3_60[5]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], stage3_62[5]},
      {stage4_64[0],stage4_63[2],stage4_62[2],stage4_61[3],stage4_60[6]}
   );
   gpc606_5 gpc4140 (
      {stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9], stage3_62[10], stage3_62[11]},
      {stage3_64[0], stage3_64[1], stage3_64[2], stage3_64[3], stage3_64[4], stage3_64[5]},
      {stage4_66[0],stage4_65[0],stage4_64[1],stage4_63[3],stage4_62[3]}
   );
   gpc606_5 gpc4141 (
      {stage3_62[12], stage3_62[13], stage3_62[14], stage3_62[15], stage3_62[16], stage3_62[17]},
      {stage3_64[6], stage3_64[7], stage3_64[8], stage3_64[9], stage3_64[10], stage3_64[11]},
      {stage4_66[1],stage4_65[1],stage4_64[2],stage4_63[4],stage4_62[4]}
   );
   gpc606_5 gpc4142 (
      {stage3_63[0], stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[2],stage4_65[2],stage4_64[3],stage4_63[5]}
   );
   gpc606_5 gpc4143 (
      {stage3_63[6], stage3_63[7], stage3_63[8], stage3_63[9], stage3_63[10], stage3_63[11]},
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage4_67[1],stage4_66[3],stage4_65[3],stage4_64[4],stage4_63[6]}
   );
   gpc1_1 gpc4144 (
      {stage3_0[6]},
      {stage4_0[2]}
   );
   gpc1_1 gpc4145 (
      {stage3_0[7]},
      {stage4_0[3]}
   );
   gpc1_1 gpc4146 (
      {stage3_1[12]},
      {stage4_1[2]}
   );
   gpc1_1 gpc4147 (
      {stage3_1[13]},
      {stage4_1[3]}
   );
   gpc1_1 gpc4148 (
      {stage3_2[7]},
      {stage4_2[3]}
   );
   gpc1_1 gpc4149 (
      {stage3_2[8]},
      {stage4_2[4]}
   );
   gpc1_1 gpc4150 (
      {stage3_2[9]},
      {stage4_2[5]}
   );
   gpc1_1 gpc4151 (
      {stage3_2[10]},
      {stage4_2[6]}
   );
   gpc1_1 gpc4152 (
      {stage3_4[11]},
      {stage4_4[6]}
   );
   gpc1_1 gpc4153 (
      {stage3_4[12]},
      {stage4_4[7]}
   );
   gpc1_1 gpc4154 (
      {stage3_4[13]},
      {stage4_4[8]}
   );
   gpc1_1 gpc4155 (
      {stage3_5[13]},
      {stage4_5[4]}
   );
   gpc1_1 gpc4156 (
      {stage3_5[14]},
      {stage4_5[5]}
   );
   gpc1_1 gpc4157 (
      {stage3_5[15]},
      {stage4_5[6]}
   );
   gpc1_1 gpc4158 (
      {stage3_5[16]},
      {stage4_5[7]}
   );
   gpc1_1 gpc4159 (
      {stage3_5[17]},
      {stage4_5[8]}
   );
   gpc1_1 gpc4160 (
      {stage3_6[11]},
      {stage4_6[5]}
   );
   gpc1_1 gpc4161 (
      {stage3_6[12]},
      {stage4_6[6]}
   );
   gpc1_1 gpc4162 (
      {stage3_6[13]},
      {stage4_6[7]}
   );
   gpc1_1 gpc4163 (
      {stage3_6[14]},
      {stage4_6[8]}
   );
   gpc1_1 gpc4164 (
      {stage3_6[15]},
      {stage4_6[9]}
   );
   gpc1_1 gpc4165 (
      {stage3_6[16]},
      {stage4_6[10]}
   );
   gpc1_1 gpc4166 (
      {stage3_6[17]},
      {stage4_6[11]}
   );
   gpc1_1 gpc4167 (
      {stage3_6[18]},
      {stage4_6[12]}
   );
   gpc1_1 gpc4168 (
      {stage3_6[19]},
      {stage4_6[13]}
   );
   gpc1_1 gpc4169 (
      {stage3_7[15]},
      {stage4_7[6]}
   );
   gpc1_1 gpc4170 (
      {stage3_7[16]},
      {stage4_7[7]}
   );
   gpc1_1 gpc4171 (
      {stage3_8[12]},
      {stage4_8[5]}
   );
   gpc1_1 gpc4172 (
      {stage3_8[13]},
      {stage4_8[6]}
   );
   gpc1_1 gpc4173 (
      {stage3_8[14]},
      {stage4_8[7]}
   );
   gpc1_1 gpc4174 (
      {stage3_8[15]},
      {stage4_8[8]}
   );
   gpc1_1 gpc4175 (
      {stage3_8[16]},
      {stage4_8[9]}
   );
   gpc1_1 gpc4176 (
      {stage3_10[14]},
      {stage4_10[8]}
   );
   gpc1_1 gpc4177 (
      {stage3_11[16]},
      {stage4_11[5]}
   );
   gpc1_1 gpc4178 (
      {stage3_11[17]},
      {stage4_11[6]}
   );
   gpc1_1 gpc4179 (
      {stage3_12[23]},
      {stage4_12[8]}
   );
   gpc1_1 gpc4180 (
      {stage3_15[32]},
      {stage4_15[12]}
   );
   gpc1_1 gpc4181 (
      {stage3_15[33]},
      {stage4_15[13]}
   );
   gpc1_1 gpc4182 (
      {stage3_15[34]},
      {stage4_15[14]}
   );
   gpc1_1 gpc4183 (
      {stage3_15[35]},
      {stage4_15[15]}
   );
   gpc1_1 gpc4184 (
      {stage3_15[36]},
      {stage4_15[16]}
   );
   gpc1_1 gpc4185 (
      {stage3_17[12]},
      {stage4_17[12]}
   );
   gpc1_1 gpc4186 (
      {stage3_17[13]},
      {stage4_17[13]}
   );
   gpc1_1 gpc4187 (
      {stage3_17[14]},
      {stage4_17[14]}
   );
   gpc1_1 gpc4188 (
      {stage3_17[15]},
      {stage4_17[15]}
   );
   gpc1_1 gpc4189 (
      {stage3_17[16]},
      {stage4_17[16]}
   );
   gpc1_1 gpc4190 (
      {stage3_19[21]},
      {stage4_19[10]}
   );
   gpc1_1 gpc4191 (
      {stage3_19[22]},
      {stage4_19[11]}
   );
   gpc1_1 gpc4192 (
      {stage3_19[23]},
      {stage4_19[12]}
   );
   gpc1_1 gpc4193 (
      {stage3_19[24]},
      {stage4_19[13]}
   );
   gpc1_1 gpc4194 (
      {stage3_19[25]},
      {stage4_19[14]}
   );
   gpc1_1 gpc4195 (
      {stage3_19[26]},
      {stage4_19[15]}
   );
   gpc1_1 gpc4196 (
      {stage3_20[22]},
      {stage4_20[10]}
   );
   gpc1_1 gpc4197 (
      {stage3_21[24]},
      {stage4_21[7]}
   );
   gpc1_1 gpc4198 (
      {stage3_22[22]},
      {stage4_22[9]}
   );
   gpc1_1 gpc4199 (
      {stage3_22[23]},
      {stage4_22[10]}
   );
   gpc1_1 gpc4200 (
      {stage3_22[24]},
      {stage4_22[11]}
   );
   gpc1_1 gpc4201 (
      {stage3_22[25]},
      {stage4_22[12]}
   );
   gpc1_1 gpc4202 (
      {stage3_22[26]},
      {stage4_22[13]}
   );
   gpc1_1 gpc4203 (
      {stage3_24[14]},
      {stage4_24[6]}
   );
   gpc1_1 gpc4204 (
      {stage3_24[15]},
      {stage4_24[7]}
   );
   gpc1_1 gpc4205 (
      {stage3_24[16]},
      {stage4_24[8]}
   );
   gpc1_1 gpc4206 (
      {stage3_24[17]},
      {stage4_24[9]}
   );
   gpc1_1 gpc4207 (
      {stage3_24[18]},
      {stage4_24[10]}
   );
   gpc1_1 gpc4208 (
      {stage3_24[19]},
      {stage4_24[11]}
   );
   gpc1_1 gpc4209 (
      {stage3_24[20]},
      {stage4_24[12]}
   );
   gpc1_1 gpc4210 (
      {stage3_24[21]},
      {stage4_24[13]}
   );
   gpc1_1 gpc4211 (
      {stage3_24[22]},
      {stage4_24[14]}
   );
   gpc1_1 gpc4212 (
      {stage3_24[23]},
      {stage4_24[15]}
   );
   gpc1_1 gpc4213 (
      {stage3_24[24]},
      {stage4_24[16]}
   );
   gpc1_1 gpc4214 (
      {stage3_24[25]},
      {stage4_24[17]}
   );
   gpc1_1 gpc4215 (
      {stage3_28[15]},
      {stage4_28[7]}
   );
   gpc1_1 gpc4216 (
      {stage3_28[16]},
      {stage4_28[8]}
   );
   gpc1_1 gpc4217 (
      {stage3_28[17]},
      {stage4_28[9]}
   );
   gpc1_1 gpc4218 (
      {stage3_28[18]},
      {stage4_28[10]}
   );
   gpc1_1 gpc4219 (
      {stage3_28[19]},
      {stage4_28[11]}
   );
   gpc1_1 gpc4220 (
      {stage3_30[17]},
      {stage4_30[7]}
   );
   gpc1_1 gpc4221 (
      {stage3_30[18]},
      {stage4_30[8]}
   );
   gpc1_1 gpc4222 (
      {stage3_30[19]},
      {stage4_30[9]}
   );
   gpc1_1 gpc4223 (
      {stage3_30[20]},
      {stage4_30[10]}
   );
   gpc1_1 gpc4224 (
      {stage3_30[21]},
      {stage4_30[11]}
   );
   gpc1_1 gpc4225 (
      {stage3_30[22]},
      {stage4_30[12]}
   );
   gpc1_1 gpc4226 (
      {stage3_30[23]},
      {stage4_30[13]}
   );
   gpc1_1 gpc4227 (
      {stage3_30[24]},
      {stage4_30[14]}
   );
   gpc1_1 gpc4228 (
      {stage3_30[25]},
      {stage4_30[15]}
   );
   gpc1_1 gpc4229 (
      {stage3_31[19]},
      {stage4_31[7]}
   );
   gpc1_1 gpc4230 (
      {stage3_31[20]},
      {stage4_31[8]}
   );
   gpc1_1 gpc4231 (
      {stage3_32[24]},
      {stage4_32[9]}
   );
   gpc1_1 gpc4232 (
      {stage3_32[25]},
      {stage4_32[10]}
   );
   gpc1_1 gpc4233 (
      {stage3_32[26]},
      {stage4_32[11]}
   );
   gpc1_1 gpc4234 (
      {stage3_32[27]},
      {stage4_32[12]}
   );
   gpc1_1 gpc4235 (
      {stage3_32[28]},
      {stage4_32[13]}
   );
   gpc1_1 gpc4236 (
      {stage3_32[29]},
      {stage4_32[14]}
   );
   gpc1_1 gpc4237 (
      {stage3_32[30]},
      {stage4_32[15]}
   );
   gpc1_1 gpc4238 (
      {stage3_32[31]},
      {stage4_32[16]}
   );
   gpc1_1 gpc4239 (
      {stage3_32[32]},
      {stage4_32[17]}
   );
   gpc1_1 gpc4240 (
      {stage3_32[33]},
      {stage4_32[18]}
   );
   gpc1_1 gpc4241 (
      {stage3_32[34]},
      {stage4_32[19]}
   );
   gpc1_1 gpc4242 (
      {stage3_33[12]},
      {stage4_33[9]}
   );
   gpc1_1 gpc4243 (
      {stage3_33[13]},
      {stage4_33[10]}
   );
   gpc1_1 gpc4244 (
      {stage3_33[14]},
      {stage4_33[11]}
   );
   gpc1_1 gpc4245 (
      {stage3_34[18]},
      {stage4_34[6]}
   );
   gpc1_1 gpc4246 (
      {stage3_34[19]},
      {stage4_34[7]}
   );
   gpc1_1 gpc4247 (
      {stage3_34[20]},
      {stage4_34[8]}
   );
   gpc1_1 gpc4248 (
      {stage3_34[21]},
      {stage4_34[9]}
   );
   gpc1_1 gpc4249 (
      {stage3_34[22]},
      {stage4_34[10]}
   );
   gpc1_1 gpc4250 (
      {stage3_35[24]},
      {stage4_35[9]}
   );
   gpc1_1 gpc4251 (
      {stage3_35[25]},
      {stage4_35[10]}
   );
   gpc1_1 gpc4252 (
      {stage3_36[16]},
      {stage4_36[9]}
   );
   gpc1_1 gpc4253 (
      {stage3_39[23]},
      {stage4_39[9]}
   );
   gpc1_1 gpc4254 (
      {stage3_40[15]},
      {stage4_40[5]}
   );
   gpc1_1 gpc4255 (
      {stage3_40[16]},
      {stage4_40[6]}
   );
   gpc1_1 gpc4256 (
      {stage3_40[17]},
      {stage4_40[7]}
   );
   gpc1_1 gpc4257 (
      {stage3_40[18]},
      {stage4_40[8]}
   );
   gpc1_1 gpc4258 (
      {stage3_40[19]},
      {stage4_40[9]}
   );
   gpc1_1 gpc4259 (
      {stage3_40[20]},
      {stage4_40[10]}
   );
   gpc1_1 gpc4260 (
      {stage3_40[21]},
      {stage4_40[11]}
   );
   gpc1_1 gpc4261 (
      {stage3_40[22]},
      {stage4_40[12]}
   );
   gpc1_1 gpc4262 (
      {stage3_40[23]},
      {stage4_40[13]}
   );
   gpc1_1 gpc4263 (
      {stage3_41[15]},
      {stage4_41[7]}
   );
   gpc1_1 gpc4264 (
      {stage3_41[16]},
      {stage4_41[8]}
   );
   gpc1_1 gpc4265 (
      {stage3_41[17]},
      {stage4_41[9]}
   );
   gpc1_1 gpc4266 (
      {stage3_41[18]},
      {stage4_41[10]}
   );
   gpc1_1 gpc4267 (
      {stage3_41[19]},
      {stage4_41[11]}
   );
   gpc1_1 gpc4268 (
      {stage3_41[20]},
      {stage4_41[12]}
   );
   gpc1_1 gpc4269 (
      {stage3_41[21]},
      {stage4_41[13]}
   );
   gpc1_1 gpc4270 (
      {stage3_41[22]},
      {stage4_41[14]}
   );
   gpc1_1 gpc4271 (
      {stage3_41[23]},
      {stage4_41[15]}
   );
   gpc1_1 gpc4272 (
      {stage3_41[24]},
      {stage4_41[16]}
   );
   gpc1_1 gpc4273 (
      {stage3_42[20]},
      {stage4_42[11]}
   );
   gpc1_1 gpc4274 (
      {stage3_42[21]},
      {stage4_42[12]}
   );
   gpc1_1 gpc4275 (
      {stage3_42[22]},
      {stage4_42[13]}
   );
   gpc1_1 gpc4276 (
      {stage3_42[23]},
      {stage4_42[14]}
   );
   gpc1_1 gpc4277 (
      {stage3_42[24]},
      {stage4_42[15]}
   );
   gpc1_1 gpc4278 (
      {stage3_42[25]},
      {stage4_42[16]}
   );
   gpc1_1 gpc4279 (
      {stage3_44[25]},
      {stage4_44[7]}
   );
   gpc1_1 gpc4280 (
      {stage3_44[26]},
      {stage4_44[8]}
   );
   gpc1_1 gpc4281 (
      {stage3_44[27]},
      {stage4_44[9]}
   );
   gpc1_1 gpc4282 (
      {stage3_44[28]},
      {stage4_44[10]}
   );
   gpc1_1 gpc4283 (
      {stage3_44[29]},
      {stage4_44[11]}
   );
   gpc1_1 gpc4284 (
      {stage3_44[30]},
      {stage4_44[12]}
   );
   gpc1_1 gpc4285 (
      {stage3_46[7]},
      {stage4_46[8]}
   );
   gpc1_1 gpc4286 (
      {stage3_46[8]},
      {stage4_46[9]}
   );
   gpc1_1 gpc4287 (
      {stage3_46[9]},
      {stage4_46[10]}
   );
   gpc1_1 gpc4288 (
      {stage3_46[10]},
      {stage4_46[11]}
   );
   gpc1_1 gpc4289 (
      {stage3_46[11]},
      {stage4_46[12]}
   );
   gpc1_1 gpc4290 (
      {stage3_46[12]},
      {stage4_46[13]}
   );
   gpc1_1 gpc4291 (
      {stage3_46[13]},
      {stage4_46[14]}
   );
   gpc1_1 gpc4292 (
      {stage3_46[14]},
      {stage4_46[15]}
   );
   gpc1_1 gpc4293 (
      {stage3_46[15]},
      {stage4_46[16]}
   );
   gpc1_1 gpc4294 (
      {stage3_46[16]},
      {stage4_46[17]}
   );
   gpc1_1 gpc4295 (
      {stage3_47[12]},
      {stage4_47[4]}
   );
   gpc1_1 gpc4296 (
      {stage3_47[13]},
      {stage4_47[5]}
   );
   gpc1_1 gpc4297 (
      {stage3_47[14]},
      {stage4_47[6]}
   );
   gpc1_1 gpc4298 (
      {stage3_47[15]},
      {stage4_47[7]}
   );
   gpc1_1 gpc4299 (
      {stage3_47[16]},
      {stage4_47[8]}
   );
   gpc1_1 gpc4300 (
      {stage3_47[17]},
      {stage4_47[9]}
   );
   gpc1_1 gpc4301 (
      {stage3_47[18]},
      {stage4_47[10]}
   );
   gpc1_1 gpc4302 (
      {stage3_47[19]},
      {stage4_47[11]}
   );
   gpc1_1 gpc4303 (
      {stage3_47[20]},
      {stage4_47[12]}
   );
   gpc1_1 gpc4304 (
      {stage3_47[21]},
      {stage4_47[13]}
   );
   gpc1_1 gpc4305 (
      {stage3_47[22]},
      {stage4_47[14]}
   );
   gpc1_1 gpc4306 (
      {stage3_47[23]},
      {stage4_47[15]}
   );
   gpc1_1 gpc4307 (
      {stage3_48[8]},
      {stage4_48[4]}
   );
   gpc1_1 gpc4308 (
      {stage3_48[9]},
      {stage4_48[5]}
   );
   gpc1_1 gpc4309 (
      {stage3_48[10]},
      {stage4_48[6]}
   );
   gpc1_1 gpc4310 (
      {stage3_48[11]},
      {stage4_48[7]}
   );
   gpc1_1 gpc4311 (
      {stage3_48[12]},
      {stage4_48[8]}
   );
   gpc1_1 gpc4312 (
      {stage3_48[13]},
      {stage4_48[9]}
   );
   gpc1_1 gpc4313 (
      {stage3_48[14]},
      {stage4_48[10]}
   );
   gpc1_1 gpc4314 (
      {stage3_48[15]},
      {stage4_48[11]}
   );
   gpc1_1 gpc4315 (
      {stage3_49[6]},
      {stage4_49[5]}
   );
   gpc1_1 gpc4316 (
      {stage3_49[7]},
      {stage4_49[6]}
   );
   gpc1_1 gpc4317 (
      {stage3_49[8]},
      {stage4_49[7]}
   );
   gpc1_1 gpc4318 (
      {stage3_49[9]},
      {stage4_49[8]}
   );
   gpc1_1 gpc4319 (
      {stage3_49[10]},
      {stage4_49[9]}
   );
   gpc1_1 gpc4320 (
      {stage3_49[11]},
      {stage4_49[10]}
   );
   gpc1_1 gpc4321 (
      {stage3_49[12]},
      {stage4_49[11]}
   );
   gpc1_1 gpc4322 (
      {stage3_49[13]},
      {stage4_49[12]}
   );
   gpc1_1 gpc4323 (
      {stage3_50[31]},
      {stage4_50[6]}
   );
   gpc1_1 gpc4324 (
      {stage3_51[12]},
      {stage4_51[7]}
   );
   gpc1_1 gpc4325 (
      {stage3_51[13]},
      {stage4_51[8]}
   );
   gpc1_1 gpc4326 (
      {stage3_52[23]},
      {stage4_52[8]}
   );
   gpc1_1 gpc4327 (
      {stage3_53[7]},
      {stage4_53[6]}
   );
   gpc1_1 gpc4328 (
      {stage3_53[8]},
      {stage4_53[7]}
   );
   gpc1_1 gpc4329 (
      {stage3_53[9]},
      {stage4_53[8]}
   );
   gpc1_1 gpc4330 (
      {stage3_53[10]},
      {stage4_53[9]}
   );
   gpc1_1 gpc4331 (
      {stage3_53[11]},
      {stage4_53[10]}
   );
   gpc1_1 gpc4332 (
      {stage3_53[12]},
      {stage4_53[11]}
   );
   gpc1_1 gpc4333 (
      {stage3_53[13]},
      {stage4_53[12]}
   );
   gpc1_1 gpc4334 (
      {stage3_53[14]},
      {stage4_53[13]}
   );
   gpc1_1 gpc4335 (
      {stage3_53[15]},
      {stage4_53[14]}
   );
   gpc1_1 gpc4336 (
      {stage3_54[12]},
      {stage4_54[6]}
   );
   gpc1_1 gpc4337 (
      {stage3_54[13]},
      {stage4_54[7]}
   );
   gpc1_1 gpc4338 (
      {stage3_54[14]},
      {stage4_54[8]}
   );
   gpc1_1 gpc4339 (
      {stage3_54[15]},
      {stage4_54[9]}
   );
   gpc1_1 gpc4340 (
      {stage3_55[5]},
      {stage4_55[4]}
   );
   gpc1_1 gpc4341 (
      {stage3_55[6]},
      {stage4_55[5]}
   );
   gpc1_1 gpc4342 (
      {stage3_55[7]},
      {stage4_55[6]}
   );
   gpc1_1 gpc4343 (
      {stage3_55[8]},
      {stage4_55[7]}
   );
   gpc1_1 gpc4344 (
      {stage3_55[9]},
      {stage4_55[8]}
   );
   gpc1_1 gpc4345 (
      {stage3_55[10]},
      {stage4_55[9]}
   );
   gpc1_1 gpc4346 (
      {stage3_55[11]},
      {stage4_55[10]}
   );
   gpc1_1 gpc4347 (
      {stage3_55[12]},
      {stage4_55[11]}
   );
   gpc1_1 gpc4348 (
      {stage3_55[13]},
      {stage4_55[12]}
   );
   gpc1_1 gpc4349 (
      {stage3_55[14]},
      {stage4_55[13]}
   );
   gpc1_1 gpc4350 (
      {stage3_55[15]},
      {stage4_55[14]}
   );
   gpc1_1 gpc4351 (
      {stage3_55[16]},
      {stage4_55[15]}
   );
   gpc1_1 gpc4352 (
      {stage3_55[17]},
      {stage4_55[16]}
   );
   gpc1_1 gpc4353 (
      {stage3_56[24]},
      {stage4_56[6]}
   );
   gpc1_1 gpc4354 (
      {stage3_56[25]},
      {stage4_56[7]}
   );
   gpc1_1 gpc4355 (
      {stage3_56[26]},
      {stage4_56[8]}
   );
   gpc1_1 gpc4356 (
      {stage3_56[27]},
      {stage4_56[9]}
   );
   gpc1_1 gpc4357 (
      {stage3_56[28]},
      {stage4_56[10]}
   );
   gpc1_1 gpc4358 (
      {stage3_56[29]},
      {stage4_56[11]}
   );
   gpc1_1 gpc4359 (
      {stage3_56[30]},
      {stage4_56[12]}
   );
   gpc1_1 gpc4360 (
      {stage3_58[18]},
      {stage4_58[6]}
   );
   gpc1_1 gpc4361 (
      {stage3_58[19]},
      {stage4_58[7]}
   );
   gpc1_1 gpc4362 (
      {stage3_58[20]},
      {stage4_58[8]}
   );
   gpc1_1 gpc4363 (
      {stage3_58[21]},
      {stage4_58[9]}
   );
   gpc1_1 gpc4364 (
      {stage3_58[22]},
      {stage4_58[10]}
   );
   gpc1_1 gpc4365 (
      {stage3_58[23]},
      {stage4_58[11]}
   );
   gpc1_1 gpc4366 (
      {stage3_58[24]},
      {stage4_58[12]}
   );
   gpc1_1 gpc4367 (
      {stage3_58[25]},
      {stage4_58[13]}
   );
   gpc1_1 gpc4368 (
      {stage3_58[26]},
      {stage4_58[14]}
   );
   gpc1_1 gpc4369 (
      {stage3_58[27]},
      {stage4_58[15]}
   );
   gpc1_1 gpc4370 (
      {stage3_58[28]},
      {stage4_58[16]}
   );
   gpc1_1 gpc4371 (
      {stage3_58[29]},
      {stage4_58[17]}
   );
   gpc1_1 gpc4372 (
      {stage3_58[30]},
      {stage4_58[18]}
   );
   gpc1_1 gpc4373 (
      {stage3_58[31]},
      {stage4_58[19]}
   );
   gpc1_1 gpc4374 (
      {stage3_58[32]},
      {stage4_58[20]}
   );
   gpc1_1 gpc4375 (
      {stage3_59[18]},
      {stage4_59[7]}
   );
   gpc1_1 gpc4376 (
      {stage3_59[19]},
      {stage4_59[8]}
   );
   gpc1_1 gpc4377 (
      {stage3_59[20]},
      {stage4_59[9]}
   );
   gpc1_1 gpc4378 (
      {stage3_59[21]},
      {stage4_59[10]}
   );
   gpc1_1 gpc4379 (
      {stage3_59[22]},
      {stage4_59[11]}
   );
   gpc1_1 gpc4380 (
      {stage3_59[23]},
      {stage4_59[12]}
   );
   gpc1_1 gpc4381 (
      {stage3_59[24]},
      {stage4_59[13]}
   );
   gpc1_1 gpc4382 (
      {stage3_59[25]},
      {stage4_59[14]}
   );
   gpc1_1 gpc4383 (
      {stage3_59[26]},
      {stage4_59[15]}
   );
   gpc1_1 gpc4384 (
      {stage3_59[27]},
      {stage4_59[16]}
   );
   gpc1_1 gpc4385 (
      {stage3_60[6]},
      {stage4_60[7]}
   );
   gpc1_1 gpc4386 (
      {stage3_60[7]},
      {stage4_60[8]}
   );
   gpc1_1 gpc4387 (
      {stage3_60[8]},
      {stage4_60[9]}
   );
   gpc1_1 gpc4388 (
      {stage3_60[9]},
      {stage4_60[10]}
   );
   gpc1_1 gpc4389 (
      {stage3_60[10]},
      {stage4_60[11]}
   );
   gpc1_1 gpc4390 (
      {stage3_60[11]},
      {stage4_60[12]}
   );
   gpc1_1 gpc4391 (
      {stage3_60[12]},
      {stage4_60[13]}
   );
   gpc1_1 gpc4392 (
      {stage3_60[13]},
      {stage4_60[14]}
   );
   gpc1_1 gpc4393 (
      {stage3_60[14]},
      {stage4_60[15]}
   );
   gpc1_1 gpc4394 (
      {stage3_61[12]},
      {stage4_61[4]}
   );
   gpc1_1 gpc4395 (
      {stage3_61[13]},
      {stage4_61[5]}
   );
   gpc1_1 gpc4396 (
      {stage3_61[14]},
      {stage4_61[6]}
   );
   gpc1_1 gpc4397 (
      {stage3_61[15]},
      {stage4_61[7]}
   );
   gpc1_1 gpc4398 (
      {stage3_61[16]},
      {stage4_61[8]}
   );
   gpc1_1 gpc4399 (
      {stage3_61[17]},
      {stage4_61[9]}
   );
   gpc1_1 gpc4400 (
      {stage3_61[18]},
      {stage4_61[10]}
   );
   gpc1_1 gpc4401 (
      {stage3_61[19]},
      {stage4_61[11]}
   );
   gpc1_1 gpc4402 (
      {stage3_61[20]},
      {stage4_61[12]}
   );
   gpc1_1 gpc4403 (
      {stage3_61[21]},
      {stage4_61[13]}
   );
   gpc1_1 gpc4404 (
      {stage3_61[22]},
      {stage4_61[14]}
   );
   gpc1_1 gpc4405 (
      {stage3_61[23]},
      {stage4_61[15]}
   );
   gpc1_1 gpc4406 (
      {stage3_61[24]},
      {stage4_61[16]}
   );
   gpc1_1 gpc4407 (
      {stage3_62[18]},
      {stage4_62[5]}
   );
   gpc1_1 gpc4408 (
      {stage3_62[19]},
      {stage4_62[6]}
   );
   gpc1_1 gpc4409 (
      {stage3_62[20]},
      {stage4_62[7]}
   );
   gpc1_1 gpc4410 (
      {stage3_63[12]},
      {stage4_63[7]}
   );
   gpc1_1 gpc4411 (
      {stage3_63[13]},
      {stage4_63[8]}
   );
   gpc1_1 gpc4412 (
      {stage3_63[14]},
      {stage4_63[9]}
   );
   gpc1_1 gpc4413 (
      {stage3_63[15]},
      {stage4_63[10]}
   );
   gpc1_1 gpc4414 (
      {stage3_63[16]},
      {stage4_63[11]}
   );
   gpc1_1 gpc4415 (
      {stage3_63[17]},
      {stage4_63[12]}
   );
   gpc1_1 gpc4416 (
      {stage3_64[12]},
      {stage4_64[5]}
   );
   gpc1_1 gpc4417 (
      {stage3_64[13]},
      {stage4_64[6]}
   );
   gpc1_1 gpc4418 (
      {stage3_64[14]},
      {stage4_64[7]}
   );
   gpc1_1 gpc4419 (
      {stage3_64[15]},
      {stage4_64[8]}
   );
   gpc1_1 gpc4420 (
      {stage3_64[16]},
      {stage4_64[9]}
   );
   gpc1_1 gpc4421 (
      {stage3_64[17]},
      {stage4_64[10]}
   );
   gpc1_1 gpc4422 (
      {stage3_64[18]},
      {stage4_64[11]}
   );
   gpc1_1 gpc4423 (
      {stage3_64[19]},
      {stage4_64[12]}
   );
   gpc1_1 gpc4424 (
      {stage3_64[20]},
      {stage4_64[13]}
   );
   gpc1_1 gpc4425 (
      {stage3_64[21]},
      {stage4_64[14]}
   );
   gpc1_1 gpc4426 (
      {stage3_64[22]},
      {stage4_64[15]}
   );
   gpc1_1 gpc4427 (
      {stage3_64[23]},
      {stage4_64[16]}
   );
   gpc1_1 gpc4428 (
      {stage3_64[24]},
      {stage4_64[17]}
   );
   gpc1_1 gpc4429 (
      {stage3_64[25]},
      {stage4_64[18]}
   );
   gpc1_1 gpc4430 (
      {stage3_64[26]},
      {stage4_64[19]}
   );
   gpc1_1 gpc4431 (
      {stage3_64[27]},
      {stage4_64[20]}
   );
   gpc1_1 gpc4432 (
      {stage3_64[28]},
      {stage4_64[21]}
   );
   gpc1_1 gpc4433 (
      {stage3_65[12]},
      {stage4_65[4]}
   );
   gpc1_1 gpc4434 (
      {stage3_65[13]},
      {stage4_65[5]}
   );
   gpc1_1 gpc4435 (
      {stage3_66[0]},
      {stage4_66[4]}
   );
   gpc1_1 gpc4436 (
      {stage3_66[1]},
      {stage4_66[5]}
   );
   gpc1_1 gpc4437 (
      {stage3_66[2]},
      {stage4_66[6]}
   );
   gpc1_1 gpc4438 (
      {stage3_66[3]},
      {stage4_66[7]}
   );
   gpc1_1 gpc4439 (
      {stage3_66[4]},
      {stage4_66[8]}
   );
   gpc1_1 gpc4440 (
      {stage3_66[5]},
      {stage4_66[9]}
   );
   gpc1_1 gpc4441 (
      {stage3_66[6]},
      {stage4_66[10]}
   );
   gpc1_1 gpc4442 (
      {stage3_66[7]},
      {stage4_66[11]}
   );
   gpc1_1 gpc4443 (
      {stage3_66[8]},
      {stage4_66[12]}
   );
   gpc1_1 gpc4444 (
      {stage3_67[0]},
      {stage4_67[2]}
   );
   gpc1_1 gpc4445 (
      {stage3_67[1]},
      {stage4_67[3]}
   );
   gpc1_1 gpc4446 (
      {stage3_67[2]},
      {stage4_67[4]}
   );
   gpc1_1 gpc4447 (
      {stage3_67[3]},
      {stage4_67[5]}
   );
   gpc1_1 gpc4448 (
      {stage3_67[4]},
      {stage4_67[6]}
   );
   gpc1_1 gpc4449 (
      {stage3_68[0]},
      {stage4_68[0]}
   );
   gpc1_1 gpc4450 (
      {stage3_68[1]},
      {stage4_68[1]}
   );
   gpc1343_5 gpc4451 (
      {stage4_0[0], stage4_0[1], stage4_0[2]},
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3]},
      {stage4_2[0], stage4_2[1], stage4_2[2]},
      {stage4_3[0]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc606_5 gpc4452 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[1]}
   );
   gpc606_5 gpc4453 (
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[1],stage5_5[1]}
   );
   gpc615_5 gpc4454 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[0]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[2]}
   );
   gpc606_5 gpc4455 (
      {stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[1],stage5_11[1],stage5_10[1],stage5_9[2]}
   );
   gpc606_5 gpc4456 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[1]}
   );
   gpc615_5 gpc4457 (
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4]},
      {stage4_15[6]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[1],stage5_16[1],stage5_15[1],stage5_14[1]}
   );
   gpc615_5 gpc4458 (
      {stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage4_16[6]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[1],stage5_17[2],stage5_16[2],stage5_15[2]}
   );
   gpc606_5 gpc4459 (
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[0],stage5_19[1],stage5_18[2],stage5_17[3]}
   );
   gpc606_5 gpc4460 (
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], 1'b0},
      {stage4_19[6], stage4_19[7], stage4_19[8], stage4_19[9], stage4_19[10], stage4_19[11]},
      {stage5_21[1],stage5_20[1],stage5_19[2],stage5_18[3],stage5_17[4]}
   );
   gpc615_5 gpc4461 (
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4]},
      {stage4_19[12]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[2],stage5_20[2],stage5_19[3],stage5_18[4]}
   );
   gpc606_5 gpc4462 (
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], 1'b0},
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage5_24[0],stage5_23[0],stage5_22[1],stage5_21[3],stage5_20[3]}
   );
   gpc7_3 gpc4463 (
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5], stage4_21[6]},
      {stage5_23[1],stage5_22[2],stage5_21[4]}
   );
   gpc606_5 gpc4464 (
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[0],stage5_25[0],stage5_24[1],stage5_23[2]}
   );
   gpc1406_5 gpc4465 (
      {stage4_24[0], stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5]},
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3]},
      {stage4_27[0]},
      {stage5_28[0],stage5_27[1],stage5_26[1],stage5_25[1],stage5_24[2]}
   );
   gpc1406_5 gpc4466 (
      {stage4_24[6], stage4_24[7], stage4_24[8], stage4_24[9], stage4_24[10], stage4_24[11]},
      {stage4_26[4], stage4_26[5], stage4_26[6], stage4_26[7]},
      {stage4_27[1]},
      {stage5_28[1],stage5_27[2],stage5_26[2],stage5_25[2],stage5_24[3]}
   );
   gpc615_5 gpc4467 (
      {stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5], stage4_27[6]},
      {stage4_28[0]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[0],stage5_29[0],stage5_28[2],stage5_27[3]}
   );
   gpc2135_5 gpc4468 (
      {stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage4_29[6], stage4_29[7], stage4_29[8]},
      {stage4_30[0]},
      {stage4_31[0], stage4_31[1]},
      {stage5_32[0],stage5_31[1],stage5_30[1],stage5_29[1],stage5_28[3]}
   );
   gpc606_5 gpc4469 (
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9], stage4_28[10], stage4_28[11]},
      {stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5], stage4_30[6]},
      {stage5_32[1],stage5_31[2],stage5_30[2],stage5_29[2],stage5_28[4]}
   );
   gpc615_5 gpc4470 (
      {stage4_30[7], stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11]},
      {stage4_31[2]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[0],stage5_32[2],stage5_31[3],stage5_30[3]}
   );
   gpc615_5 gpc4471 (
      {stage4_30[12], stage4_30[13], stage4_30[14], stage4_30[15], 1'b0},
      {stage4_31[3]},
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11]},
      {stage5_34[1],stage5_33[1],stage5_32[3],stage5_31[4],stage5_30[4]}
   );
   gpc615_5 gpc4472 (
      {stage4_31[4], stage4_31[5], stage4_31[6], stage4_31[7], stage4_31[8]},
      {stage4_32[12]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[2],stage5_33[2],stage5_32[4],stage5_31[5]}
   );
   gpc1343_5 gpc4473 (
      {stage4_33[6], stage4_33[7], stage4_33[8]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3]},
      {stage4_35[0], stage4_35[1], stage4_35[2]},
      {stage4_36[0]},
      {stage5_37[0],stage5_36[0],stage5_35[1],stage5_34[3],stage5_33[3]}
   );
   gpc1343_5 gpc4474 (
      {stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage4_34[4], stage4_34[5], stage4_34[6], stage4_34[7]},
      {stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage4_36[1]},
      {stage5_37[1],stage5_36[1],stage5_35[2],stage5_34[4],stage5_33[4]}
   );
   gpc615_5 gpc4475 (
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10]},
      {stage4_36[2]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage5_39[0],stage5_38[0],stage5_37[2],stage5_36[2],stage5_35[3]}
   );
   gpc606_5 gpc4476 (
      {stage4_36[3], stage4_36[4], stage4_36[5], stage4_36[6], stage4_36[7], stage4_36[8]},
      {stage4_38[0], stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4], stage4_38[5]},
      {stage5_40[0],stage5_39[1],stage5_38[1],stage5_37[3],stage5_36[3]}
   );
   gpc207_4 gpc4477 (
      {stage4_39[0], stage4_39[1], stage4_39[2], stage4_39[3], stage4_39[4], stage4_39[5], stage4_39[6]},
      {stage4_41[0], stage4_41[1]},
      {stage5_42[0],stage5_41[0],stage5_40[1],stage5_39[2]}
   );
   gpc606_5 gpc4478 (
      {stage4_40[0], stage4_40[1], stage4_40[2], stage4_40[3], stage4_40[4], stage4_40[5]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[0],stage5_42[1],stage5_41[1],stage5_40[2]}
   );
   gpc606_5 gpc4479 (
      {stage4_40[6], stage4_40[7], stage4_40[8], stage4_40[9], stage4_40[10], stage4_40[11]},
      {stage4_42[6], stage4_42[7], stage4_42[8], stage4_42[9], stage4_42[10], stage4_42[11]},
      {stage5_44[1],stage5_43[1],stage5_42[2],stage5_41[2],stage5_40[3]}
   );
   gpc606_5 gpc4480 (
      {stage4_41[2], stage4_41[3], stage4_41[4], stage4_41[5], stage4_41[6], stage4_41[7]},
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], stage4_43[5]},
      {stage5_45[0],stage5_44[2],stage5_43[2],stage5_42[3],stage5_41[3]}
   );
   gpc615_5 gpc4481 (
      {stage4_42[12], stage4_42[13], stage4_42[14], stage4_42[15], stage4_42[16]},
      {stage4_43[6]},
      {stage4_44[0], stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage5_46[0],stage5_45[1],stage5_44[3],stage5_43[3],stage5_42[4]}
   );
   gpc606_5 gpc4482 (
      {stage4_44[6], stage4_44[7], stage4_44[8], stage4_44[9], stage4_44[10], stage4_44[11]},
      {stage4_46[0], stage4_46[1], stage4_46[2], stage4_46[3], stage4_46[4], stage4_46[5]},
      {stage5_48[0],stage5_47[0],stage5_46[1],stage5_45[2],stage5_44[4]}
   );
   gpc23_3 gpc4483 (
      {stage4_45[0], stage4_45[1], stage4_45[2]},
      {stage4_46[6], stage4_46[7]},
      {stage5_47[1],stage5_46[2],stage5_45[3]}
   );
   gpc606_5 gpc4484 (
      {stage4_45[3], stage4_45[4], stage4_45[5], stage4_45[6], stage4_45[7], stage4_45[8]},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4], stage4_47[5]},
      {stage5_49[0],stage5_48[1],stage5_47[2],stage5_46[3],stage5_45[4]}
   );
   gpc615_5 gpc4485 (
      {stage4_46[8], stage4_46[9], stage4_46[10], stage4_46[11], stage4_46[12]},
      {stage4_47[6]},
      {stage4_48[0], stage4_48[1], stage4_48[2], stage4_48[3], stage4_48[4], stage4_48[5]},
      {stage5_50[0],stage5_49[1],stage5_48[2],stage5_47[3],stage5_46[4]}
   );
   gpc615_5 gpc4486 (
      {stage4_46[13], stage4_46[14], stage4_46[15], stage4_46[16], stage4_46[17]},
      {stage4_47[7]},
      {stage4_48[6], stage4_48[7], stage4_48[8], stage4_48[9], stage4_48[10], stage4_48[11]},
      {stage5_50[1],stage5_49[2],stage5_48[3],stage5_47[4],stage5_46[5]}
   );
   gpc135_4 gpc4487 (
      {stage4_49[0], stage4_49[1], stage4_49[2], stage4_49[3], stage4_49[4]},
      {stage4_50[0], stage4_50[1], stage4_50[2]},
      {stage4_51[0]},
      {stage5_52[0],stage5_51[0],stage5_50[2],stage5_49[3]}
   );
   gpc606_5 gpc4488 (
      {stage4_49[5], stage4_49[6], stage4_49[7], stage4_49[8], stage4_49[9], stage4_49[10]},
      {stage4_51[1], stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5], stage4_51[6]},
      {stage5_53[0],stage5_52[1],stage5_51[1],stage5_50[3],stage5_49[4]}
   );
   gpc615_5 gpc4489 (
      {stage4_50[3], stage4_50[4], stage4_50[5], stage4_50[6], 1'b0},
      {stage4_51[7]},
      {stage4_52[0], stage4_52[1], stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5]},
      {stage5_54[0],stage5_53[1],stage5_52[2],stage5_51[2],stage5_50[4]}
   );
   gpc606_5 gpc4490 (
      {stage4_53[0], stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5]},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5]},
      {stage5_57[0],stage5_56[0],stage5_55[0],stage5_54[1],stage5_53[2]}
   );
   gpc606_5 gpc4491 (
      {stage4_53[6], stage4_53[7], stage4_53[8], stage4_53[9], stage4_53[10], stage4_53[11]},
      {stage4_55[6], stage4_55[7], stage4_55[8], stage4_55[9], stage4_55[10], stage4_55[11]},
      {stage5_57[1],stage5_56[1],stage5_55[1],stage5_54[2],stage5_53[3]}
   );
   gpc615_5 gpc4492 (
      {stage4_54[0], stage4_54[1], stage4_54[2], stage4_54[3], stage4_54[4]},
      {stage4_55[12]},
      {stage4_56[0], stage4_56[1], stage4_56[2], stage4_56[3], stage4_56[4], stage4_56[5]},
      {stage5_58[0],stage5_57[2],stage5_56[2],stage5_55[2],stage5_54[3]}
   );
   gpc606_5 gpc4493 (
      {stage4_56[6], stage4_56[7], stage4_56[8], stage4_56[9], stage4_56[10], stage4_56[11]},
      {stage4_58[0], stage4_58[1], stage4_58[2], stage4_58[3], stage4_58[4], stage4_58[5]},
      {stage5_60[0],stage5_59[0],stage5_58[1],stage5_57[3],stage5_56[3]}
   );
   gpc1343_5 gpc4494 (
      {stage4_57[0], stage4_57[1], stage4_57[2]},
      {stage4_58[6], stage4_58[7], stage4_58[8], stage4_58[9]},
      {stage4_59[0], stage4_59[1], stage4_59[2]},
      {stage4_60[0]},
      {stage5_61[0],stage5_60[1],stage5_59[1],stage5_58[2],stage5_57[4]}
   );
   gpc1343_5 gpc4495 (
      {stage4_57[3], stage4_57[4], stage4_57[5]},
      {stage4_58[10], stage4_58[11], stage4_58[12], stage4_58[13]},
      {stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage4_60[1]},
      {stage5_61[1],stage5_60[2],stage5_59[2],stage5_58[3],stage5_57[5]}
   );
   gpc606_5 gpc4496 (
      {stage4_58[14], stage4_58[15], stage4_58[16], stage4_58[17], stage4_58[18], stage4_58[19]},
      {stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5], stage4_60[6], stage4_60[7]},
      {stage5_62[0],stage5_61[2],stage5_60[3],stage5_59[3],stage5_58[4]}
   );
   gpc606_5 gpc4497 (
      {stage4_59[6], stage4_59[7], stage4_59[8], stage4_59[9], stage4_59[10], stage4_59[11]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[1],stage5_61[3],stage5_60[4],stage5_59[4]}
   );
   gpc606_5 gpc4498 (
      {stage4_59[12], stage4_59[13], stage4_59[14], stage4_59[15], stage4_59[16], 1'b0},
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], stage4_61[10], stage4_61[11]},
      {stage5_63[1],stage5_62[2],stage5_61[4],stage5_60[5],stage5_59[5]}
   );
   gpc606_5 gpc4499 (
      {stage4_60[8], stage4_60[9], stage4_60[10], stage4_60[11], stage4_60[12], stage4_60[13]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[2],stage5_62[3],stage5_61[5],stage5_60[6]}
   );
   gpc135_4 gpc4500 (
      {stage4_63[0], stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4]},
      {stage4_64[0], stage4_64[1], stage4_64[2]},
      {stage4_65[0]},
      {stage5_66[0],stage5_65[0],stage5_64[1],stage5_63[3]}
   );
   gpc606_5 gpc4501 (
      {stage4_64[3], stage4_64[4], stage4_64[5], stage4_64[6], stage4_64[7], stage4_64[8]},
      {stage4_66[0], stage4_66[1], stage4_66[2], stage4_66[3], stage4_66[4], stage4_66[5]},
      {stage5_68[0],stage5_67[0],stage5_66[1],stage5_65[1],stage5_64[2]}
   );
   gpc606_5 gpc4502 (
      {stage4_64[9], stage4_64[10], stage4_64[11], stage4_64[12], stage4_64[13], stage4_64[14]},
      {stage4_66[6], stage4_66[7], stage4_66[8], stage4_66[9], stage4_66[10], stage4_66[11]},
      {stage5_68[1],stage5_67[1],stage5_66[2],stage5_65[2],stage5_64[3]}
   );
   gpc606_5 gpc4503 (
      {stage4_65[1], stage4_65[2], stage4_65[3], stage4_65[4], stage4_65[5], 1'b0},
      {stage4_67[0], stage4_67[1], stage4_67[2], stage4_67[3], stage4_67[4], stage4_67[5]},
      {stage5_69[0],stage5_68[2],stage5_67[2],stage5_66[3],stage5_65[3]}
   );
   gpc1_1 gpc4504 (
      {stage4_0[3]},
      {stage5_0[1]}
   );
   gpc1_1 gpc4505 (
      {stage4_2[3]},
      {stage5_2[1]}
   );
   gpc1_1 gpc4506 (
      {stage4_2[4]},
      {stage5_2[2]}
   );
   gpc1_1 gpc4507 (
      {stage4_2[5]},
      {stage5_2[3]}
   );
   gpc1_1 gpc4508 (
      {stage4_2[6]},
      {stage5_2[4]}
   );
   gpc1_1 gpc4509 (
      {stage4_3[1]},
      {stage5_3[1]}
   );
   gpc1_1 gpc4510 (
      {stage4_3[2]},
      {stage5_3[2]}
   );
   gpc1_1 gpc4511 (
      {stage4_3[3]},
      {stage5_3[3]}
   );
   gpc1_1 gpc4512 (
      {stage4_3[4]},
      {stage5_3[4]}
   );
   gpc1_1 gpc4513 (
      {stage4_4[6]},
      {stage5_4[2]}
   );
   gpc1_1 gpc4514 (
      {stage4_4[7]},
      {stage5_4[3]}
   );
   gpc1_1 gpc4515 (
      {stage4_4[8]},
      {stage5_4[4]}
   );
   gpc1_1 gpc4516 (
      {stage4_5[6]},
      {stage5_5[2]}
   );
   gpc1_1 gpc4517 (
      {stage4_5[7]},
      {stage5_5[3]}
   );
   gpc1_1 gpc4518 (
      {stage4_5[8]},
      {stage5_5[4]}
   );
   gpc1_1 gpc4519 (
      {stage4_6[6]},
      {stage5_6[2]}
   );
   gpc1_1 gpc4520 (
      {stage4_6[7]},
      {stage5_6[3]}
   );
   gpc1_1 gpc4521 (
      {stage4_6[8]},
      {stage5_6[4]}
   );
   gpc1_1 gpc4522 (
      {stage4_6[9]},
      {stage5_6[5]}
   );
   gpc1_1 gpc4523 (
      {stage4_6[10]},
      {stage5_6[6]}
   );
   gpc1_1 gpc4524 (
      {stage4_6[11]},
      {stage5_6[7]}
   );
   gpc1_1 gpc4525 (
      {stage4_6[12]},
      {stage5_6[8]}
   );
   gpc1_1 gpc4526 (
      {stage4_6[13]},
      {stage5_6[9]}
   );
   gpc1_1 gpc4527 (
      {stage4_7[6]},
      {stage5_7[2]}
   );
   gpc1_1 gpc4528 (
      {stage4_7[7]},
      {stage5_7[3]}
   );
   gpc1_1 gpc4529 (
      {stage4_8[5]},
      {stage5_8[3]}
   );
   gpc1_1 gpc4530 (
      {stage4_8[6]},
      {stage5_8[4]}
   );
   gpc1_1 gpc4531 (
      {stage4_8[7]},
      {stage5_8[5]}
   );
   gpc1_1 gpc4532 (
      {stage4_8[8]},
      {stage5_8[6]}
   );
   gpc1_1 gpc4533 (
      {stage4_8[9]},
      {stage5_8[7]}
   );
   gpc1_1 gpc4534 (
      {stage4_10[6]},
      {stage5_10[2]}
   );
   gpc1_1 gpc4535 (
      {stage4_10[7]},
      {stage5_10[3]}
   );
   gpc1_1 gpc4536 (
      {stage4_10[8]},
      {stage5_10[4]}
   );
   gpc1_1 gpc4537 (
      {stage4_11[6]},
      {stage5_11[2]}
   );
   gpc1_1 gpc4538 (
      {stage4_12[0]},
      {stage5_12[2]}
   );
   gpc1_1 gpc4539 (
      {stage4_12[1]},
      {stage5_12[3]}
   );
   gpc1_1 gpc4540 (
      {stage4_12[2]},
      {stage5_12[4]}
   );
   gpc1_1 gpc4541 (
      {stage4_12[3]},
      {stage5_12[5]}
   );
   gpc1_1 gpc4542 (
      {stage4_12[4]},
      {stage5_12[6]}
   );
   gpc1_1 gpc4543 (
      {stage4_12[5]},
      {stage5_12[7]}
   );
   gpc1_1 gpc4544 (
      {stage4_12[6]},
      {stage5_12[8]}
   );
   gpc1_1 gpc4545 (
      {stage4_12[7]},
      {stage5_12[9]}
   );
   gpc1_1 gpc4546 (
      {stage4_12[8]},
      {stage5_12[10]}
   );
   gpc1_1 gpc4547 (
      {stage4_13[6]},
      {stage5_13[2]}
   );
   gpc1_1 gpc4548 (
      {stage4_13[7]},
      {stage5_13[3]}
   );
   gpc1_1 gpc4549 (
      {stage4_13[8]},
      {stage5_13[4]}
   );
   gpc1_1 gpc4550 (
      {stage4_13[9]},
      {stage5_13[5]}
   );
   gpc1_1 gpc4551 (
      {stage4_14[5]},
      {stage5_14[2]}
   );
   gpc1_1 gpc4552 (
      {stage4_14[6]},
      {stage5_14[3]}
   );
   gpc1_1 gpc4553 (
      {stage4_14[7]},
      {stage5_14[4]}
   );
   gpc1_1 gpc4554 (
      {stage4_14[8]},
      {stage5_14[5]}
   );
   gpc1_1 gpc4555 (
      {stage4_14[9]},
      {stage5_14[6]}
   );
   gpc1_1 gpc4556 (
      {stage4_14[10]},
      {stage5_14[7]}
   );
   gpc1_1 gpc4557 (
      {stage4_15[12]},
      {stage5_15[3]}
   );
   gpc1_1 gpc4558 (
      {stage4_15[13]},
      {stage5_15[4]}
   );
   gpc1_1 gpc4559 (
      {stage4_15[14]},
      {stage5_15[5]}
   );
   gpc1_1 gpc4560 (
      {stage4_15[15]},
      {stage5_15[6]}
   );
   gpc1_1 gpc4561 (
      {stage4_15[16]},
      {stage5_15[7]}
   );
   gpc1_1 gpc4562 (
      {stage4_16[7]},
      {stage5_16[3]}
   );
   gpc1_1 gpc4563 (
      {stage4_16[8]},
      {stage5_16[4]}
   );
   gpc1_1 gpc4564 (
      {stage4_16[9]},
      {stage5_16[5]}
   );
   gpc1_1 gpc4565 (
      {stage4_16[10]},
      {stage5_16[6]}
   );
   gpc1_1 gpc4566 (
      {stage4_16[11]},
      {stage5_16[7]}
   );
   gpc1_1 gpc4567 (
      {stage4_16[12]},
      {stage5_16[8]}
   );
   gpc1_1 gpc4568 (
      {stage4_18[5]},
      {stage5_18[5]}
   );
   gpc1_1 gpc4569 (
      {stage4_19[13]},
      {stage5_19[4]}
   );
   gpc1_1 gpc4570 (
      {stage4_19[14]},
      {stage5_19[5]}
   );
   gpc1_1 gpc4571 (
      {stage4_19[15]},
      {stage5_19[6]}
   );
   gpc1_1 gpc4572 (
      {stage4_21[7]},
      {stage5_21[5]}
   );
   gpc1_1 gpc4573 (
      {stage4_22[6]},
      {stage5_22[3]}
   );
   gpc1_1 gpc4574 (
      {stage4_22[7]},
      {stage5_22[4]}
   );
   gpc1_1 gpc4575 (
      {stage4_22[8]},
      {stage5_22[5]}
   );
   gpc1_1 gpc4576 (
      {stage4_22[9]},
      {stage5_22[6]}
   );
   gpc1_1 gpc4577 (
      {stage4_22[10]},
      {stage5_22[7]}
   );
   gpc1_1 gpc4578 (
      {stage4_22[11]},
      {stage5_22[8]}
   );
   gpc1_1 gpc4579 (
      {stage4_22[12]},
      {stage5_22[9]}
   );
   gpc1_1 gpc4580 (
      {stage4_22[13]},
      {stage5_22[10]}
   );
   gpc1_1 gpc4581 (
      {stage4_23[6]},
      {stage5_23[3]}
   );
   gpc1_1 gpc4582 (
      {stage4_23[7]},
      {stage5_23[4]}
   );
   gpc1_1 gpc4583 (
      {stage4_23[8]},
      {stage5_23[5]}
   );
   gpc1_1 gpc4584 (
      {stage4_23[9]},
      {stage5_23[6]}
   );
   gpc1_1 gpc4585 (
      {stage4_24[12]},
      {stage5_24[4]}
   );
   gpc1_1 gpc4586 (
      {stage4_24[13]},
      {stage5_24[5]}
   );
   gpc1_1 gpc4587 (
      {stage4_24[14]},
      {stage5_24[6]}
   );
   gpc1_1 gpc4588 (
      {stage4_24[15]},
      {stage5_24[7]}
   );
   gpc1_1 gpc4589 (
      {stage4_24[16]},
      {stage5_24[8]}
   );
   gpc1_1 gpc4590 (
      {stage4_24[17]},
      {stage5_24[9]}
   );
   gpc1_1 gpc4591 (
      {stage4_29[9]},
      {stage5_29[3]}
   );
   gpc1_1 gpc4592 (
      {stage4_32[13]},
      {stage5_32[5]}
   );
   gpc1_1 gpc4593 (
      {stage4_32[14]},
      {stage5_32[6]}
   );
   gpc1_1 gpc4594 (
      {stage4_32[15]},
      {stage5_32[7]}
   );
   gpc1_1 gpc4595 (
      {stage4_32[16]},
      {stage5_32[8]}
   );
   gpc1_1 gpc4596 (
      {stage4_32[17]},
      {stage5_32[9]}
   );
   gpc1_1 gpc4597 (
      {stage4_32[18]},
      {stage5_32[10]}
   );
   gpc1_1 gpc4598 (
      {stage4_32[19]},
      {stage5_32[11]}
   );
   gpc1_1 gpc4599 (
      {stage4_34[8]},
      {stage5_34[5]}
   );
   gpc1_1 gpc4600 (
      {stage4_34[9]},
      {stage5_34[6]}
   );
   gpc1_1 gpc4601 (
      {stage4_34[10]},
      {stage5_34[7]}
   );
   gpc1_1 gpc4602 (
      {stage4_36[9]},
      {stage5_36[4]}
   );
   gpc1_1 gpc4603 (
      {stage4_39[7]},
      {stage5_39[3]}
   );
   gpc1_1 gpc4604 (
      {stage4_39[8]},
      {stage5_39[4]}
   );
   gpc1_1 gpc4605 (
      {stage4_39[9]},
      {stage5_39[5]}
   );
   gpc1_1 gpc4606 (
      {stage4_40[12]},
      {stage5_40[4]}
   );
   gpc1_1 gpc4607 (
      {stage4_40[13]},
      {stage5_40[5]}
   );
   gpc1_1 gpc4608 (
      {stage4_41[8]},
      {stage5_41[4]}
   );
   gpc1_1 gpc4609 (
      {stage4_41[9]},
      {stage5_41[5]}
   );
   gpc1_1 gpc4610 (
      {stage4_41[10]},
      {stage5_41[6]}
   );
   gpc1_1 gpc4611 (
      {stage4_41[11]},
      {stage5_41[7]}
   );
   gpc1_1 gpc4612 (
      {stage4_41[12]},
      {stage5_41[8]}
   );
   gpc1_1 gpc4613 (
      {stage4_41[13]},
      {stage5_41[9]}
   );
   gpc1_1 gpc4614 (
      {stage4_41[14]},
      {stage5_41[10]}
   );
   gpc1_1 gpc4615 (
      {stage4_41[15]},
      {stage5_41[11]}
   );
   gpc1_1 gpc4616 (
      {stage4_41[16]},
      {stage5_41[12]}
   );
   gpc1_1 gpc4617 (
      {stage4_44[12]},
      {stage5_44[5]}
   );
   gpc1_1 gpc4618 (
      {stage4_47[8]},
      {stage5_47[5]}
   );
   gpc1_1 gpc4619 (
      {stage4_47[9]},
      {stage5_47[6]}
   );
   gpc1_1 gpc4620 (
      {stage4_47[10]},
      {stage5_47[7]}
   );
   gpc1_1 gpc4621 (
      {stage4_47[11]},
      {stage5_47[8]}
   );
   gpc1_1 gpc4622 (
      {stage4_47[12]},
      {stage5_47[9]}
   );
   gpc1_1 gpc4623 (
      {stage4_47[13]},
      {stage5_47[10]}
   );
   gpc1_1 gpc4624 (
      {stage4_47[14]},
      {stage5_47[11]}
   );
   gpc1_1 gpc4625 (
      {stage4_47[15]},
      {stage5_47[12]}
   );
   gpc1_1 gpc4626 (
      {stage4_49[11]},
      {stage5_49[5]}
   );
   gpc1_1 gpc4627 (
      {stage4_49[12]},
      {stage5_49[6]}
   );
   gpc1_1 gpc4628 (
      {stage4_51[8]},
      {stage5_51[3]}
   );
   gpc1_1 gpc4629 (
      {stage4_52[6]},
      {stage5_52[3]}
   );
   gpc1_1 gpc4630 (
      {stage4_52[7]},
      {stage5_52[4]}
   );
   gpc1_1 gpc4631 (
      {stage4_52[8]},
      {stage5_52[5]}
   );
   gpc1_1 gpc4632 (
      {stage4_53[12]},
      {stage5_53[4]}
   );
   gpc1_1 gpc4633 (
      {stage4_53[13]},
      {stage5_53[5]}
   );
   gpc1_1 gpc4634 (
      {stage4_53[14]},
      {stage5_53[6]}
   );
   gpc1_1 gpc4635 (
      {stage4_54[5]},
      {stage5_54[4]}
   );
   gpc1_1 gpc4636 (
      {stage4_54[6]},
      {stage5_54[5]}
   );
   gpc1_1 gpc4637 (
      {stage4_54[7]},
      {stage5_54[6]}
   );
   gpc1_1 gpc4638 (
      {stage4_54[8]},
      {stage5_54[7]}
   );
   gpc1_1 gpc4639 (
      {stage4_54[9]},
      {stage5_54[8]}
   );
   gpc1_1 gpc4640 (
      {stage4_55[13]},
      {stage5_55[3]}
   );
   gpc1_1 gpc4641 (
      {stage4_55[14]},
      {stage5_55[4]}
   );
   gpc1_1 gpc4642 (
      {stage4_55[15]},
      {stage5_55[5]}
   );
   gpc1_1 gpc4643 (
      {stage4_55[16]},
      {stage5_55[6]}
   );
   gpc1_1 gpc4644 (
      {stage4_56[12]},
      {stage5_56[4]}
   );
   gpc1_1 gpc4645 (
      {stage4_58[20]},
      {stage5_58[5]}
   );
   gpc1_1 gpc4646 (
      {stage4_60[14]},
      {stage5_60[7]}
   );
   gpc1_1 gpc4647 (
      {stage4_60[15]},
      {stage5_60[8]}
   );
   gpc1_1 gpc4648 (
      {stage4_61[12]},
      {stage5_61[6]}
   );
   gpc1_1 gpc4649 (
      {stage4_61[13]},
      {stage5_61[7]}
   );
   gpc1_1 gpc4650 (
      {stage4_61[14]},
      {stage5_61[8]}
   );
   gpc1_1 gpc4651 (
      {stage4_61[15]},
      {stage5_61[9]}
   );
   gpc1_1 gpc4652 (
      {stage4_61[16]},
      {stage5_61[10]}
   );
   gpc1_1 gpc4653 (
      {stage4_62[6]},
      {stage5_62[4]}
   );
   gpc1_1 gpc4654 (
      {stage4_62[7]},
      {stage5_62[5]}
   );
   gpc1_1 gpc4655 (
      {stage4_63[5]},
      {stage5_63[4]}
   );
   gpc1_1 gpc4656 (
      {stage4_63[6]},
      {stage5_63[5]}
   );
   gpc1_1 gpc4657 (
      {stage4_63[7]},
      {stage5_63[6]}
   );
   gpc1_1 gpc4658 (
      {stage4_63[8]},
      {stage5_63[7]}
   );
   gpc1_1 gpc4659 (
      {stage4_63[9]},
      {stage5_63[8]}
   );
   gpc1_1 gpc4660 (
      {stage4_63[10]},
      {stage5_63[9]}
   );
   gpc1_1 gpc4661 (
      {stage4_63[11]},
      {stage5_63[10]}
   );
   gpc1_1 gpc4662 (
      {stage4_63[12]},
      {stage5_63[11]}
   );
   gpc1_1 gpc4663 (
      {stage4_64[15]},
      {stage5_64[4]}
   );
   gpc1_1 gpc4664 (
      {stage4_64[16]},
      {stage5_64[5]}
   );
   gpc1_1 gpc4665 (
      {stage4_64[17]},
      {stage5_64[6]}
   );
   gpc1_1 gpc4666 (
      {stage4_64[18]},
      {stage5_64[7]}
   );
   gpc1_1 gpc4667 (
      {stage4_64[19]},
      {stage5_64[8]}
   );
   gpc1_1 gpc4668 (
      {stage4_64[20]},
      {stage5_64[9]}
   );
   gpc1_1 gpc4669 (
      {stage4_64[21]},
      {stage5_64[10]}
   );
   gpc1_1 gpc4670 (
      {stage4_66[12]},
      {stage5_66[4]}
   );
   gpc1_1 gpc4671 (
      {stage4_67[6]},
      {stage5_67[3]}
   );
   gpc1_1 gpc4672 (
      {stage4_68[0]},
      {stage5_68[3]}
   );
   gpc1_1 gpc4673 (
      {stage4_68[1]},
      {stage5_68[4]}
   );
   gpc615_5 gpc4674 (
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], 1'b0},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc1415_5 gpc4675 (
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4]},
      {stage5_7[0]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3]},
      {stage5_9[0]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1]}
   );
   gpc1415_5 gpc4676 (
      {stage5_6[5], stage5_6[6], stage5_6[7], stage5_6[8], stage5_6[9]},
      {stage5_7[1]},
      {stage5_8[4], stage5_8[5], stage5_8[6], stage5_8[7]},
      {stage5_9[1]},
      {stage6_10[1],stage6_9[1],stage6_8[1],stage6_7[2],stage6_6[2]}
   );
   gpc606_5 gpc4677 (
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage6_16[0],stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[0]}
   );
   gpc606_5 gpc4678 (
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[1],stage6_13[1]}
   );
   gpc606_5 gpc4679 (
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5]},
      {stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[1],stage6_16[2]}
   );
   gpc2135_5 gpc4680 (
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4]},
      {stage5_20[0], stage5_20[1], stage5_20[2]},
      {stage5_21[0]},
      {stage5_22[0], stage5_22[1]},
      {stage6_23[0],stage6_22[0],stage6_21[0],stage6_20[1],stage6_19[1]}
   );
   gpc1163_5 gpc4681 (
      {stage5_22[2], stage5_22[3], stage5_22[4]},
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3], stage5_23[4], stage5_23[5]},
      {stage5_24[0]},
      {stage5_25[0]},
      {stage6_26[0],stage6_25[0],stage6_24[0],stage6_23[1],stage6_22[1]}
   );
   gpc615_5 gpc4682 (
      {stage5_22[5], stage5_22[6], stage5_22[7], stage5_22[8], stage5_22[9]},
      {stage5_23[6]},
      {stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], stage5_24[6]},
      {stage6_26[1],stage6_25[1],stage6_24[1],stage6_23[2],stage6_22[2]}
   );
   gpc1343_5 gpc4683 (
      {stage5_24[7], stage5_24[8], stage5_24[9]},
      {stage5_25[1], stage5_25[2], 1'b0, 1'b0},
      {stage5_26[0], stage5_26[1], stage5_26[2]},
      {stage5_27[0]},
      {stage6_28[0],stage6_27[0],stage6_26[2],stage6_25[2],stage6_24[2]}
   );
   gpc3_2 gpc4684 (
      {stage5_27[1], stage5_27[2], stage5_27[3]},
      {stage6_28[1],stage6_27[1]}
   );
   gpc606_5 gpc4685 (
      {stage5_28[0], stage5_28[1], stage5_28[2], stage5_28[3], stage5_28[4], 1'b0},
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], 1'b0},
      {stage6_32[0],stage6_31[0],stage6_30[0],stage6_29[0],stage6_28[2]}
   );
   gpc606_5 gpc4686 (
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], 1'b0, 1'b0},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[1],stage6_31[1],stage6_30[1],stage6_29[1]}
   );
   gpc606_5 gpc4687 (
      {stage5_32[0], stage5_32[1], stage5_32[2], stage5_32[3], stage5_32[4], stage5_32[5]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5]},
      {stage6_36[0],stage6_35[0],stage6_34[0],stage6_33[1],stage6_32[2]}
   );
   gpc615_5 gpc4688 (
      {stage5_33[0], stage5_33[1], stage5_33[2], stage5_33[3], stage5_33[4]},
      {stage5_34[6]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3], 1'b0, 1'b0},
      {stage6_37[0],stage6_36[1],stage6_35[1],stage6_34[1],stage6_33[2]}
   );
   gpc615_5 gpc4689 (
      {stage5_38[0], stage5_38[1], 1'b0, 1'b0, 1'b0},
      {stage5_39[0]},
      {stage5_40[0], stage5_40[1], stage5_40[2], stage5_40[3], stage5_40[4], stage5_40[5]},
      {stage6_42[0],stage6_41[0],stage6_40[0],stage6_39[0],stage6_38[0]}
   );
   gpc606_5 gpc4690 (
      {stage5_39[1], stage5_39[2], stage5_39[3], stage5_39[4], stage5_39[5], 1'b0},
      {stage5_41[0], stage5_41[1], stage5_41[2], stage5_41[3], stage5_41[4], stage5_41[5]},
      {stage6_43[0],stage6_42[1],stage6_41[1],stage6_40[1],stage6_39[1]}
   );
   gpc606_5 gpc4691 (
      {stage5_41[6], stage5_41[7], stage5_41[8], stage5_41[9], stage5_41[10], stage5_41[11]},
      {stage5_43[0], stage5_43[1], stage5_43[2], stage5_43[3], 1'b0, 1'b0},
      {stage6_45[0],stage6_44[0],stage6_43[1],stage6_42[2],stage6_41[2]}
   );
   gpc606_5 gpc4692 (
      {stage5_44[0], stage5_44[1], stage5_44[2], stage5_44[3], stage5_44[4], stage5_44[5]},
      {stage5_46[0], stage5_46[1], stage5_46[2], stage5_46[3], stage5_46[4], stage5_46[5]},
      {stage6_48[0],stage6_47[0],stage6_46[0],stage6_45[1],stage6_44[1]}
   );
   gpc606_5 gpc4693 (
      {stage5_45[0], stage5_45[1], stage5_45[2], stage5_45[3], stage5_45[4], 1'b0},
      {stage5_47[0], stage5_47[1], stage5_47[2], stage5_47[3], stage5_47[4], stage5_47[5]},
      {stage6_49[0],stage6_48[1],stage6_47[1],stage6_46[1],stage6_45[2]}
   );
   gpc615_5 gpc4694 (
      {stage5_47[6], stage5_47[7], stage5_47[8], stage5_47[9], stage5_47[10]},
      {stage5_48[0]},
      {stage5_49[0], stage5_49[1], stage5_49[2], stage5_49[3], stage5_49[4], stage5_49[5]},
      {stage6_51[0],stage6_50[0],stage6_49[1],stage6_48[2],stage6_47[2]}
   );
   gpc1343_5 gpc4695 (
      {stage5_50[0], stage5_50[1], stage5_50[2]},
      {stage5_51[0], stage5_51[1], stage5_51[2], stage5_51[3]},
      {stage5_52[0], stage5_52[1], stage5_52[2]},
      {stage5_53[0]},
      {stage6_54[0],stage6_53[0],stage6_52[0],stage6_51[1],stage6_50[1]}
   );
   gpc223_4 gpc4696 (
      {stage5_53[1], stage5_53[2], stage5_53[3]},
      {stage5_54[0], stage5_54[1]},
      {stage5_55[0], stage5_55[1]},
      {stage6_56[0],stage6_55[0],stage6_54[1],stage6_53[1]}
   );
   gpc207_4 gpc4697 (
      {stage5_54[2], stage5_54[3], stage5_54[4], stage5_54[5], stage5_54[6], stage5_54[7], stage5_54[8]},
      {stage5_56[0], stage5_56[1]},
      {stage6_57[0],stage6_56[1],stage6_55[1],stage6_54[2]}
   );
   gpc615_5 gpc4698 (
      {stage5_55[2], stage5_55[3], stage5_55[4], stage5_55[5], stage5_55[6]},
      {stage5_56[2]},
      {stage5_57[0], stage5_57[1], stage5_57[2], stage5_57[3], stage5_57[4], stage5_57[5]},
      {stage6_59[0],stage6_58[0],stage6_57[1],stage6_56[2],stage6_55[2]}
   );
   gpc606_5 gpc4699 (
      {stage5_58[0], stage5_58[1], stage5_58[2], stage5_58[3], stage5_58[4], stage5_58[5]},
      {stage5_60[0], stage5_60[1], stage5_60[2], stage5_60[3], stage5_60[4], stage5_60[5]},
      {stage6_62[0],stage6_61[0],stage6_60[0],stage6_59[1],stage6_58[1]}
   );
   gpc606_5 gpc4700 (
      {stage5_59[0], stage5_59[1], stage5_59[2], stage5_59[3], stage5_59[4], stage5_59[5]},
      {stage5_61[0], stage5_61[1], stage5_61[2], stage5_61[3], stage5_61[4], stage5_61[5]},
      {stage6_63[0],stage6_62[1],stage6_61[1],stage6_60[1],stage6_59[2]}
   );
   gpc606_5 gpc4701 (
      {stage5_61[6], stage5_61[7], stage5_61[8], stage5_61[9], stage5_61[10], 1'b0},
      {stage5_63[0], stage5_63[1], stage5_63[2], stage5_63[3], stage5_63[4], stage5_63[5]},
      {stage6_65[0],stage6_64[0],stage6_63[1],stage6_62[2],stage6_61[2]}
   );
   gpc606_5 gpc4702 (
      {stage5_62[0], stage5_62[1], stage5_62[2], stage5_62[3], stage5_62[4], stage5_62[5]},
      {stage5_64[0], stage5_64[1], stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5]},
      {stage6_66[0],stage6_65[1],stage6_64[1],stage6_63[2],stage6_62[3]}
   );
   gpc606_5 gpc4703 (
      {stage5_63[6], stage5_63[7], stage5_63[8], stage5_63[9], stage5_63[10], stage5_63[11]},
      {stage5_65[0], stage5_65[1], stage5_65[2], stage5_65[3], 1'b0, 1'b0},
      {stage6_67[0],stage6_66[1],stage6_65[2],stage6_64[2],stage6_63[3]}
   );
   gpc606_5 gpc4704 (
      {stage5_64[6], stage5_64[7], stage5_64[8], stage5_64[9], stage5_64[10], 1'b0},
      {stage5_66[0], stage5_66[1], stage5_66[2], stage5_66[3], stage5_66[4], 1'b0},
      {stage6_68[0],stage6_67[1],stage6_66[2],stage6_65[3],stage6_64[3]}
   );
   gpc1_1 gpc4705 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc4706 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc4707 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc4708 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc4709 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc4710 (
      {stage5_2[2]},
      {stage6_2[2]}
   );
   gpc1_1 gpc4711 (
      {stage5_2[3]},
      {stage6_2[3]}
   );
   gpc1_1 gpc4712 (
      {stage5_2[4]},
      {stage6_2[4]}
   );
   gpc1_1 gpc4713 (
      {stage5_4[1]},
      {stage6_4[1]}
   );
   gpc1_1 gpc4714 (
      {stage5_4[2]},
      {stage6_4[2]}
   );
   gpc1_1 gpc4715 (
      {stage5_4[3]},
      {stage6_4[3]}
   );
   gpc1_1 gpc4716 (
      {stage5_4[4]},
      {stage6_4[4]}
   );
   gpc1_1 gpc4717 (
      {stage5_7[2]},
      {stage6_7[3]}
   );
   gpc1_1 gpc4718 (
      {stage5_7[3]},
      {stage6_7[4]}
   );
   gpc1_1 gpc4719 (
      {stage5_9[2]},
      {stage6_9[2]}
   );
   gpc1_1 gpc4720 (
      {stage5_10[0]},
      {stage6_10[2]}
   );
   gpc1_1 gpc4721 (
      {stage5_10[1]},
      {stage6_10[3]}
   );
   gpc1_1 gpc4722 (
      {stage5_10[2]},
      {stage6_10[4]}
   );
   gpc1_1 gpc4723 (
      {stage5_10[3]},
      {stage6_10[5]}
   );
   gpc1_1 gpc4724 (
      {stage5_10[4]},
      {stage6_10[6]}
   );
   gpc1_1 gpc4725 (
      {stage5_11[0]},
      {stage6_11[0]}
   );
   gpc1_1 gpc4726 (
      {stage5_11[1]},
      {stage6_11[1]}
   );
   gpc1_1 gpc4727 (
      {stage5_11[2]},
      {stage6_11[2]}
   );
   gpc1_1 gpc4728 (
      {stage5_12[6]},
      {stage6_12[1]}
   );
   gpc1_1 gpc4729 (
      {stage5_12[7]},
      {stage6_12[2]}
   );
   gpc1_1 gpc4730 (
      {stage5_12[8]},
      {stage6_12[3]}
   );
   gpc1_1 gpc4731 (
      {stage5_12[9]},
      {stage6_12[4]}
   );
   gpc1_1 gpc4732 (
      {stage5_12[10]},
      {stage6_12[5]}
   );
   gpc1_1 gpc4733 (
      {stage5_14[6]},
      {stage6_14[2]}
   );
   gpc1_1 gpc4734 (
      {stage5_14[7]},
      {stage6_14[3]}
   );
   gpc1_1 gpc4735 (
      {stage5_15[6]},
      {stage6_15[2]}
   );
   gpc1_1 gpc4736 (
      {stage5_15[7]},
      {stage6_15[3]}
   );
   gpc1_1 gpc4737 (
      {stage5_16[6]},
      {stage6_16[3]}
   );
   gpc1_1 gpc4738 (
      {stage5_16[7]},
      {stage6_16[4]}
   );
   gpc1_1 gpc4739 (
      {stage5_16[8]},
      {stage6_16[5]}
   );
   gpc1_1 gpc4740 (
      {stage5_17[0]},
      {stage6_17[2]}
   );
   gpc1_1 gpc4741 (
      {stage5_17[1]},
      {stage6_17[3]}
   );
   gpc1_1 gpc4742 (
      {stage5_17[2]},
      {stage6_17[4]}
   );
   gpc1_1 gpc4743 (
      {stage5_17[3]},
      {stage6_17[5]}
   );
   gpc1_1 gpc4744 (
      {stage5_17[4]},
      {stage6_17[6]}
   );
   gpc1_1 gpc4745 (
      {stage5_19[5]},
      {stage6_19[2]}
   );
   gpc1_1 gpc4746 (
      {stage5_19[6]},
      {stage6_19[3]}
   );
   gpc1_1 gpc4747 (
      {stage5_20[3]},
      {stage6_20[2]}
   );
   gpc1_1 gpc4748 (
      {stage5_21[1]},
      {stage6_21[1]}
   );
   gpc1_1 gpc4749 (
      {stage5_21[2]},
      {stage6_21[2]}
   );
   gpc1_1 gpc4750 (
      {stage5_21[3]},
      {stage6_21[3]}
   );
   gpc1_1 gpc4751 (
      {stage5_21[4]},
      {stage6_21[4]}
   );
   gpc1_1 gpc4752 (
      {stage5_21[5]},
      {stage6_21[5]}
   );
   gpc1_1 gpc4753 (
      {stage5_22[10]},
      {stage6_22[3]}
   );
   gpc1_1 gpc4754 (
      {stage5_32[6]},
      {stage6_32[3]}
   );
   gpc1_1 gpc4755 (
      {stage5_32[7]},
      {stage6_32[4]}
   );
   gpc1_1 gpc4756 (
      {stage5_32[8]},
      {stage6_32[5]}
   );
   gpc1_1 gpc4757 (
      {stage5_32[9]},
      {stage6_32[6]}
   );
   gpc1_1 gpc4758 (
      {stage5_32[10]},
      {stage6_32[7]}
   );
   gpc1_1 gpc4759 (
      {stage5_32[11]},
      {stage6_32[8]}
   );
   gpc1_1 gpc4760 (
      {stage5_34[7]},
      {stage6_34[2]}
   );
   gpc1_1 gpc4761 (
      {stage5_36[0]},
      {stage6_36[2]}
   );
   gpc1_1 gpc4762 (
      {stage5_36[1]},
      {stage6_36[3]}
   );
   gpc1_1 gpc4763 (
      {stage5_36[2]},
      {stage6_36[4]}
   );
   gpc1_1 gpc4764 (
      {stage5_36[3]},
      {stage6_36[5]}
   );
   gpc1_1 gpc4765 (
      {stage5_36[4]},
      {stage6_36[6]}
   );
   gpc1_1 gpc4766 (
      {stage5_37[0]},
      {stage6_37[1]}
   );
   gpc1_1 gpc4767 (
      {stage5_37[1]},
      {stage6_37[2]}
   );
   gpc1_1 gpc4768 (
      {stage5_37[2]},
      {stage6_37[3]}
   );
   gpc1_1 gpc4769 (
      {stage5_37[3]},
      {stage6_37[4]}
   );
   gpc1_1 gpc4770 (
      {stage5_41[12]},
      {stage6_41[3]}
   );
   gpc1_1 gpc4771 (
      {stage5_42[0]},
      {stage6_42[3]}
   );
   gpc1_1 gpc4772 (
      {stage5_42[1]},
      {stage6_42[4]}
   );
   gpc1_1 gpc4773 (
      {stage5_42[2]},
      {stage6_42[5]}
   );
   gpc1_1 gpc4774 (
      {stage5_42[3]},
      {stage6_42[6]}
   );
   gpc1_1 gpc4775 (
      {stage5_42[4]},
      {stage6_42[7]}
   );
   gpc1_1 gpc4776 (
      {stage5_47[11]},
      {stage6_47[3]}
   );
   gpc1_1 gpc4777 (
      {stage5_47[12]},
      {stage6_47[4]}
   );
   gpc1_1 gpc4778 (
      {stage5_48[1]},
      {stage6_48[3]}
   );
   gpc1_1 gpc4779 (
      {stage5_48[2]},
      {stage6_48[4]}
   );
   gpc1_1 gpc4780 (
      {stage5_48[3]},
      {stage6_48[5]}
   );
   gpc1_1 gpc4781 (
      {stage5_49[6]},
      {stage6_49[2]}
   );
   gpc1_1 gpc4782 (
      {stage5_50[3]},
      {stage6_50[2]}
   );
   gpc1_1 gpc4783 (
      {stage5_50[4]},
      {stage6_50[3]}
   );
   gpc1_1 gpc4784 (
      {stage5_52[3]},
      {stage6_52[1]}
   );
   gpc1_1 gpc4785 (
      {stage5_52[4]},
      {stage6_52[2]}
   );
   gpc1_1 gpc4786 (
      {stage5_52[5]},
      {stage6_52[3]}
   );
   gpc1_1 gpc4787 (
      {stage5_53[4]},
      {stage6_53[2]}
   );
   gpc1_1 gpc4788 (
      {stage5_53[5]},
      {stage6_53[3]}
   );
   gpc1_1 gpc4789 (
      {stage5_53[6]},
      {stage6_53[4]}
   );
   gpc1_1 gpc4790 (
      {stage5_56[3]},
      {stage6_56[3]}
   );
   gpc1_1 gpc4791 (
      {stage5_56[4]},
      {stage6_56[4]}
   );
   gpc1_1 gpc4792 (
      {stage5_60[6]},
      {stage6_60[2]}
   );
   gpc1_1 gpc4793 (
      {stage5_60[7]},
      {stage6_60[3]}
   );
   gpc1_1 gpc4794 (
      {stage5_60[8]},
      {stage6_60[4]}
   );
   gpc1_1 gpc4795 (
      {stage5_67[0]},
      {stage6_67[2]}
   );
   gpc1_1 gpc4796 (
      {stage5_67[1]},
      {stage6_67[3]}
   );
   gpc1_1 gpc4797 (
      {stage5_67[2]},
      {stage6_67[4]}
   );
   gpc1_1 gpc4798 (
      {stage5_67[3]},
      {stage6_67[5]}
   );
   gpc1_1 gpc4799 (
      {stage5_68[0]},
      {stage6_68[1]}
   );
   gpc1_1 gpc4800 (
      {stage5_68[1]},
      {stage6_68[2]}
   );
   gpc1_1 gpc4801 (
      {stage5_68[2]},
      {stage6_68[3]}
   );
   gpc1_1 gpc4802 (
      {stage5_68[3]},
      {stage6_68[4]}
   );
   gpc1_1 gpc4803 (
      {stage5_68[4]},
      {stage6_68[5]}
   );
   gpc1_1 gpc4804 (
      {stage5_69[0]},
      {stage6_69[0]}
   );
   gpc1415_5 gpc4805 (
      {stage6_2[0], stage6_2[1], stage6_2[2], stage6_2[3], stage6_2[4]},
      {stage6_3[0]},
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3]},
      {stage6_5[0]},
      {stage7_6[0],stage7_5[0],stage7_4[0],stage7_3[0],stage7_2[0]}
   );
   gpc23_3 gpc4806 (
      {stage6_6[0], stage6_6[1], stage6_6[2]},
      {stage6_7[0], stage6_7[1]},
      {stage7_8[0],stage7_7[0],stage7_6[1]}
   );
   gpc223_4 gpc4807 (
      {stage6_7[2], stage6_7[3], stage6_7[4]},
      {stage6_8[0], stage6_8[1]},
      {stage6_9[0], stage6_9[1]},
      {stage7_10[0],stage7_9[0],stage7_8[1],stage7_7[1]}
   );
   gpc207_4 gpc4808 (
      {stage6_10[0], stage6_10[1], stage6_10[2], stage6_10[3], stage6_10[4], stage6_10[5], stage6_10[6]},
      {stage6_12[0], stage6_12[1]},
      {stage7_13[0],stage7_12[0],stage7_11[0],stage7_10[1]}
   );
   gpc1343_5 gpc4809 (
      {stage6_11[0], stage6_11[1], stage6_11[2]},
      {stage6_12[2], stage6_12[3], stage6_12[4], stage6_12[5]},
      {stage6_13[0], stage6_13[1], 1'b0},
      {stage6_14[0]},
      {stage7_15[0],stage7_14[0],stage7_13[1],stage7_12[1],stage7_11[1]}
   );
   gpc1343_5 gpc4810 (
      {stage6_14[1], stage6_14[2], stage6_14[3]},
      {stage6_15[0], stage6_15[1], stage6_15[2], stage6_15[3]},
      {stage6_16[0], stage6_16[1], stage6_16[2]},
      {stage6_17[0]},
      {stage7_18[0],stage7_17[0],stage7_16[0],stage7_15[1],stage7_14[1]}
   );
   gpc1163_5 gpc4811 (
      {stage6_16[3], stage6_16[4], stage6_16[5]},
      {stage6_17[1], stage6_17[2], stage6_17[3], stage6_17[4], stage6_17[5], stage6_17[6]},
      {stage6_18[0]},
      {stage6_19[0]},
      {stage7_20[0],stage7_19[0],stage7_18[1],stage7_17[1],stage7_16[1]}
   );
   gpc1343_5 gpc4812 (
      {stage6_19[1], stage6_19[2], stage6_19[3]},
      {stage6_20[0], stage6_20[1], stage6_20[2], 1'b0},
      {stage6_21[0], stage6_21[1], stage6_21[2]},
      {stage6_22[0]},
      {stage7_23[0],stage7_22[0],stage7_21[0],stage7_20[1],stage7_19[1]}
   );
   gpc1343_5 gpc4813 (
      {stage6_21[3], stage6_21[4], stage6_21[5]},
      {stage6_22[1], stage6_22[2], stage6_22[3], 1'b0},
      {stage6_23[0], stage6_23[1], stage6_23[2]},
      {stage6_24[0]},
      {stage7_25[0],stage7_24[0],stage7_23[1],stage7_22[1],stage7_21[1]}
   );
   gpc1343_5 gpc4814 (
      {stage6_24[1], stage6_24[2], 1'b0},
      {stage6_25[0], stage6_25[1], stage6_25[2], 1'b0},
      {stage6_26[0], stage6_26[1], stage6_26[2]},
      {stage6_27[0]},
      {stage7_28[0],stage7_27[0],stage7_26[0],stage7_25[1],stage7_24[1]}
   );
   gpc15_3 gpc4815 (
      {stage6_28[0], stage6_28[1], stage6_28[2], 1'b0, 1'b0},
      {stage6_29[0]},
      {stage7_30[0],stage7_29[0],stage7_28[1]}
   );
   gpc615_5 gpc4816 (
      {stage6_30[0], stage6_30[1], 1'b0, 1'b0, 1'b0},
      {stage6_31[0]},
      {stage6_32[0], stage6_32[1], stage6_32[2], stage6_32[3], stage6_32[4], stage6_32[5]},
      {stage7_34[0],stage7_33[0],stage7_32[0],stage7_31[0],stage7_30[1]}
   );
   gpc1343_5 gpc4817 (
      {stage6_32[6], stage6_32[7], stage6_32[8]},
      {stage6_33[0], stage6_33[1], stage6_33[2], 1'b0},
      {stage6_34[0], stage6_34[1], stage6_34[2]},
      {stage6_35[0]},
      {stage7_36[0],stage7_35[0],stage7_34[1],stage7_33[1],stage7_32[1]}
   );
   gpc7_3 gpc4818 (
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3], stage6_36[4], stage6_36[5], stage6_36[6]},
      {stage7_38[0],stage7_37[0],stage7_36[1]}
   );
   gpc2135_5 gpc4819 (
      {stage6_37[0], stage6_37[1], stage6_37[2], stage6_37[3], stage6_37[4]},
      {stage6_38[0], 1'b0, 1'b0},
      {stage6_39[0]},
      {stage6_40[0], stage6_40[1]},
      {stage7_41[0],stage7_40[0],stage7_39[0],stage7_38[1],stage7_37[1]}
   );
   gpc135_4 gpc4820 (
      {stage6_41[0], stage6_41[1], stage6_41[2], stage6_41[3], 1'b0},
      {stage6_42[0], stage6_42[1], stage6_42[2]},
      {stage6_43[0]},
      {stage7_44[0],stage7_43[0],stage7_42[0],stage7_41[1]}
   );
   gpc615_5 gpc4821 (
      {stage6_42[3], stage6_42[4], stage6_42[5], stage6_42[6], stage6_42[7]},
      {stage6_43[1]},
      {stage6_44[0], stage6_44[1], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage7_46[0],stage7_45[0],stage7_44[1],stage7_43[1],stage7_42[1]}
   );
   gpc2223_5 gpc4822 (
      {stage6_45[0], stage6_45[1], stage6_45[2]},
      {stage6_46[0], stage6_46[1]},
      {stage6_47[0], stage6_47[1]},
      {stage6_48[0], stage6_48[1]},
      {stage7_49[0],stage7_48[0],stage7_47[0],stage7_46[1],stage7_45[1]}
   );
   gpc1343_5 gpc4823 (
      {stage6_47[2], stage6_47[3], stage6_47[4]},
      {stage6_48[2], stage6_48[3], stage6_48[4], stage6_48[5]},
      {stage6_49[0], stage6_49[1], stage6_49[2]},
      {stage6_50[0]},
      {stage7_51[0],stage7_50[0],stage7_49[1],stage7_48[1],stage7_47[1]}
   );
   gpc1343_5 gpc4824 (
      {stage6_50[1], stage6_50[2], stage6_50[3]},
      {stage6_51[0], stage6_51[1], 1'b0, 1'b0},
      {stage6_52[0], stage6_52[1], stage6_52[2]},
      {stage6_53[0]},
      {stage7_54[0],stage7_53[0],stage7_52[0],stage7_51[1],stage7_50[1]}
   );
   gpc1343_5 gpc4825 (
      {stage6_52[3], 1'b0, 1'b0},
      {stage6_53[1], stage6_53[2], stage6_53[3], stage6_53[4]},
      {stage6_54[0], stage6_54[1], stage6_54[2]},
      {stage6_55[0]},
      {stage7_56[0],stage7_55[0],stage7_54[1],stage7_53[1],stage7_52[1]}
   );
   gpc1163_5 gpc4826 (
      {stage6_55[1], stage6_55[2], 1'b0},
      {stage6_56[0], stage6_56[1], stage6_56[2], stage6_56[3], stage6_56[4], 1'b0},
      {stage6_57[0]},
      {stage6_58[0]},
      {stage7_59[0],stage7_58[0],stage7_57[0],stage7_56[1],stage7_55[1]}
   );
   gpc1343_5 gpc4827 (
      {stage6_59[0], stage6_59[1], stage6_59[2]},
      {stage6_60[0], stage6_60[1], stage6_60[2], stage6_60[3]},
      {stage6_61[0], stage6_61[1], stage6_61[2]},
      {stage6_62[0]},
      {stage7_63[0],stage7_62[0],stage7_61[0],stage7_60[0],stage7_59[1]}
   );
   gpc1343_5 gpc4828 (
      {stage6_62[1], stage6_62[2], stage6_62[3]},
      {stage6_63[0], stage6_63[1], stage6_63[2], stage6_63[3]},
      {stage6_64[0], stage6_64[1], stage6_64[2]},
      {stage6_65[0]},
      {stage7_66[0],stage7_65[0],stage7_64[0],stage7_63[1],stage7_62[1]}
   );
   gpc1343_5 gpc4829 (
      {stage6_65[1], stage6_65[2], stage6_65[3]},
      {stage6_66[0], stage6_66[1], stage6_66[2], 1'b0},
      {stage6_67[0], stage6_67[1], stage6_67[2]},
      {stage6_68[0]},
      {stage7_69[0],stage7_68[0],stage7_67[0],stage7_66[1],stage7_65[1]}
   );
   gpc1163_5 gpc4830 (
      {stage6_67[3], stage6_67[4], stage6_67[5]},
      {stage6_68[1], stage6_68[2], stage6_68[3], stage6_68[4], stage6_68[5], 1'b0},
      {stage6_69[0]},
      {1'b0},
      {stage7_71[0],stage7_70[0],stage7_69[1],stage7_68[1],stage7_67[1]}
   );
   gpc1_1 gpc4831 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc4832 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc4833 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc4834 (
      {stage6_4[4]},
      {stage7_4[1]}
   );
   gpc1_1 gpc4835 (
      {stage6_9[2]},
      {stage7_9[1]}
   );
   gpc1_1 gpc4836 (
      {stage6_27[1]},
      {stage7_27[1]}
   );
   gpc1_1 gpc4837 (
      {stage6_29[1]},
      {stage7_29[1]}
   );
   gpc1_1 gpc4838 (
      {stage6_31[1]},
      {stage7_31[1]}
   );
   gpc1_1 gpc4839 (
      {stage6_35[1]},
      {stage7_35[1]}
   );
   gpc1_1 gpc4840 (
      {stage6_39[1]},
      {stage7_39[1]}
   );
   gpc1_1 gpc4841 (
      {stage6_57[1]},
      {stage7_57[1]}
   );
   gpc1_1 gpc4842 (
      {stage6_58[1]},
      {stage7_58[1]}
   );
   gpc1_1 gpc4843 (
      {stage6_60[4]},
      {stage7_60[1]}
   );
   gpc1_1 gpc4844 (
      {stage6_64[3]},
      {stage7_64[1]}
   );
endmodule

module testbench();
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    reg [161:0] src16;
    reg [161:0] src17;
    reg [161:0] src18;
    reg [161:0] src19;
    reg [161:0] src20;
    reg [161:0] src21;
    reg [161:0] src22;
    reg [161:0] src23;
    reg [161:0] src24;
    reg [161:0] src25;
    reg [161:0] src26;
    reg [161:0] src27;
    reg [161:0] src28;
    reg [161:0] src29;
    reg [161:0] src30;
    reg [161:0] src31;
    reg [161:0] src32;
    reg [161:0] src33;
    reg [161:0] src34;
    reg [161:0] src35;
    reg [161:0] src36;
    reg [161:0] src37;
    reg [161:0] src38;
    reg [161:0] src39;
    reg [161:0] src40;
    reg [161:0] src41;
    reg [161:0] src42;
    reg [161:0] src43;
    reg [161:0] src44;
    reg [161:0] src45;
    reg [161:0] src46;
    reg [161:0] src47;
    reg [161:0] src48;
    reg [161:0] src49;
    reg [161:0] src50;
    reg [161:0] src51;
    reg [161:0] src52;
    reg [161:0] src53;
    reg [161:0] src54;
    reg [161:0] src55;
    reg [161:0] src56;
    reg [161:0] src57;
    reg [161:0] src58;
    reg [161:0] src59;
    reg [161:0] src60;
    reg [161:0] src61;
    reg [161:0] src62;
    reg [161:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [0:0] dst71;
    wire [71:0] srcsum;
    wire [71:0] dstsum;
    wire test;
    compressor_CLA162_64 compressor_CLA162_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70),
        .dst71(dst71));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127] + src32[128] + src32[129] + src32[130] + src32[131] + src32[132] + src32[133] + src32[134] + src32[135] + src32[136] + src32[137] + src32[138] + src32[139] + src32[140] + src32[141] + src32[142] + src32[143] + src32[144] + src32[145] + src32[146] + src32[147] + src32[148] + src32[149] + src32[150] + src32[151] + src32[152] + src32[153] + src32[154] + src32[155] + src32[156] + src32[157] + src32[158] + src32[159] + src32[160] + src32[161])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127] + src33[128] + src33[129] + src33[130] + src33[131] + src33[132] + src33[133] + src33[134] + src33[135] + src33[136] + src33[137] + src33[138] + src33[139] + src33[140] + src33[141] + src33[142] + src33[143] + src33[144] + src33[145] + src33[146] + src33[147] + src33[148] + src33[149] + src33[150] + src33[151] + src33[152] + src33[153] + src33[154] + src33[155] + src33[156] + src33[157] + src33[158] + src33[159] + src33[160] + src33[161])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127] + src34[128] + src34[129] + src34[130] + src34[131] + src34[132] + src34[133] + src34[134] + src34[135] + src34[136] + src34[137] + src34[138] + src34[139] + src34[140] + src34[141] + src34[142] + src34[143] + src34[144] + src34[145] + src34[146] + src34[147] + src34[148] + src34[149] + src34[150] + src34[151] + src34[152] + src34[153] + src34[154] + src34[155] + src34[156] + src34[157] + src34[158] + src34[159] + src34[160] + src34[161])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127] + src35[128] + src35[129] + src35[130] + src35[131] + src35[132] + src35[133] + src35[134] + src35[135] + src35[136] + src35[137] + src35[138] + src35[139] + src35[140] + src35[141] + src35[142] + src35[143] + src35[144] + src35[145] + src35[146] + src35[147] + src35[148] + src35[149] + src35[150] + src35[151] + src35[152] + src35[153] + src35[154] + src35[155] + src35[156] + src35[157] + src35[158] + src35[159] + src35[160] + src35[161])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127] + src36[128] + src36[129] + src36[130] + src36[131] + src36[132] + src36[133] + src36[134] + src36[135] + src36[136] + src36[137] + src36[138] + src36[139] + src36[140] + src36[141] + src36[142] + src36[143] + src36[144] + src36[145] + src36[146] + src36[147] + src36[148] + src36[149] + src36[150] + src36[151] + src36[152] + src36[153] + src36[154] + src36[155] + src36[156] + src36[157] + src36[158] + src36[159] + src36[160] + src36[161])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127] + src37[128] + src37[129] + src37[130] + src37[131] + src37[132] + src37[133] + src37[134] + src37[135] + src37[136] + src37[137] + src37[138] + src37[139] + src37[140] + src37[141] + src37[142] + src37[143] + src37[144] + src37[145] + src37[146] + src37[147] + src37[148] + src37[149] + src37[150] + src37[151] + src37[152] + src37[153] + src37[154] + src37[155] + src37[156] + src37[157] + src37[158] + src37[159] + src37[160] + src37[161])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127] + src38[128] + src38[129] + src38[130] + src38[131] + src38[132] + src38[133] + src38[134] + src38[135] + src38[136] + src38[137] + src38[138] + src38[139] + src38[140] + src38[141] + src38[142] + src38[143] + src38[144] + src38[145] + src38[146] + src38[147] + src38[148] + src38[149] + src38[150] + src38[151] + src38[152] + src38[153] + src38[154] + src38[155] + src38[156] + src38[157] + src38[158] + src38[159] + src38[160] + src38[161])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127] + src39[128] + src39[129] + src39[130] + src39[131] + src39[132] + src39[133] + src39[134] + src39[135] + src39[136] + src39[137] + src39[138] + src39[139] + src39[140] + src39[141] + src39[142] + src39[143] + src39[144] + src39[145] + src39[146] + src39[147] + src39[148] + src39[149] + src39[150] + src39[151] + src39[152] + src39[153] + src39[154] + src39[155] + src39[156] + src39[157] + src39[158] + src39[159] + src39[160] + src39[161])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127] + src40[128] + src40[129] + src40[130] + src40[131] + src40[132] + src40[133] + src40[134] + src40[135] + src40[136] + src40[137] + src40[138] + src40[139] + src40[140] + src40[141] + src40[142] + src40[143] + src40[144] + src40[145] + src40[146] + src40[147] + src40[148] + src40[149] + src40[150] + src40[151] + src40[152] + src40[153] + src40[154] + src40[155] + src40[156] + src40[157] + src40[158] + src40[159] + src40[160] + src40[161])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127] + src41[128] + src41[129] + src41[130] + src41[131] + src41[132] + src41[133] + src41[134] + src41[135] + src41[136] + src41[137] + src41[138] + src41[139] + src41[140] + src41[141] + src41[142] + src41[143] + src41[144] + src41[145] + src41[146] + src41[147] + src41[148] + src41[149] + src41[150] + src41[151] + src41[152] + src41[153] + src41[154] + src41[155] + src41[156] + src41[157] + src41[158] + src41[159] + src41[160] + src41[161])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127] + src42[128] + src42[129] + src42[130] + src42[131] + src42[132] + src42[133] + src42[134] + src42[135] + src42[136] + src42[137] + src42[138] + src42[139] + src42[140] + src42[141] + src42[142] + src42[143] + src42[144] + src42[145] + src42[146] + src42[147] + src42[148] + src42[149] + src42[150] + src42[151] + src42[152] + src42[153] + src42[154] + src42[155] + src42[156] + src42[157] + src42[158] + src42[159] + src42[160] + src42[161])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127] + src43[128] + src43[129] + src43[130] + src43[131] + src43[132] + src43[133] + src43[134] + src43[135] + src43[136] + src43[137] + src43[138] + src43[139] + src43[140] + src43[141] + src43[142] + src43[143] + src43[144] + src43[145] + src43[146] + src43[147] + src43[148] + src43[149] + src43[150] + src43[151] + src43[152] + src43[153] + src43[154] + src43[155] + src43[156] + src43[157] + src43[158] + src43[159] + src43[160] + src43[161])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127] + src44[128] + src44[129] + src44[130] + src44[131] + src44[132] + src44[133] + src44[134] + src44[135] + src44[136] + src44[137] + src44[138] + src44[139] + src44[140] + src44[141] + src44[142] + src44[143] + src44[144] + src44[145] + src44[146] + src44[147] + src44[148] + src44[149] + src44[150] + src44[151] + src44[152] + src44[153] + src44[154] + src44[155] + src44[156] + src44[157] + src44[158] + src44[159] + src44[160] + src44[161])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127] + src45[128] + src45[129] + src45[130] + src45[131] + src45[132] + src45[133] + src45[134] + src45[135] + src45[136] + src45[137] + src45[138] + src45[139] + src45[140] + src45[141] + src45[142] + src45[143] + src45[144] + src45[145] + src45[146] + src45[147] + src45[148] + src45[149] + src45[150] + src45[151] + src45[152] + src45[153] + src45[154] + src45[155] + src45[156] + src45[157] + src45[158] + src45[159] + src45[160] + src45[161])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127] + src46[128] + src46[129] + src46[130] + src46[131] + src46[132] + src46[133] + src46[134] + src46[135] + src46[136] + src46[137] + src46[138] + src46[139] + src46[140] + src46[141] + src46[142] + src46[143] + src46[144] + src46[145] + src46[146] + src46[147] + src46[148] + src46[149] + src46[150] + src46[151] + src46[152] + src46[153] + src46[154] + src46[155] + src46[156] + src46[157] + src46[158] + src46[159] + src46[160] + src46[161])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127] + src47[128] + src47[129] + src47[130] + src47[131] + src47[132] + src47[133] + src47[134] + src47[135] + src47[136] + src47[137] + src47[138] + src47[139] + src47[140] + src47[141] + src47[142] + src47[143] + src47[144] + src47[145] + src47[146] + src47[147] + src47[148] + src47[149] + src47[150] + src47[151] + src47[152] + src47[153] + src47[154] + src47[155] + src47[156] + src47[157] + src47[158] + src47[159] + src47[160] + src47[161])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127] + src48[128] + src48[129] + src48[130] + src48[131] + src48[132] + src48[133] + src48[134] + src48[135] + src48[136] + src48[137] + src48[138] + src48[139] + src48[140] + src48[141] + src48[142] + src48[143] + src48[144] + src48[145] + src48[146] + src48[147] + src48[148] + src48[149] + src48[150] + src48[151] + src48[152] + src48[153] + src48[154] + src48[155] + src48[156] + src48[157] + src48[158] + src48[159] + src48[160] + src48[161])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127] + src49[128] + src49[129] + src49[130] + src49[131] + src49[132] + src49[133] + src49[134] + src49[135] + src49[136] + src49[137] + src49[138] + src49[139] + src49[140] + src49[141] + src49[142] + src49[143] + src49[144] + src49[145] + src49[146] + src49[147] + src49[148] + src49[149] + src49[150] + src49[151] + src49[152] + src49[153] + src49[154] + src49[155] + src49[156] + src49[157] + src49[158] + src49[159] + src49[160] + src49[161])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127] + src50[128] + src50[129] + src50[130] + src50[131] + src50[132] + src50[133] + src50[134] + src50[135] + src50[136] + src50[137] + src50[138] + src50[139] + src50[140] + src50[141] + src50[142] + src50[143] + src50[144] + src50[145] + src50[146] + src50[147] + src50[148] + src50[149] + src50[150] + src50[151] + src50[152] + src50[153] + src50[154] + src50[155] + src50[156] + src50[157] + src50[158] + src50[159] + src50[160] + src50[161])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127] + src51[128] + src51[129] + src51[130] + src51[131] + src51[132] + src51[133] + src51[134] + src51[135] + src51[136] + src51[137] + src51[138] + src51[139] + src51[140] + src51[141] + src51[142] + src51[143] + src51[144] + src51[145] + src51[146] + src51[147] + src51[148] + src51[149] + src51[150] + src51[151] + src51[152] + src51[153] + src51[154] + src51[155] + src51[156] + src51[157] + src51[158] + src51[159] + src51[160] + src51[161])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127] + src52[128] + src52[129] + src52[130] + src52[131] + src52[132] + src52[133] + src52[134] + src52[135] + src52[136] + src52[137] + src52[138] + src52[139] + src52[140] + src52[141] + src52[142] + src52[143] + src52[144] + src52[145] + src52[146] + src52[147] + src52[148] + src52[149] + src52[150] + src52[151] + src52[152] + src52[153] + src52[154] + src52[155] + src52[156] + src52[157] + src52[158] + src52[159] + src52[160] + src52[161])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127] + src53[128] + src53[129] + src53[130] + src53[131] + src53[132] + src53[133] + src53[134] + src53[135] + src53[136] + src53[137] + src53[138] + src53[139] + src53[140] + src53[141] + src53[142] + src53[143] + src53[144] + src53[145] + src53[146] + src53[147] + src53[148] + src53[149] + src53[150] + src53[151] + src53[152] + src53[153] + src53[154] + src53[155] + src53[156] + src53[157] + src53[158] + src53[159] + src53[160] + src53[161])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127] + src54[128] + src54[129] + src54[130] + src54[131] + src54[132] + src54[133] + src54[134] + src54[135] + src54[136] + src54[137] + src54[138] + src54[139] + src54[140] + src54[141] + src54[142] + src54[143] + src54[144] + src54[145] + src54[146] + src54[147] + src54[148] + src54[149] + src54[150] + src54[151] + src54[152] + src54[153] + src54[154] + src54[155] + src54[156] + src54[157] + src54[158] + src54[159] + src54[160] + src54[161])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127] + src55[128] + src55[129] + src55[130] + src55[131] + src55[132] + src55[133] + src55[134] + src55[135] + src55[136] + src55[137] + src55[138] + src55[139] + src55[140] + src55[141] + src55[142] + src55[143] + src55[144] + src55[145] + src55[146] + src55[147] + src55[148] + src55[149] + src55[150] + src55[151] + src55[152] + src55[153] + src55[154] + src55[155] + src55[156] + src55[157] + src55[158] + src55[159] + src55[160] + src55[161])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127] + src56[128] + src56[129] + src56[130] + src56[131] + src56[132] + src56[133] + src56[134] + src56[135] + src56[136] + src56[137] + src56[138] + src56[139] + src56[140] + src56[141] + src56[142] + src56[143] + src56[144] + src56[145] + src56[146] + src56[147] + src56[148] + src56[149] + src56[150] + src56[151] + src56[152] + src56[153] + src56[154] + src56[155] + src56[156] + src56[157] + src56[158] + src56[159] + src56[160] + src56[161])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127] + src57[128] + src57[129] + src57[130] + src57[131] + src57[132] + src57[133] + src57[134] + src57[135] + src57[136] + src57[137] + src57[138] + src57[139] + src57[140] + src57[141] + src57[142] + src57[143] + src57[144] + src57[145] + src57[146] + src57[147] + src57[148] + src57[149] + src57[150] + src57[151] + src57[152] + src57[153] + src57[154] + src57[155] + src57[156] + src57[157] + src57[158] + src57[159] + src57[160] + src57[161])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127] + src58[128] + src58[129] + src58[130] + src58[131] + src58[132] + src58[133] + src58[134] + src58[135] + src58[136] + src58[137] + src58[138] + src58[139] + src58[140] + src58[141] + src58[142] + src58[143] + src58[144] + src58[145] + src58[146] + src58[147] + src58[148] + src58[149] + src58[150] + src58[151] + src58[152] + src58[153] + src58[154] + src58[155] + src58[156] + src58[157] + src58[158] + src58[159] + src58[160] + src58[161])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127] + src59[128] + src59[129] + src59[130] + src59[131] + src59[132] + src59[133] + src59[134] + src59[135] + src59[136] + src59[137] + src59[138] + src59[139] + src59[140] + src59[141] + src59[142] + src59[143] + src59[144] + src59[145] + src59[146] + src59[147] + src59[148] + src59[149] + src59[150] + src59[151] + src59[152] + src59[153] + src59[154] + src59[155] + src59[156] + src59[157] + src59[158] + src59[159] + src59[160] + src59[161])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127] + src60[128] + src60[129] + src60[130] + src60[131] + src60[132] + src60[133] + src60[134] + src60[135] + src60[136] + src60[137] + src60[138] + src60[139] + src60[140] + src60[141] + src60[142] + src60[143] + src60[144] + src60[145] + src60[146] + src60[147] + src60[148] + src60[149] + src60[150] + src60[151] + src60[152] + src60[153] + src60[154] + src60[155] + src60[156] + src60[157] + src60[158] + src60[159] + src60[160] + src60[161])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127] + src61[128] + src61[129] + src61[130] + src61[131] + src61[132] + src61[133] + src61[134] + src61[135] + src61[136] + src61[137] + src61[138] + src61[139] + src61[140] + src61[141] + src61[142] + src61[143] + src61[144] + src61[145] + src61[146] + src61[147] + src61[148] + src61[149] + src61[150] + src61[151] + src61[152] + src61[153] + src61[154] + src61[155] + src61[156] + src61[157] + src61[158] + src61[159] + src61[160] + src61[161])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127] + src62[128] + src62[129] + src62[130] + src62[131] + src62[132] + src62[133] + src62[134] + src62[135] + src62[136] + src62[137] + src62[138] + src62[139] + src62[140] + src62[141] + src62[142] + src62[143] + src62[144] + src62[145] + src62[146] + src62[147] + src62[148] + src62[149] + src62[150] + src62[151] + src62[152] + src62[153] + src62[154] + src62[155] + src62[156] + src62[157] + src62[158] + src62[159] + src62[160] + src62[161])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127] + src63[128] + src63[129] + src63[130] + src63[131] + src63[132] + src63[133] + src63[134] + src63[135] + src63[136] + src63[137] + src63[138] + src63[139] + src63[140] + src63[141] + src63[142] + src63[143] + src63[144] + src63[145] + src63[146] + src63[147] + src63[148] + src63[149] + src63[150] + src63[151] + src63[152] + src63[153] + src63[154] + src63[155] + src63[156] + src63[157] + src63[158] + src63[159] + src63[160] + src63[161])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70) + ((dst71[0])<<71);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2c2a74a92ba9e81283fa9b0075e615921e724aff03ad8d170fbd998c88ef6c574ab584921a7c60696a065384666f2eb33e94258d5ca98ba33af3e4c46ae4385ab127cc4aa58a11d9d88003ecec8507a7e2898e7f2df8612ed1260bd0d4cb56f0805de511f5aabf9a5a500373c14938f8d9bacb52529fda14ec2f468a02af9499caf4450bf6ca6fe863c5d066479b56621e25458beb30e42e41f9e89622c0a6caacff7a6be63b61c5647c07e4b39a54b9b79666fd6d4e047f79c7717e31132a9c421033d51c36f0f1ae45587f8bc97732be3707196eeb5af9bada84daffbd32d041121886f1258d261d54648c4ca2a19c318645597fba7f360c90c5cfe1283f9ed60fccc95226e9b0e7ba34a5a607b666b352c229cace1be5698900606af98b600d2bbe086448eb6e09ca7b500942bbfa804c4caac2f936dd0aea8d9c99ffb95148a0c812e3624de2fcd4e8b639b73a8b8f96f6cd5b11573e0e17a3d10cc6181ea0a37e09d956aecde8156463e05d5d50d46918164badd4cea5d29cbd76aed892e45506f1cb223e628a53e19b7ec8477c7e6bd11cebec2965615992c17ac2ca29c0ecd4687ae25f132938c37dbb97c7e0146f6c56e86a5583599f3c4a92ae31b16791cf9dd5d52176aa5c922f0bf1c3e3f32e1d8a319813b340d2eea2ac54bda02053864cfb1fa2540fd9f8135c72009012bd2fa0dfecd9e124ad44599e80031508db90bf11c3501bd70f6a9a026f13380d4592b48296d45ea97e6b710c272936b56c5d868c492b0defcd9e72254b3867ca167e89a1735df08bf1fc1ea262525a6f9b959ccfad0f2ad83f8ff0870461a9819629af6d1108009bef94467966e93d8e59f8ca729e6429127ee512c5c6ef4830e3202d7ef681a80f994d420844980a728f22480990058444dd3e3d9b41517d3d14d3b2e07360dd2cb301d70f6fb2fe37db98c771922477dacac077d6b87f2f1d2bc1c933f60d905e62c1ff66ad2f90b54bd633954dfbf0795dfb6ff8109dd92671af2693ca1d5137938582aa9c6303317015e960e7df056468a73cbb527035be31c2ed0e8d0fa69ac648130d79c147b166b3e0a8d78c4037b9cb38842d05b686ff55d34b870dbb413201d38ca1edb72e3e9c3f967dd35b5bfe3af5855189c456191b6325213606a6fe28ad934fe53b37e0f0e456937919a2b1879b2d08144dc1b2c9766810d14a98eb59fe5ec6a93d61dc0e355733bdba9635ead1080bf19653b0b116f9d88db28aee8675b20e2e7e8f9161a074fbb95e92a5477b5892acdd8c0034f8a7477b16152eccfa0ef3a2a7cf651b891f4603e4b2b99532d362945915c61a85f7d5e9b1fba83f4d0b5756ec5bc5b6705106e4f877a9c0b76c91c9bb439f06a4e7a3300c7f713042261ae2a490c9b7964cb81df2ec133b12651cff04e29394140dfe403c6a0d370972eda5a6f0b5c8ee4be06275d68e2ce242bb5f5c893011cd6339b039267a7b5002d1204cafb07eb2b008a824e7af223e6554166b796f77f62a698e73cf52beabd3673d08d3b0dbf6c950ff830f7b4eadf6754e040c6011ba5c20423dbf0d15501639234cf0cd72e6f1e309cbfd091b333e88f447ab820d01888f404a8631649231b02604517c401f9da6675d8d177dd0ca8b262f31e5ee9667e41ba00403ed278a2dae4aef1e4752e0fa0a34160e2f824a1862921c52c6795ad12cafd01ac4119c4130e30da8bb01b045f84274424483dc85fbe61a309f88e119c8a9a241f90aefb4c3a7e3ab940554e701805db2e1f22251e2d8dd1bdce329b673e4d988a60b689c93ea5a9c0f38a9814863caa50799f3da3d95;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h20a653ad72a2b80b453bf31d4c7947b0bf1a7b259e201d22d2c62508e5bc97c99dcbb6e5463d7a6d410449344fc102630fdf5b38b2d42115733a17cfc44c7dd619326c270100a3ab5a267f712a1039819bf59435f0c5f3bc3c60fc5d86cd93c3df71a9a90e1827394a8ce6daaf100784086331127325627b3a81d2f48f76011e0f95ad4f823cba75a880f467e09e742fd26be8313393bbd5926efbf179f9b26f5133c0c12d4361bdc4d409d59c373363ccf0b439e09237d1028387c9c160d4c44e7f8b7e9340f82bafa97277d73014b806f6a5a69cc007a272be568a2e92ab3fc6c7056777dc960d70613e52ba0fee47c7e6ea5ec695a0700748cadb3c4f5825e610cf9ce5f455fe9f3313ab46bdac4fbd87ff35ad0ad7ba8ee117161a5988395f7077663f6e391132b2e1761d84101142fe885586a1c1490d04983ce96186d586e964f6095b9a4be358abe1ea6b39e2026ca2802f00df50db77cc2bf8a76113e022f859e89f8751c053e3d2440daea96fcdd434a54ffa056da29bdd8f4aa0150d69c4742b17e0e2910592dca2de3b4a5e0dc885291cd3b4c556289d63f8f2934ef1747e8d7f822d83b311dad60b53a0fc0a7482f3ed2332faba0ab540604da96313659e9e992e58ccc60932ca69be9fe428a9f62a8661989354ee8443c642c81dd697c921df0ddf50b5812c1ba01ac3f63bc895566f6297615046fed4c8ba17aee0a0126a05a41bb782e3a00cd2f8ad105235cddecafc7ffcfaaaee97b045223f3e0fb79a5223fef0a3eede71f2f2655ebb921a113ec25233627f8e7123ea9ed9850df410361fd3ac8856f196f4ecd80fbdb1b6d6b92f9711cf2394402a22ac5dd679a419a3b95f0bda0a94c2c5df5e25569dff3523f06bcd1f917f2c6c456ccb5c80e2c7a5da3ebd991e834123b3c919d65214f49680f5ea7800c1713032cc657c410cd12422240863c8bdd5772331a066289124a728b5c7804d5ff5041b2f0850c99085d70bc6fb639b3da7649bdfc4bf444b50ab0b90b66cbc3c1b61752ee5038e6c50893e5660e170fa0743ea03b307b660f8f624b5b9461f56b433852bad32d7e57d57b4a224f2712902a7e5ed97ababcb166388cdd1c060cd6eacb38175e4fa8e191e260d70d005c90e1be0046f04b9c11665cc7dc1d32970614e6a02e19d691000c4300f0b69edd521d78d7affa5ddf3b0e91d3632e51856eeb8830667c84a16e0a2748e5c0a369aea9e327b037577b50998e19d32bf85f8fd4e017ade7b85bb0ded43ec7c00dde06533778849bb8bc764b3e28903d038de336dd0bac0f308e6d66040d470f26c73561cec199ebb6ea695a0a4d6b814de21efbbef6caceb9f76ecbb2ad1560c0a1304b9e0c3541b52cbe7a739ca6be68031029e1752c11f3f25d8d6593634d2fbccd1277ca44b254e0761f182c0ad319067208b002c24e55191e764b776a1ff5057eba4fc411034d0ab484f5426b0c9398fb8912a73a8f5511bba5561aec6eb2593ba7bb86cdf77185c6be871a1235214b32b34c545be2ebca7e9a6149eac3008bc6ae0c210a63e8ad723a14e3ed3859fad5a12732a34d7f51ba9be4f06eb181dd0590b39535d07e30dd10a241de99432c1ff2f4a5e325245c168b5f59ed370da25198516263d99b8058b59b06ac9a663cbfc57dc3ab88e993eab019bf3bcbe5acf0d8f1c74d539f08d394bdc105a43b1ad07624fc1f31ba07dc0759a24d3ec2772ffed2ef6f9b19a1c3598b156bfb04c5e85e14c3a2740c46876afd70e60797ccd9e79868a0644a3d5d7c887d43636316efaddf21fb92041db058b778853f5ce97216c8c29;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hb571f6eec9a5dc003a2b51b7cdb10b5cc6ee0fd3091e5afc1c48e148898a96fb1edca59e66254cee7129863001196ce47ea5bce0a62c5d92ef53093c42b9b96f19d8a0a031e72d9b74d226dd54b86b2e45cc23861bc112e80efdf4be61ce3c20e6fac31eeed5a75ed0c7b3cde2769a1a1ecf4010a46713fd8fe38cebedbdb62fccd8e3376e03f0ceeb849e98dbc0d44e3406199961b4499b4bad73a58c8c35718b982a8ff3b36b691c01567a2897e3aa02938a44aa0c1561b66593323a79e36c7c40b4592aa213e64f2de52746068407e2a2757b648d5f9fcf5ccff8732021b4fa85c0a4048dae67c02561a3e7ab2e690860a9f442b7dcd3cd14840eb32cdd9feb00b9e9f4fe1f84704ebf09533bf81338b8e208c83b7a7300674feaa433aa9671039cd8009829fea95db4c02f1631a1062c3a09041a4ae623fdec8e83cab6673d205d3d6e2dbbe2fb592bb78016070531fc02fddebccf98d8aec89f9047125d3f7d7d35ca5c45a0600bcc3e93fba1fcef19f71f065ecbc9f5fb9ffe32ced7c15feaf805a0337ee83a87e84aef42c41b0cb55009e746196eadfe9e80413810f8efea91b2d12294fd22df1f37ca8ced9525f6f35c3c6ce0c07c62316d05a72e5d0949006740ea99d5d01def72ff4eca210d84d79cf8d66eca8892538fa4f231377608f1dc093b6fd3a81d6fe7e2962fa1b9eff4d70bd8aef1d5fbcedae14455692d02bb5b3a95eced1df712926326c4da1c96643e83646488770b54abe4b89eb0dee59b5f1ca5176ebea8b52aff3857167d6e8d7aba909fdfea6d38d1440aab5e9fff2f75c6515a8ae1c733c3ddc738a6be7769c0e3cfbd35cb7efc02bec5fb6414363ca5380d81e811a22fa40ca6949e7540adef2a0e11ab1fa6c816d7a9e0c480df8d83f2b6d7c5e9d474b2d3e8a01ef7d77d14e0ccc21a97b700632705077667f9fe86f87cb208a73491df7cda2708bfd19947bac36db69b6486073b909a60d18d77bcd68c8879e1748aea644039a353fc9a0fa75ace619db613635279a60d0e24467c7e40cef84be16e2dfcadd0a1843c5c70d9215ee765cbf16a0f0d7667c6290d1fbf6ae0e9b16f5aa7c0467cee2012865061b5b4fb08f42d7221513226223c68b14420a9968b64278f8aefd3705f47c176be062276770752efe981da74d8bd56256add4ffc527e241721064025e6977871e736e35b6433bec042b4f564120969916ed883175e4642615ae2108c956b5e2172a60320ae084187ed1e3a3417ca553cc1bcf2451470b9703619418d6db51f4ffeefd2a7e7732d04d27ab42872b692134b9ce3694a198a0a6d9525816dcaa7d3c9dd6635286ce1e8738637b805869359326ae1e707e29162470fc4f5bc694e3b984e8891dbaacd3030a2ed25c9323d49438c41a29e7c557042721f89df9020ffd264cb566106189e72804336fbdaf1247efaac18f3d13a8c72197779e7af2754626002d7c270e1b4ae5531f6a03c3c3b388569b2a25bf699cb5921f2ea748424548498a35373f8db762752bd0fea82b7de5436fdd83015d06ba29089c508a6c9d3a80367dfc6d43dfc7cdafd5b53d612511591f659ddcddcab8bea37a0bfaca2409e87143dbc4eb786466299610235b576e7bd7929665a8cd7d2e12c38973da37148f4f5944ee12d1367741a736b471a8b6564c572f92be1b42feb052f2f211d58f7fa8f12958e605425fd3c235983415a31281d466e364460959a31e7ebd5a523d0f6ca396d1dba13807e5c58b55eff1afd5918c385bb78bb938d2b474c1d51d23543127791e18a39a4d06cdf518bef24ace8d17ff8aeb28a428c44;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h4584e6345f5ee01a760930c441e638fa961831bc4e98cb2e8739cbd9a76fc614d6fcb6ac6977840123fd358f42e35341d6377582b66033430dba6f2589bcb8a2a7c746d8be7dabd92fa25632d7e0bcc42dd68ab0e2179527c02c7221451913c779cbbd24809fcc0a2bb8ca3fb482573fa15f3833f61d83037b565cb9f8a1a2147bc4bde86e3a7a73c6ddd267212909a6e4e03fad4c289f689f25412cf467784e40f839dfb683254d1dff63abc6cf234308bfbaba594d83e97ae08f9a6285e4a06d270a6de75b018b457066e2c453f0a8d1ca53bd5a3384a0c08ee48ca35b31a1b07b3fb2c5f02d5ddb0cb9b555e109cff6a5b261c94a0af35599815891449cf34ea94a1bd5596a8b2bfec3551af39417a2b6ff8dfb1e749551665f2604e544018eef144081a1947161e9166e2d1798cf9e4b5d74d951061f1462f959b945b68839519a41656aba3db44a67f0c1122db37123c1cc6a130102cc54ffa5950b93c87ca69e8163ccf3de222156d2c65b594bda0d69b35b66ee38c7fe0364447624ae9fd24c259f1a496d3c1e1a223b71fc68e5644d81722e26d623206118dd2cce4c9d08292824378d6a246f743474df6ebfd9a4901404c049c98e8b881e7f661e0d0248a97b475aada5accabbb065c5b9b21eed6a200a58e4f59890a384d67497a6cd30ad2f039a69afb101138a378fee565ba74dc6b6f15135199ac032c58570cf09ac4808da331261039049da3913266ba048d51b30dc3b9287d38efdf81b2a301b79b834c49accf058967cd48c734bfd2d3aa34b2ab90ba90e0bbb69fb9aa133daa0d1df0762680b1b27a8dc62dc64a77b7202e433fbe6f1ab2041ce5ee31a007265cf796d75f4bd1f4d024d4b384596ac7981799b4f9339f29faec711ad51f058e295d5e3cdf74f1b2e514ce5e507fe783832689b38cba1b478473d6b6c283566cac546a7c0130837c896c86ae23ea3d8b1d0d460b39d2899ead5437f6f6c1e8cb76600d053bdfbbd5b98b9127887df1c7fa02598391dbfe7c599448ccfb9d1ffd557107c6cf44bd99b8b3eb6c72edcdb1997987b1e5a77370050990735d9e3bb26a6a1ef321d18ba40f62f625483d1e09339f0bce03ce10418155d33cd0c087b878b991618e3e6d3219437de96469bacdaa52f6b2b9b07d3ba4305ada2270124c9c41ac747cabf7294daebdbca2d8b81c1a67664cbbd6839f37ba80b404276cdc4bad7838841aa67e20875adafe5abf671f04743ffcbf889055b4f85bf62381bea9bfd240e966c2da132afcfa52ad3d7b820a4b569a0f78bcc05e03dce1a22b8a52ffbf7d257e869c6bbff6bb10a99da186cd0ee70104a9d74163b1b36423bf18f32e62b86f64376b961708b941909167501fcf4e99368528f63907cf2ac07ace6c8d94b6577678f94f85089895ddb78b6452382313b02c672074102ce4a46fafb909a4e03d23b6dd4b5f8e8aeace79f6ad7f2ac50b617b796744b2394c301d2ade933a63656286e73e36cc137a235a884470c61e24b8e589409207b7faf7f55f8c838bb661270ad673e3c2456beb71f4a376d2dad6ca48a4bc41d4da36b3895ce246a6c931ce2e2352db6c38fb096ff100d8667c0426e0979e13c2ee5f58cc26156daccdb54456aab449d03433bf07794750d30abe281b5f354d1a2ac53bd27d1b29fd7b4ed2516a46253b99e966fd1c7eed55e5c4ecd44aa569089bd2a34162d09075bf7a70660c2f6247d4dbf8f88b68d18bcc7315ea38c9aff1b0c3773fdfc7015a04de088422b821322e114ba3cdd3497274464d9ec6f2cca34856490aeb1a5f7d2baa0c54300d859cdd91adb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h735d8c1ce94b80f78fa94e7141006307c5952dd337fabc944261a70a0d705c0199c1c4a208b04041552526113cb0a860da7414c4397be2830a373ecf95565c79c972fa5d993f6c8e86c86c394851530b4ade36f3c537c1ed0071d4498e6a88522138b1fa4660e4d36d48da9a030b9456a460a189b9291dd81dac033ba378436acaec02d54abeb6eb2f4d82444e256b4d98b5591087a0db3b3e97b5d6cebfca1dc50de3ec80280dc4ee74be77486a9f556b18790110c47ddad89ec162a437127f180005db81894edb3421bda6697b16d7ff182be5a146cdf1f4d5ed1639a49ca49b2cb289d504dce909e3db95249552515f2bf29143f81ea27c56689ccb2d288e2164358ebdae5a0c68754bc81c7af0b89c736d735d1149dea5e47af103588e6d0b657d16e452a335fa3615dc2dc487bdf7a0dd50bc71958531139355e9144b014d3c40f923cfa7be5c2caccbafae3b11b8034756b021f382a781f6cd289833c4e0888d9a2b306671dced5145811d0d92fe77d40a8e2a2a1f4f1aa1f5c182074c241eebeba2c04a59edb441233e3070cf70060ea4eb3b1283dbe99bc554247d96b285f0f91456812ce734268d29c915752df1b9a3926caf76e23a52ef95dc2c03ce2a0423609ce5e0ac88bb7a9725073e4c79f77c823f58c3a7977b8a978200cd64161613310b0cff23a1cbe39f0abcf314e1ec6235d29a399133c82b42fb535f06c22bd92ce0b6b288d5fceaf138640f5906395d8fae8ef0890be95bbd17bef56d383407e3de548740ed4ea93d3f0f2f4babb474513a58d4c04eed0ad8a8c2a3af52b9ee908825f99b96fa5958e493ceac10748d72bf1b712e21f3088a9a0f6a85a30c8cfe2370440823512fe1e2b278b56d0a588468a51219f9c38651ee7c756bf09a9a9fc3a6ad0144fd6c6d3af4405c9f85116178bdece0fa0f78695e48307a97695eec8d6815e161b8c56a85a4663de4c4c0359574b020c3584fb1eb2353f6b9e27db0a4c12e6e2b885afc471d9e18bfc7b615594054cd3bd18dc076bb1ea7516e0faaae75e2d6f950637276582868a06c83acd42f7c15585d345ac3422912336c5052d5955ed421531cd67617b9330814f2174c0b1cf1ff0ba6e55618da2d435e7abbd12bfe56c7cf28d650db38e80f35cd6ebeb6ed607e284327ec9205bff379a517f6a6c8bc41cdb4e51e4137609811c2d6cb30344a59ab6ee909ea9328336d471d90eb0edf35426f58c72e13e8efebfe1ae839079c12f1a792e127cb38919d826d71b563ab57e452c0ac130c393a608722378b6cec94b076418ccf55d877bf310e40470e2870a10b16636d041b572b7ed80eb3d3baf7e4df34a0859e4a093a32426feb354f405f4e0f4e87a4d921ae6f8f2485c2898b65d54172ebf49ffe2e4028df6a44a4bf4d90b0e499ea07f94da2d74f070d4591c09ad4650c567a13f0744485ac1ccb01ac8169b6d20133a96539fb609f058081e641d04b481b5163e67402f50e6763c82715129f67d97b525c34c4f8f3fb9a40e05de50cc9c6619a58f5cc8745533f6d2f0d9e331b93d314dffe10c8d6634a88ba4317870c4c673bc362298f1fd013cc9ab04a69ee091abcc49d64ee74d75937e8a23f57d231a235643e8d2dfd62a1df9dd00930878d91a98747755b651944eba4acd09ac53c3ccd30f683c2f5b56893870d425dc41a87806bf1124813ebf1f9f286625fc96c8ae1258aef0b11ca508d0ee7dc83b0e9f1ca97bcfcb5625fcf9868b084bedd3cbbe8684850e139213775d072283848d735269062712373d527135ca6c411399ba0df96d34264df1e4d234087b6d1858b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h6ec76607fc89f7b1d4c17d760ac80dc6bf42378db4bea70a29a605561f8ae00842e61e84e6950693c557d3c63a5374e8b03abc81758b2219de579df7c4dc104ed0b924650e077f8de1837b662e78b6c74b98d3e69ea24c211483d33a42c723924c2516304e280f2bce4b61caf9bfe802c612d524411c441bb3b877e693a7d6d8c5e1897383659832655034597ec970dfba3b8f1210cef9a447c76d0d0a74a8adcc5c6fbfb6ccccdf31368d4700935f03ba7d242904c1395dd836f0ac2dca726c6c9dca83266342abd95d7fd16ceba3b8a5be0631d8b51307819c8e754d4d27f6dc1dacb232d1e3690ae4954b519055ed24ee209e38172cb42acde9874d5dca551125c8fe00a36f0680b989cd9f007b6686eeb546e23ae769058e20e2395b608959cd870f2044e68ef061fd48604a29fd7e36e3451f00371c457f7a9099724a2e68995e4ebe7e05d5d81d05c3b9f71d71e776b7245470920fca5f89a02c083716ff39e95054d4ae41154224137492a0540fc0309d9809e3d43e73d3fe92f3fbac03af60a8f109a13072c65c3ecaf63a1ac54c0c1ed016c076d05a3a202fe6150648ebc84bdefdafc7c743db7b9f7a6ffe04b0f0f736528c26b0b03438449ba45a742edd9cab4fe340aa778c182f221de71da9076ebc24dc7264bbf967bd74f2352bae965f7f8291780e214393ff9639c9ff5d8612e8c2236437e2208d60aed7501f03ae312f78aa99abf626cc6f523f3543dc94fee1f74e43fbec309e5e80183c94c8b6fd77cf28e486c475ae415ec11fe1135149988903e00739cac5a0644985fadb13ffcd410a915850a52355944046530d93f0339764e5b30cfdba755352df554fdf6d6a627a76883615e1dd242d85af868b30b084f9e643efc02862623abf87c2ae1fc0a4cd25e5ec59a82109ba7195fee1969493078e10b2de6cb3bb24f3f23d98a34aa6a83dbee7763bdf1c046e4fbdbf1afbe19bae3d856c6bcce3af78214ef9e0bee99afa147d00744ac0e77cc34e8b7da95aafc6c84549f319489db20c95b0de5b9fc063d7f406eb2419564911638e8a20a88f0c359cb1a64ac0d121346055aef6db6128cf96f1fbf8980fdc5d65328d4cd596fce193a61a6a7a2d13f8b35f1d8b967faddb76e7228a2b6abf23318bf599c7bfb183e6d3fac907dd747da9f85b5bba0b9e19353cd51f43c6a537fbbb1d84e49927f68d355e35affae811a9bcd1abd61e3c84e4dcb71dd363c1af00f5945ea7ff364d1ed411388079dfc0963fa1e8c0e8eb5110ba3a3e3cd4edb729db160407480f3af07634a72f3fa343dafba7e6052ceedc1290a3b69b9ff9f55c91c525f61ac004c85c3e5236296029326ffe95c780caa8252cf57e50a8c817274ce99aea43e942c18a2ee4c10a01d05a0b5938e8eb1b97ae30cb4145ed4fb7a81ddd73daa6d1c38413500acf9226adc516f39edeff1349ab94585fea9ed732fe17a51492baf4f5bc4c68bcf06acc5442cd5e32ec30beeaf777a659c653c32e41c43acd529050f8b8ce1034d5b1e64a6583950d8cbe4f307a3090a0bb9b83bad3959a8a9c0f2277e4e1dac28babc379f42ed0381f7907d98068cdc8e6cdfbcd919d064c84d1029917fa9c6ff6d6a8a3b507d63aa881234d1fd2dfd5fd496aaeb9ce0603d006ecfd915e9209911684343ad423e2eacd0364ff6b29416cf9e37d0f3a800964b9433932c4888a0dd71560b2a140c94a8a49d52db6fdaca1e7f1a435c672278fa3319ce214abbbe991e4f9f8825a3cb0bb39f7ee9aa830fa5b710b210ecd76166f9d869440980f2456d191fd0bab76f1740bcacc19c488820cc8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h10e81a13d2c450f0f73bb57ac94faebfa69d8ba650d2b5e1104faeed802fafbc90965b17e7c62ce3b11f619deb107d013d707619d75461c0c22c39cd2a706bfe6e6574b0dd1621beb9e8839ac41470ac74261936623302545aa06ff027455322c02198e849e7151bfd556ee0208e0c8e7d8af391978dc9fd26cb763988f139bf45d36a4989a308ea1802f7c269229703879eb99d750626fb5e462085427d0a4b60c9754d4735b6a8179a88ab2af3534237bee480ebb0a41833e884a79ea6c210d568b62ec38239723b8b7a26b59e19e3034e0e64c339264b05d7468c68e9dcb2a2689d9b6ca420329f3f2eb145c051e8fe361bd09451c6973ee0f19abe30db6e1f721af5a2c83ce72e926cdac103257842eda4efa0cf60230d22b8cfc62a76121e9d2c1f0692f1e3e76f6c2bbe5e751d09037e30956c959db9a47d67fe8100ba9f18b022a1a902d93239d421e94159165dde23ef7dadda422f800d28a182a6edc1e294102068735b8cb224b710f29a0fdbe810538bc4adddbf3e33e7a2902c5884429c6bf4fa69c763ac900e7c1bed0ac483c93c473c987662e2311f1adca1c8b28be113f5c8b70fdf2c7e94b35643b5bfdb91e1091604bf1c49c9a8c9d5e27a20aa8f941c1bcb4829daf53fe7c38ba118be4ce4f3f0a6257b7d26612f7483b111e24e3641d224a2f175a1e17e8878fe8eafb34dd3e000523743ddf43630ff040c4b008feb75a7816d605eb9a58c907b36f274bc4ab821bac4de81d3d2f20e09a840ab35ae8289b13d7356645620108a417758f126900686d1eda994681a5b08bdeb747a729a585dda0c5ef6d9da7267d89449a25f5f6d12806da78142e47167480a8a22063e5727905bb2713e0ebfbb09a307a29d07723b237b611c2ce81f72d213977a317a54c8fa84ad41655e5228d23ed2577d34efeb582b6eeb647df8165ab2ab31762dc9f0870eba682340dbf90b583779621aea05fbdfcd75833f5214217c98b1b051dba499a30fd039304cbd7c83ad3bc48c147bf32ddcacdf0f8dca91c5bddbc6949d6e2e8967f0a4309b8eede84d33601321c6a90e3336e6ead4886cd7a950f69bd985e0b8b803deedb6a4fd82ad8ab5447915817bdf137c24d8e52227362740d701df5915903de41e85e340eaa48b23fc58f8b8c13bd0a0877738c70fab973cc621059aeb32136483305e3069c9011771405bc4526b4685dd46aa69f1ab585006e23b0bbd7d9bc26064f3d0246686e6161869fe607d4510bef7ea54eff5b4ca4e1a277b32e9f9aeaee1854e4c97c2e229f3ce4be9d369ba524085767e1f13e940ff75143580c945dd731f8de1141828b3ced5af9ec63a94e7a7ec96d3493ec141ff74acaed0951e67b0e2fdba78cdcb90ac9ec852c36b039f9923730b309aa913639e3dd1d3e85fbb7019e74f976727ee159ad3f25495402476d14fd3763751867f2394a2565dc67ca5581498d3ae171f5a5ea6948536cb0ebcc7d363c960872a1d1ba99ca2f44e393e464e68a9c4af2b753d4116d6175a98abd3f500ee3e8d2fe31eefb380c7550df7520d050e59a0f6eaca1a5cc4305852b7f3fe24a74810baddc611b08e160bc119e375027c84b157eefea844814da7984355322dcfa73eb2017850b0213d443f37ab6a1b959dfd1a9ff4a8aacf1d5be4acaa32a1a861e6c05f0c1a6cfc65c594aaa67a18415fadba50d98bdf16c656fa73a96e7274fa9e5f977001f736af2753a410c9f858c92af582a52efd66c3d5914725f7a41669bf5e98659326804c82a99aa93bbc89c552e255c5a489f77caf86cc6661b5348bc1991e950816ba40f74787eb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h31d291fcbd28659c68251f0b24335206d9dc2f4b38d57ff78cae2f410e03a6424ea7b29f02e787051058265910f1b9b537ef8f028a361d16e8223d10ba2fd01d1670b75ffbdf8979acf2ccb1dae50d0657d7579d2d433f667347061b6b42bca4deee23b3dcd8af2f396a6b296bc67814b38962a23cddb66854e5de10f5993233b00eaafdbdcab7996f2648dc47e1557fc1e7e4b4d9718b8766aa4ac35d146c2f2ca2436bbfda92e82db46ed8d417a67690001712e09971edf6b8ca30fd060aa5fdb9d8bed086821b5743a73eb83175d71e8b707ec5e585c4e253bf5064cd95c66c98ddeb95cfd1e6e9fedca6d86c115a8c96877b4fbee133ba5d9e42bcc70dc489e08781b80d70c6145af2e6ced9a6f215d308a53f4f1eb20dc1b94b5f7c12ce1856d94e21dfb5db70ed50724233b42d2a07ef7d95f405588e73f52faf5e7d0f855f190c373b30c0aa50cccd6acf6cd5d7ff5724e21747d0137fbfa49abd749f056c79ddf6b323932ae34ab3e47a3e57da197901a8552c5e0601bc91aab249842ab3ebf2a4eac01b87bf5270081d7ab2401fb60e2fc11b9d5fd50b205ac408f87f35489cf6d338544111971fc3d5ab38de3b54ca563cc87ad3d107b972684d48ad4e8f9535046510f8c3f3f623677e2d63202f2492c66744660bb4d3ccd6ac4a6789275959065f36fd16652227ea91595bac8811e7afaa492cb1061093a649dac5ed358259f1270b860e105bb66751185fb4fdaddd4536761de283abe63f4cf157fbdf4861d053bbcc166cab99f4e61a2559fd098ddd0b61c14a3baca7464b3d2dd26a616e0049ff3a9fa2d0c7d04ee80a7157fa9a484a5a34213bebc88afc24c2f10cd45495158031d4f2f6f88b14dd504eec705ded023df4939705858dfa5424ea2361ebe4f2382737734fd3204394a8515f69a06dc53d61fc07debd45828ffd8093fb17356452cbdecf9974fae2d71034c9ce9440964e1af4d0a621789a5816c48b5f769e7aef6c6739d825e6032221f91caba26c07306a2698b446af9c855149a0ec576b2758682d5de8d3590f74936c12f4844c01b72b7d2c4f044aefb695b4b858bdf6783ff7aa380ecd472a45b503987a8aec045734b9e21b6b131ed3dd9b49e751262e2feb57f402ba8355d36c744f4150c2b2c6d50cd4d2c36de0635c011c5bfee149384b1522f869c9b331b9376496063a152d9caf5d84a35a233ed7396d1c03da92f5ce6a12266e24e11bdf7f31fd4947a4fb6bf4d3ebd28786ccfa2986e4e45d9b6e178c4ee6f3ab0415117504b8acb66537ab10922bc753f877b823e02dc2f6b6f100f1425e55b44ba6b6f7fd6f544e1cb67899b95bc43a05961d6b898006a5b6b74033e13a51b89c06671d821c113cd8e5506cbde4c1801fdd3f31a34418aba70e8261fb8d1eafa50f38bc1b683e5683c6d2f4782b06feacf0ee40cb92bfba001c29ec42c85de91e97b0c05c6a2693676c47d0ce7dc564f3065a2a151128dcf3b5833511d72c77190d8ac3e8cc299a5c70a756cc33750b55a94810e4abc4668189af973763a5c29b98b3553a9a3bafe52e9275bcc9b061a8ddcfdf68bd3166ef059f13b5307aa2dc7ada1f53093bc1075a9d5d342d447cc624829064feba8001117da56bf4d09e105674d9da13da50022be18655a2455d8357251a5a20a0122bb84a54d37ebedba8c4a327e4beae7295c23468d8c2a404ba9623f3c87a0d3b9fedd81fd129b4c8f19808488225da0d9b1b034d069b5d91267228db9e6b81a2ce710d773eddd219e189b321afe3c7faf2e894f1ec4cf45a980c29a5efdf13698a294411aea3fedd6d35;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hf06494a85d1c391a7ea8b79513bdf6563aa87a1e1b6389d5f7ce7cac91decbecc671e7368576dcf9e4b0b17156186f56e36d039683026910f112bdb0f07d9b6230568816ff66f1f494c60088f2c63dc94acb8474b874ddec08cf3d58f8842f878ec1acb093a914a7e5e78f00100be89a0af0e7a99a2caedd6c5619ef15371604efab929ce7eda6581bc85714260335cb80da5fa81a4f94a452c30a129dbba3b4a452eeaba1feeab1f17ffa6e5f3eabcf988d338a8653008af764be03eac77b337323d5a7e8117c048d3269a179b83a0478e4ec186bc81b1e848d3ad0c7ee1150241652c974b5b0cf2d2b099e30d400535a4dab7699427dc47a4cd22b7542e92451be65a8ad20bdb0d11b62613b94bcbc3e9a4714955e232392523e03b337a9193ad1628f93be416d2337291710dc61155ae551e2529613b62ad05a9ecac1ff7c9ce6f085f52085477395deaf953b56b286727661139a6465e787beba2633c594c6862d00ba59ca225da4ed05a41f633d514bddf62ef1c04c6529b6ea1726d9b1eb34dc790274cda24d4918b0ea5cdd1c8e5113a5de6df38fc67769431791ca8293b39e098b77287017fc38009b3eba9451194a0e285648e07714de2f77ed0c83cf4d3c51c622fb07fe2c727d151f164220462170c74a02aef53cf9e7b8dc83c2efad530cf1fb0715ba976b8b769ce044b980f4f776713db3539f2d97c047c6934785e28daffe77b822cd2da4e262151479972113f4d116f43601d5cd08694cc3105f8a61c8f16af8d4c3d35e364d3925ccb48b2fbbef94f0666ec8766d29027bf18e67ae2013a03bf6dea3bc7ad67a90adcad1971265ed0dc072dedd37ef7665256a2c22cfab55fabe12b23be3f35dfc07986d7b4036ba7f2b16b27366ff746f9b14661a80f7f60149a972614f2c4f252f9ff70836edfcba52e1e65b7025be6fc9d5f2ae2b53cab46f82986c9c85ad760ba5b5aeda2bd9d229de51bd708f1a1d3058b0f2b33a6a513a20c76b4adbe4b4c37a337720facacebf63f84f68d2f7e32ff01c3c5cd73817fae20a740cf274569e9143a502b556a0440b896e2ed05b0d044cdbbf840a78a8b4799b3261545b0f2d0dbdc8f8456937048a135f510020c001c7fdc41635d148d11c7d5d7652f6c439a932883fdc9b84e0bfdd141cc70fc498d260d948df681c8b2e5430bbbeee69d1830053220f1f04eeccb889d3f00808964c2ff27245c064b5931d84f19cd7af17bce99b4e8cad12c6eac046ca0fa00af51966d8697a9653006f5f5e023dba7af771777aaeb5456da29212d626347f08a589badb8d0886392af31a8dda0f61888d85241731cc4c964205ede9ebb70388a7318401d86ab03691a22bca3b6e20b569c6c67f3b5112c7f280470b9a986db8ef94af26d758436dadc350a7c9c518b1914c795706d14e1bd4e7222cd90bc3bc0f7e4988320a3634ccde61e084a1403f12ef50e4568e336de8b59b7de53ce80fc532839cb4b9ad087257903aa6306077f66bb8d8e6a725532cd12bdccdbb9c80d724f318b5797e9b712b31b545d89acb64d7379952a9c5347cd0e413be2160ac51b15bf9d840d0987baf5c2937902a0e837ad5a17af8ee800c99a4f6ce62dac8a5cbeb65375ab7a431b7d6769940ddba5f62059d7054fa4eb00f8abb1b98555baeb95240a93a50e9937bfc03da707bcbf93090c8569a82c774932aa73c4a1fd4fceed8dfa421554658bec0444a86c74aa89020c90ff41a8dec6e3ac1ad9756dbc96ee0bd3ca1eb93a69da210d94bb3d45aedea6cfcf59c22fb74af12fbe99c355458d91e04f3e0773669034acb032484;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'he53af9be108f48f6f8bc68ce16d2e8aa47e302cbb43f31f125e372ddd53cca658bed948349fa63c2b258b9130b3a93dcb7692ac89500a36338331bfaf22e2f353aabd07b21f5846038a0b925ab5a4e34ce721e999d99ed07634737a4549531e90539d93ae178b1388b3e0b8d1251c3b78bb464ee32fe8534f2e77dfeb7bb5b47be158a35276959f0d7f414ff8584700ca43fa18929b31aa251ab0b235ed398505b7358f9ee119e3fe3b09f54a5d31efe8981e3bf807ec0dbbbb480f2b4fe34ce3ab3add8726d21b83b3cd951235bab1bd3ec37e299822b12bb2cbba2c706571ce7555d61c2439c95f63b687c607f6cf8d7932cec245c24413c9915f21300e10279f8993ef8e292e554bb43e570e70b42d4989c2ea63259b2271f384e6911a57f3d4a47eb7a5767d32a3f1e5908d6f2db6ddba70630a23b09a65e4bd9480622a85c5c9faea5fc29fe04d979462073557eb3749648050e45a8ba0133d292cbf1a78eeddad3f18d1eaffb34adbe9f53efa12689f08a189b4b8a051370901c44db0b99ac2eb93d74a0a131e712aaf60e2aa35ac31401b021acc02a89f487287e44b04ee4068d0d080b7de1b6109920fc60cfa331150a63c17ef4dd6dfba71488e4cb9b1da0c4e9f42c1c5bb4e7578f19e729827835407b66bff1e0bd6f464f647e807d449a59a9fdc4c65464998499d0f6bc480063b600d3ac6ebbdc57aa84adb690f135ad43c25da5771803f7bb29c6cbba87db69e7b6eb6fd2c651ffce41ac47537071533c124ef0b59b8f188bbecca7262ec4226c161856b6c0e92b01007db81095b1096738b6baf6fdf70e8ce81da873a0f8825ac0a5304da90085ad736c1c8cfd8503d8296d6a043873cb7b9a97192d74c4dabbb333ed4d1a4c98caa422efd97350a69d7d319050483777f34fa5566790c56dec3b9d7f252f8c6fa87c699a07e346ccc67f7698a73d31ec0e49cd94f7f1bc473617e73eb5eea7481dbfa7f4028f9d08ae1a74e8132bac1a8f07d5a68e065b860aa5afcbe292e30fb3d258f86d3790c274b047ba8073874564904c0e441f9a5b68387a61bc8d9b9710b79faec97ed9abcb5e9431b51901597ce7ac2f817bff823bc1727e7851f2a8fd46a1117f23cd4168375b56fb40d1bb2c63e11e0886637edb30ca0676773aa0c83523a9a3d6b1474113ac1980e6f7fbf3d4764bad14ed855cb5dcf0f1af21673a02be176001e5618b07172700b837a4d84ac386e85393423004c4b57d2a190df3abeb3ca01076286c1681f499d7088b44321835586867d0eedd3f17ec29b001cb034ac8e0a2eb0da7ea154bd26fe89e3e03cd30378069639386a47d53b6ceec196da268172c245e75434555d4252ae469e53dbacceb8915bcc7896d442b55da78671ef8ac19bbd9e1cb597ba7b7048968a9ac943e8e7830da8052b543957e1c69124bcacf6a5d468283079b13c79537ab2c5db00fba9fa7df04e581453d841eccf7994d16bd11c14053b19860486543f53f6a94313edec5f16a88ee87dfb898da26746445b65e3045055eef9dad93b833f375087f657c897d0b018806fa197adf17df1b88ee38abb271376f3466d4b93945284930183a5acfb71c378a390384f3e337db13a5b2077911e7435f6e93119a1eefbe4f7539049191d7222f94ddce8f271fab6c78dffff5764bad02d3c330896b16a4bb11d25ce4f093ed1075a8e9138015c404cc27e52e8c2fc636700aed839daac66b7e0abafa929ff174d6a227f02b389a2193cfdd6b676d58a24ee2bd3f07a80f57c3fa72bd3e3b431374588eb0d95432c3d6070c495af0e943e95ff7c57060624e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hbe087f76fcea826481d8fa5b75d122db9704431536adfac6d1bdb606e614ebb2313dd3f3225dd92fb3dfc3e68302e9abec895084177987f59255cd4af44766a0d49fded60086da4a375971da5a9291e9d5514dd9f1261dd0638b07ad2b5016201dc9e391c35fc590f004b4df3a65719f9ec73ac5749f0d01387d9e6ece229435fd2343dd3468d5c6dcb490f5feed9a4cb72b645c094dd0b63c4bf2b8f361a6ab404082f2f6187417cdb64c835b4b54bbce9258a73668c2e44fb57e50363954f47cdaee81c94d85eeff3c8880884da372bf573439f59c0e386d5a63b0b1737c516e94e56d52448252899c14b772ec4e82bc5d9ac78691424458a7ac52f2fe61591368a3dd9b53fe179b23129d71b361e855191d577d578181ab60e1ac38a3a4626314300489315984ded2b42a74e82d2a0e9b34eee9a406820b6feec826d19a4a6cda4bf3e11a6a66ce71097525c75d7488ec04d024bd95dbbc30a307176c4556627a04d99349d7bf5809e35a99bf5cfda2c0b06f2774214e434ddce4a9867c3e3689ced0e38c622816aa2ef1d8e0834b36a1490521cdaef23880387b803d5d9d72bbb1815ff17e9f57372600a977d93c4c4f67ceafac88add5a4eed4bb67f65cb9693931d2823d04546f90b0d1ea8d52a7aeaa6836783469433782ba10e96b9051cb32e9cb9efdc6842cb4960d256e633c3b62d4ff632e90d269cd7fef4d03643667cf894ef287b65ca040b0ee9262d2f9a2c56ca189951cec728b4f0e4015ad798a86a1471237b96301b50974d8bf10950f51188d1af57dacad1f482edff339d2f60b22556477085964c5221adc11f6dc8f3775876b12e16ca8b26a374dafa15bb2243c2f6c1d108c5c73db9351f97003e35d10906890f93cd89d06c1c377dadd48f24c5c34e77b5e160af34e1a1821cc9b6fa557b78d76af673378f209bc08b5436b22e118292a767c19520ba707b25f1081aea23af3d52ab61cccb0566c584a78e4e8296bc9c39ee2410dcc13e12b59a5644249b2eba2eb7db1931b22888a3559d70b22c8607fca0b3a2777c6f1a5235db0f6a6a1dc55ffd307e163d1fe5836bf94eddf35a05707025933c2793882046b693d95d68715c7e30253c4faa4e8a43a59c39560ef58d9759f841b4fe9c1c6f746e4ebdb5ca6312d4b74c838f477fa89d9039c2f22d34c7c4cd5e9484800a2a3db7d4d6474d69d6fbaaee10ae2186e74c054f8006b41cc88d8f1314a70304fc57bf823783d7ca86acefb6cebde0ad977b8008cb140ff9f4ec17c1768dfd8b388f3b71be2d6256c2009643d71172621b0ee25cb5b823febfb06711fe7e41704923881104fb64e70efcc5ce3a5adebc832145282a6e32deab55f62c5617bcd12f02e50075c416d49defeb0973a26379eb349a2bf0cb4c0ebe35ca2d2eab8a7924dda73636f6aab38ebf80da4a8523dc7f112ea19eba5049b0764257ec3d0da1b222a86b3cf697715a8b2e8aa7336d44ef71f931b32f76f220e80b0722730f3ee6b5039facbf04a331f60cf77c040f4bb9e0e168ef044f0d204cf706b3c360876ee95b53fd0ce94e9719f4e72881a7d2856a822461ae2311b7e805a5021eec5c6fe761f59f193b8ee6d0233962ee587aebccd071cfb39fab23294a9a2d7e31cdb1411e2614647bfe1161eda5b5580d9cf044780d67905af933e3baa74aa74891f940ee2680bc924c9148eeff7602988e8e8ddd747dca80bff33c9feb742f2656823af95eb472616cb40f98f4ae9165a4dd38cb0a169d2abe4b8606e001b5f6a16324e8b8b5e00a7a5fc95045c3eccfe04d9920045ea2a301777924ffa4dc87e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h553203d4a7a961e21cfe3e1fdeb6e5f181fb0561aece250cce6e125e1fd782ad46333ce3cf407916deb19090f0f0740db83d77ce211731d25b45bca57ebfcf117d4e49585d9018f34ddb1a53d160ef654ebf43448fdd950433a763a008f293e6f85881571aa87b5f8520c7812afe956918c404a9d4897c9baaed5b5cc04e51d7b16deaa0f8d4cc0ed7e04b9df8e7defa1bcd69a5d50487be2dfe7ca1512e95af2b9c2bd9c6b852e18bfd74daacb596c6c5742524a404efd00b1a1d21351e5fd802fbd54bf7b1942bb7c296491fd5cb1798ef4260b3ca6519ccbd402845d8439c86357526dbc8d49021d5a1e84ce2531e6c6668dad2c1212ada6331d7d03048c37b48bd36270ed8cdb910a606e74314ca1dd288c49439fc5a8830c3b3268ad120504bceb8cdc2831393507b3eca37a1eca0c75a7f269f10151785e05835f42842b62653a6158ca28fd09ebd1014888c0671acb85a919973cc5091a98e190d2f0be0116c7565e63c9889bc0d47eaebe1571cc5fa963f8b469807ad6cf07399a308f11139721f25d482fdd6a13db2ebb705878892c968520d51ffacc1a35d9ce0aea362114ebd81cebc534d5edc640c34943d9023015424d680d012b6f50f044ee7bfaae17662546b0a0d3833cbfee94e1eadb4c11df6f8e1c9496b4df2d71472d88c85776f5df3513d9c86ee595df970e780e656cc1adf49113057b5c828812ab2158922c72e661f98db663e0c690e6f0d78860102e8b870721cf92d998779c2d3417ad06f1d384a66a1ef883a50d5e796b706db2b320ddf20dfd3771c78e750acd8b6741e639b3d34040550028fa001feee85d12946024f2192fa032866c4d10d40b07b87982897e0989b92c7737fa7d730a0d376e2b2bd707d102b35f0404c7aa0650fcb83353cde91d863a957fabaa0d3df8007ae1605e9a3ebf2bb07ffdcd92a1c3e82ff072be87ba4b29f160a99be2e3072648acda20d151711e87bb1ec1f8ff68a4af94e6dddb190ddb0df500b62a793b6d28f275536ebc1c3cbbdcc7d627e07bb5ced7fb2981c968f70b26322c2a8ab6a20a654857887009bac9fea6d503d9ed652450ddcb5ca8c70aa0f59b4df30997b9fa42d25415c6333a1ee14de895ab81d44e7c5df720d1de32154b1ab20e9d5e23c5348bde5acc54f5630c54182f7053bafa7163fa7ccc55c0c206fa9ee30e2bf3d9436ae48044ff1e1b47418b12615814e82802da5a70ab139dc0b49a904808d0551eea12197bb8b389e23c79532cbd8895e5d97c4c02b756b323e6ce5ca99d3f6336750ba9c42555f382b5dc037e5c827359cd35da3b95901e756e323a3764081532d2c798bb8f57c0d659fbe085381f36ca0daf77f1d2e418c9fdcc519912a0cf30971a43dd40c3937a8eab5b7cb7ff07b3920d59ec5fb4e123714854b085848101bc761d8bfe47a16d56513d6ed1c0c715b2360a36dce80d19b1081ba4ee1ba4338f4e43f01aaaf94c23fd1a1897a1ed9c7c8d9142da66045aba49aecc83b126f65ff9ebbf82e650c147cb28566b5de93de537a98f5ffc9aa24c5875e043ba0078be4533157fb3fe4c47602bae4426db18802556887fdf8054809439611d9381b8f1a521180cc481fc058a14db22e12332b15ced6af721c8779fe5c9de13cfb66df4019fb50ac30b040953e08031001ad77fdfc142a1a2b2d80ca7a44141d8e7b381f1ba77d2d51c6a682a128debea0892bd2a9fafeff5b9479d20159a8a1b1b12f2c036ca878ef178183401e49e3b4cfa1e6f472b98e01086ed7ff9e8d2e33c0769f51e074334cf2af4b9e7bdfcba894cb419310fb0a8c6f9de20a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h144d5fe4b158658e6f4d3dfd9866df99fa8018d71ee446fb76086f5bc6989b138892cd6e088a1f89ee864d03ed7ea57153a40b42d8c0ef8fa315db305ab757f4c5a6e988c32cfd93895d14e9606ad285a2c693bc177353888bfcca5506ac7e8824a7e17452fd3588af252f8013d8761a8ccbb72b6bb317e51dd2b13fd2ab50e6ebb2e76d97135b5bb41c8c4c177cbb86ca4918f9f2af4c050b021260e3815ab7c61fcad41f94df374fbc8d6ce9f99f6de6b815da536ab3ac37ea7f054b5c5bdad2645055137a262cf3e2949940e506f06edaf4138620d92dda3d4c46a2f0079037d304e2d813135f944a78ed70818d5c6f35e9e9cf97b8eef155c2854c5f954d149d623d31bd3d6b40f9eb5e5ea34e14ca4f760982274c72f2b323999cc8161b5cedc7bf2591703a38ef61b20898e8d70de0ac1fc2fa460e7d98a9651fa33696cccce0acd8ccbdaf8ff69c05103ec101de1c79fa6dcba2436f9d0a8a028147853cb6908c79fe1c52f5aab4a9d5bc269d3fd9e91717f75236e33f119f1c456c2d98e356610f8cca60371e0bb3fc96a6447a4cea57520ae2911b1cea994c03d61bd549c76b6c1999de3e0696911f0ba16f3ca4890517eac8ff695fc8d45f9ef08c51044d4fe4dd8f4c9a5e84d3cfe1d6c5635691064e5866078c86ea03d2f2dbe0ea73455c51a49b218ec15757bb90ee28c70b3fe7457defe486c005514ce0f197cf94444ba7cdb2931f151b77a97a6732a5cd4e2e61d53010aadec411db01fe58194171ad66746daee0b4f4116154886f11073fb658ddf48057231525c01bf7d67549438e21ef7b560872ddf5682ff10826afbdc22fc6c89d9fb068ebcd39b8c83213726e1ffff0a7b9f4eb4d3dd8dd552bdb3ca77d01c5e35a6fc12a2f34f79c505f452e76f50d9beb7dbf657c9e47c161936b11585e68e04540133a32e58e4965ce6a584d1bbc7c6470cb38cd56d939baee74398ce9a52690b12d8205158d5c6de40b9d9a15d253c47b57c1d2766b5031df4bac8a87b2e33798fb4cd25d6080607a324cadd2926df710a2e0d4a0e28f34d347a751b849f130bc68d2e6a30b1a872f5114208833dca1da18ccf7c7844a225bc768bd6372889210b48b0eb2475cd05fd3327fc80e02b7c00500e2576abb48fb28f4cd5ff593f0ef05c09a29a19f9600aa160199d9e6c1467c2508407ca80a6f1738b4d004cb90e0ad6283f3dd92fd26c75fcbfd19e162649681d0d93b1f3ddfbc0beb11b8adb1dddb8cafbe2cd3178b2046d80f12cddd212f867dc2225790e449ec22b2fd4e9ddf8b5d6f479e6113175c03173dfdd440dd5a330c64f5a169db9992711e65c83f6901d083c15ff97f8ff8459edffa98c85adcc1afb3339a789ac08c762dcbfdf1faf04712751b31a9367f8a98fe51faeee62bc3d5bba3a3bcbf7ee79a9e3271ba669c4604599e2013eb98ec4b517288e09b8f49fc52b52a496240fa6aec2a622eed373c6f63b56fbd791971306900cf7ca6a12d58d304b261e9618783295fd1dbbfef0d3f117645c0dd2847c98da733ffc7cbfa105b34564e64cf0c97ea6ba820c621002a946e63617d9115295c8e9d971cd9510a5d8a129d11f667cade71d63938f17115997b65e94e43fd97f9815cb2256b9831bd4e0eafc559e91ca0d8f832d324f9eee2cae3051f2bcbd69eb3e6864345f8ada6c1d251e343f1253a43b3b0b7268ebfd4c345a38aa17c048e0fd0132c140aeec05109471d4ae194ce138d647e937542e9d02f44ae523bd6e72188bbbbc72367419ac8d253d7444ca118d16279392f2daa112aa06405f1304dfa8133d7c78194407a6a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hccd9a5baaaabc049f5bbdc49994a700d4ac4cbbfbe9b35f6b3878ea136b57ce0301f664d5a1d3f93beca00c5eb04277d1c0b3b0fa7d3ad3c03b56afbba5a5bb50e91614d632dd62c656da8a1c26dd494f3ab6215afc4ab5daace47b9f5a86f2762294b7efd07910276095d7a7aecd0a93282b8cc17cf0c69532add4e61593dfc7c2bc26a05b8f9305ebfb4e77aa045a0a2e9cf872dd309a6c0b9ee3a18ca5120b9fece584f00e0d3433dbfca40cff355f8c5dc043100b8b6d69c73b1065776ec382aa0e5fe80d0cafeebbe44dcd26053b9d2d933a63d62cde0785977a2f88465e264a5eeae243fdd6f46415b082c7f465accbb4583cdb5cb7f9549aad55ac911196cf1aca364e45ccaf1a17b50ecc138f123663a634f833713ada06ba13588fdd33cf5efcf83b7bf2cf06a1997a9d291c4bafec2cd19dcbf3dac627f208abe9514c67c5b35557702313c025a4286b3d26dc4fee08fb4dbbb9a996831a03cc5fbd687c7f700578b5088f19ffe80bfb8465f57f1264b37f211360a19b6220d6aaabbd1ecb89d831fe46ca0784f128650e9d54618a57336e7008b440e3b6c1111c11b196eca1463c78ae35bb984a5a19ea6ece92aea3c69f844254d7e595b557c3f626d8608aadd5a754bddc23d3b7ba842699a0e177295d886d2814f12142e9171070c1c27c34b263eb3074e64a38fca2a04860777299316e317918587998f773d36af87306d8df976564ef7cd1cae6efb746dc3dc706de163abfa286af7474014100216453042baecd51725d04ce9bafb87c19da3344b0c0e7e5c45fab1131c37f66eb94e7dc6267f174cb164b618b8d959b1e67498fe95f4385dd81ef793008192e67989b5480578370484aeaf6c57414e17287939da4b1ef63a2db930ec899e3892355cf48291b7800e9dcd3ac49b700e840879dec9ea761ea38b8e3fbc2b90ce5bd1dec81927df6214f062299a96847494d7b8345d7284475aaf138baadda25bc4d357a2b59bf543e5a87687939de0a2d484f4ef314829e09f47bf7736b8bdbc6c53b0482b534bf59458bcab0d7e8b06e0f111ab2b63824cbedfcfb848f524920e067be8d4cb6b9e7f93369043dc9329a7dcfbbbc297c8b79404da5309bab5c271688d62173852ac51d318325bb0a7240cdc71959785866ec79059d53bd036c396f323a87acde0ce6577fc9534301c22a07edcb1da690e4a923548dd5f66118a7803d2bce74d04bfbb5a23bcc8061c608de1eb6493953bd979a84b00d2524a1034f4dd1ea9d8004af450332ebeaafcf3009b63a8daa7c7b2972d8e4821868069a0312ca2a71e1b555b0b197bfcb6b7effc03290a6bb84d82a550e7e1dc5f2758b296d17f006d507422cda1138768fec2983219df3498bfccfe9862ebda7917b3c8aac973b4ca3183878e3877610580fae3232dfdaea6c22141661ec7945157581896966d4ed031b3d5bda934aa39b9a5215fa4e33aa5d3660fb5fca7a6d47f4a08f9babea720a2b37ae559d6cc51bb975c956713eda29da6beb69b8bcf34eeef9186a1d690eac79caddb07fb797f3f3b9e1fc064bade07a44d14e2d619edff9eb85ea5f384afa7071af9da8cb4a30367a40a1c172201688f7e31d57aa92e84c580d7ea0cd64bf40ec75d4ad59a4962a2c382c2336cd4aca858eee219088ed60c34bdc6cbd8e1b06bd41d844259e333801893faebd3d321e0dde07a84fd28719be810c18edf752feb32e2a705313b792d5521a1e9fdeb3a74ac97031d7f6d4f716e3ce679e5dd4615f6ee0b174913520ed9ee89873c72eb1b6c519c28b7fca8fcec4169e0750cff7c80d41a00970c5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8ad42fe4993369cb9a23e64c19e5f5037d0f8dc6407174353613ba2b5e79527c35ed2a5ef8fc6d53e3ef5affacbfe707f0f7dd612f65e5e17e3b1159e742f29f77995d2079d7b6f35ebfab91ace1f0cac5722dc5dcefc04bbcfbf9653210dcd863a1ee2a5263af32cddab67953ac920d0a2c28ec48cab17dede6bbbf7826073aa9fe50a071d7a368d6ad21ec8293ce18c0d436bccbbd2ff8766fd7f8df473bd15e08d05ebb6046afd0a46d2ec3bfaed5346d38fa3fe35dfa38fa34c6c0ed22f4a8ce722667588bd4d39df713f9a429f9bbcbc3ca62b87aacd0f48892244548c6b56d1b1d8afc0c654dc46c37dc97ade5bdad9205f213e2e3a1f580f1bddaa0dbdba10bb0c792a739de9f6c87268dc7600c95d2eef7286fa133a17b7ebc82658850785d68cc506cd373dfecb66754f3532b2ce8a369874aac120bb1cefc52b235627b943e9ebf27d5e26f58d1992cc968588b4d2df6243be59824baf1a8a2e47b577fdefb027f126c2c7507403d065bc23be7caff7768ea76eaee930a9e513f240b7e57a4925ed7b1198444ac86a7d0e0520c735b1ef1940931cee3f881c36e8e4aef6094529bbfdd3487ca33249757b6a6ef1b517b0ebaa91ea72da3c6f9675bc2a892c7b0b9b5b955a3a40ef8e05f1ac360aa7292d8b494a3f22ace5451544364f2d86a2c66ec12c355c3c47a26fb49e9735674362abb4648dddc851b55e4d6491b39de40909b5779515e09f09f0213b7365b94ba4af31c9602ef4cf67a870d690f07ec8d3eef4ba603ab468f2e8d55c34c489552e4dd54bd9c87da9af278577d58f3991900065e0cba553846397f1e65a3767321d8a32653004857b481bb6d85a1084b0f36c29a4e389b1f83453f1a6386bba4cde7f17796ed427f44cdd842394d6924a85a844aa243326bcfd3d31f72a887bc0a4b9295479c1224fe208375d5a60ab769e0ae593955ef51ecaa0892b14b615a37bb89d307255597d744223f7c130378e914cdb82593ba4769c82095a3132f0dc969c5b638c1d3ff910e37a47ae899e41f5e9718fec2d32ce4506feac097b3f668c1953f02a91b4b7059eff85de05309f458f05af82d45e91e50d15de9ce72219f3b35ac5fd9c5accbcfe206a4489e060d43047046b69d62d5cafe431a122e8cf6b865bd5e0ead134b7f25d3c7058e50ec6c9095c68bac7943c6b67993d3664ba74046c07b59fe3d7bc68195c95c9f8b2e33aa1813b6ec4837b23cb709cb7250eeb19b484e4ed85923f6679b6d6b67e54a0cf9b85e9d550c5bc0cacc683693d0b181b5799123b631e3d5e1ef5cd5edd707b57a09170b7f0a956d23fc4d0e1acb92835d359605d9663d46fb36853dde1058f958ae17a6088ad5bd794aedfe41a7c92361f033aee899af407a927858f6243736f99b99ba8ab6d66f7ba06d2c1676c911660b2ee019eab237b17454817fe6f08a505f7c565eee3501f80d1852811bc7121c40b18dc5c46410e885540c42af344bb95c1fb7380d43a89159d7c5e6969d8f3a04801de3e39db75f7b49b0856816c49720d6b12c5484e257a83f9d15c49e0e28ac6642275f9202d1ca59e4cef542b3c6337805dcbc3f5888d552f35a2a473f7a6d6e3e676df99ec4c2b9510029af96e3b1343bf15ac14367178d172f28606f79c3072fedc0096c7d011d22571230da1d3b430e57ba5fab22fb8f597f28dca003129a46b8e0f3303b16a88d1721bb3f89f1c299713d165a9d257c59c3e787f99b922457485470e6df9d6d765de5e7e2a5ea1429b7f6c307e98c3a90f9e557c6ab4e082a4ef69d56ed37842fda7045dd9c6ead3970ed84bea442;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h4c4afe5e38f93ade2d3db0d8fcfd641ea6c5b1c4c3d640e0e70cb9167ce4e164db268fece4d9bb58ce7b7214960a3c7d832fe3562d5fef27385a5b5cbf79e00e77d6e9343c5f50dc881438cb7441e910910aae46fbb32f806035bd329bab73e7d420ade7cdaa029a001fc4d9d2733676c727be1fd3ceb83862c96d99ccb0af6582d80480d2bd9b2a5d0b7e824dd2355314da27940dcc0060dc5167611909320d69bb68c35965ffeae5a279005405babfc86ccd5e2d17afcaaebb77d757d50c71f55f07121b052ed67122fe7163500ed1842ef3aa7b20a5dff4ae6c255ba862d4e7c2b4f24a36d9fdd987445a5dab7edc7358c746c59cbb9f99fa8f264fa6bc846a584ed9f6c5e80d7c1b8482b13781d44330265ca1ded4980b23cab29f0ffc55f150121ac8815312add27b26b14a44c0a70ac0396e43677572286a5ffdb184c8732bb1bcdbadee62ae6196e1df5427bdf5dd3c78a43f5e085f1b58f715d3b9a1b1552ce44cd00179924f8e0f43b236b16e9e0a430dd37b72a619337c1cbbdaa9be8c21d78c608a5f89c0764b694ad3d1ea5be166a4fac010cec5fbe5bfa196154bf66d1d00dd7177a7c521a68a345d204689a1a5f45927f8894bb64dd83dab62f4114610fcbc52dfa714649a1c409b8b03dc1e76166fdfc296e38afaf8bbe4c7a4cbd25fb4629ae02e39bc88e84e74abb01e196ec6d7a963056aa17919ba6891ded6c92d3d2c19f22193371f98795cbf02e8ef18e67cc3a50540d0102615af75edfac3a9ca86859cd3e198224acd9023d375bb9816da67763eae9c845b1fc66b43e3f5789d083c41df4ec76bb2bce161ddc7c0df642fac28f33f6a8dc88ef8081f158ea645453ba39675c623ba78091004009b608c13d0aae5ed021eb7647cb01eeb43a2f218b235c84256d70d91d229bb086f10f2131bd08f856fbe3eab06e1db38be1f9301f08e39c526e18cc084c361e85239aca35f4ab54e37c570d95c2ecf8cbf1b15ce164ac08b7dc745a778d559be1a3a80039a3bed98902b1c08ab2b04b9912c14a895a7666145b0b606c8d9bc98658a222d20aa66042b4938e29b053d9c49ebd9884e1d1000098bb6dbbcc29d7d47066c8eff7127814ebe8836e0b49fbc81804768d3754bcfbe1268f4db499c8128d656790608e55c65d51392aa5292710881686edb5085bd57fd34e2c5c4982cf64ad5f5beaefeb99dc477c1efc09aeacfb5c872e14071b17f0e637a45ccdbf9b541b038068b02ab1af20a4630015184697bc76208c84f782fb0ee741ffa04c839e3fea72cb9d3622eee5f6fe9f2d114b1f56f7b5e62aef0e55e422600fc45a273a35504265f0eb143f4cf539c9e4f178ae2c7d2dcd539d236e431dd838e48d26690f3341985bf8bca2642546d3d4e6c76ffcbc7b692f20b3c6103669c0d32c1e4de71ef03ed5192eb2524ac353484901cb946abe7d18382c6a60e53b8701f68d6b47ab720a9c79fa6eb6f81fae8cfd5e0ee6697aa3394a51e32c3f2e124734b5f6b588936363c0dec480bc77eb0cb4fd41636a9834a0fcafc51b76c08d6dfae5346978658f71cb3036980297d8db0ad5e478481eb021ec6af5c588b0933a98342eb56a94db3c0e1e4b6faebc5cde8e437b11dd8f6e5187b1659ebab9404cb35f39c962a6f7c1c173a56a4901ab3946baf860cecab2d509ceb8e35a98c3b24c82571cb4648b8b2af3ab570e3a1be3bd50935fd7ac29548ec8d8c443513356865baf375b0ab77870dfa76f9e669a23f5c1312ee8b56addeba834af121bf9a236fc19569be5796f86d4dc6f70a9e385c2d6d980712f6220fe88f494f29e1fb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hdcb6e780c1841add59b2faac5cbae35e09e626926726efbe01445c2553cd3c793d2a93eba63a18596bd8c8662a842da8efb4233ce61030220d202d7c4cfa21903e75352a58cdf0955c911924ae74644e1b4ef77b1b87e234f8097ac994dd84125e36635695476c9f53e09e9c8d88152408eecc24f86d1ef590de14649e2705b6dda7b768ee771850a2cf011b911f9e5fe989987acb41230cd9fa747b38cb1f93b542c9bfd8716b41692b4efd77c76623826d77d00562625a3485b677776443577dd94761602d0498449846382deaa7ebffc1478319264abedd7b28d809fb608e07b7c29d5ef015346a26c7e05e7cdee45ee882fdffd27dcde8413fead2994bda6ba36a60d365d4d87cc153fc53238d0ec0750d80e4beebefea36ab0445081d50dc5bafcdc0ca25c5c5a59a84ca791486a985ccdab630d3439c5f612fbbc37b087385bb87d71b526108fe817ea96d7362194639c14d702c56b413fee4edeb1c1a72005563c22bced14c27339074ab28ed911a5609966ee7d2ff65b8091a0e95eff961309ee72077686fa6e35d49c231ae780ee46e25796bc62711c334abcc73d6d2b98d21ec6ed833fdf29b757e36a99fc43c4bc44e4ce68c8ada2ff5a72c5736da63ba443c42ece033056f10cdcf15193237210f8de993ca4721f5af4229cd0c1f5fbe4b5c66a197e81ec41db1d83b8acca962cee8ea0eb4bcdcd6f799bfef7a754e04df70cd01adcd8b2df622935f179858ec9830bf7a4f7824440bb3f4fbe00ae03b29f11239e817f4c121404087aec80dc7fbc42ce08cf6e405a0b89b02e59fead61043f875266b1af491df5857f7a5728507ce9fbd3df2700b4c63d73d73f5d8e6dc8ae97c73002e1c5c7074cf35eecb88ae94d414f607e0df10be6e412e77747fca280f1516eae3228b6a33d19b851ea4f3aa0107e19d73c5acc452d72aa714c34b6134b4ed40712e02937a94d80debe72d7529ec28e32f6134cdcefd497c497a070d00aef56687ccf0ddad3fc24cb2207823366946317848bc272f93730991fe576ab5b19c96e2b9fda82b06aaeb055bcdf7f405424b6323cfbf4f90acc811c5dae571e81f9838771649120f3b237c89b89208f4fd9c6839f72cac33e641d386ad4f052d8ec8aa3e50184cd9c27fd9d74dbe99616a4b72ed6af264ad22a8caef46e6718d9e859b92f8d10f217a45252b1fc79f6a726319e5b6cd57739ee215d61f048093de83d6d1e288a223b1e379c844b37441856be1366f7c0e76f373c0487ddc0c6fade36b0268a17d1a2f4df35861261b16eec60c15ce1274aef90a1b9efb359ea2f359a210c73d1b91fc842c9dc01dba3d0b23bf856272ba71ac1c80a4e29aad17bd457cf4b6fd2eb3c7e49ebfa1a6d592924b8af2c42bd2c2bbe94926b362f630b60902745f1e8439e394606cc7efee9272737d79845e27b8d0879ddfe62f08c06eb01bb5b18e6baaf2885a8d9835972fa12f28fc23c63e2f64b3d4b14035b6991434b517adbde3ca177054efabfbbbfbbd1fb71999d61db8b79f975f4d5a2e847a384e6f5085d36285cf4ca52a9273f9224838bb5e12a5c90f9b6adf6ced8ff0a26ea26b89dbac047b56f1f23645b80b286cbf5d17e3f110840a055d8625caf2d5e91d1dddad16b81ea334fc64deab590e0c16ba8b84cd0c83cc41b0b5236d193e82937d381064330bd78023497c44b0552dd6ebf0b7cfe47a2c033acb2f298ec0b236a7c00b3b4f65e71353e21c53781b7680dd761063a51913a39471722cef5aaffe10c53583ec9907f66e78c906395ccd91d1ca0e0313169b14d4f3858428d47d376a66e5cf41c7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h641370ea4a103b8eb916b4d2b18908bdf26d14cb5d1005890a46c6212e0acacd68024d4d96dbca5365a0ad8c2a197847e01fe40b46d108441afa2fc44aa3eebb70c0e8fb275ca2dbea98c5343405ab9d6da7c13be2bbb6b784643c61b53d577e5926e0d8cec6337dd07bce908e3e9cc64bd2896f4b714cfee2fb4609de3473b4a768d0148470a3db5d54c9dd102f545e1cba06144b616c621563d33cd155fd7009c030f2f9cf6498249f1281ece7fbbbea34279861cc3fcf0492b6fc6f676c1aa1e0ea803e644a2f7e839137b3c5317814db38bb67ba60a81a852a0c09dc77e008687149c0e06c9c157935399696ffc0406c8f110b03bc7c44111e2e807c5e9451452d16481cbf679954bcc940653d84366a5d299560968bed00edfe82a736f24de6c9da413f71395335c4860ad5c0e39a2ae29bd95befb76982c7b2f6b5a38338d9224924b8eb6fe96e55cb88f5f5a20209d62ad2db011ebf5c7d80b42d4a22528f4cacb1aa34919c26b1853a120b0e5e3abca9a08db08dcb51f6885ed6f532eb0530df9e8a616f31f6549be967164245a601b07c100294363aece5ecea303967d6e2b3acec2d9bfae116cb42df7f127d83f4bdb51d7dfba289f50e6aa7f2481c69262494f1dc4ab11bdddbffdc8000a5e01f1e94534fc0c79d33686dee5b15f133c5041ba716310f2f0d5afe99b91b1a3c7cc10e2c33108f99c9f80a5966c9ee5836d2f77aeecb0ee7d74fc1b1811839261a086235c637bb372f0a5eeb2aec973a0675af9bd588f2676f80a1f958e0b15b3219db021e7d0c0b1ec440a67c2b8e8b94d18dfffad035897508aa7467b139357eaf929f123526dfafd1d926cd03c850013097b63fcc370a3144128a882fe094e2506c63311e4dee332c3973867d120970e5009692b0d3227e71f647b43bcda09c33c2129ee6600fc0d6cfa88281b7fbbd170631f8808dcaafb659b3915baa73ec30fd5a4d121b98f73a641a759e7b2f3feb1b8ce8bac628db3972ebc76c94bddade9a12e3e2ef037617fcc5804261448eafd399223dc5b2287bf25db189d8f288757ee4dc94966c1b7b9911652da0e96940c68b31218ce6d99aad2de08abd572c46e1897ebd24b52930a4508b24259861270d0ba7e5515edc9d90b6bd794789d0374d578fbccf4890c7ee0cfdf64425ed9733db56ed1c55f59d3e7e24eee85010c3bee5afc7df803cce5786a907da2d6ebc198c27c8f093a266fe1e5e06549deac2f72db97b91fe3568e65889749f6fb8b235223272f1c948e241f5b25d45f9b23483feb97cfb881c9f07808dfb3565bb10efaf377e5afe55f59ca244838d2bf7f37765c0e7746464d62b85564ff25095a402afe5ddd4a1e4931ef9a268dc0930b295d0ac647311da963ab1d960cfd0c56fd29b5d45bd4fc9b1a5e2d8f51e194359c183e4ff4ea88b45959e1c8c1d3f142f04106f2a69fe7a754b06f645aafbfd539c9e6688910741c649281e8e5fbca910581e4415745f70bce644306236adf82cbcb2722bfe0b4069cde9d14abeb534f64a1d8a16dad6d03d75b00e22d89c1987f848ae0abf09b2b53825823555ef6e9b7c4c8a4b1490c2d8ea4d1f65deccb942bd1b6145f7202d7f29a6d6a8c2244ad5fc210af106e946e022ff54b1e83102166a1efeb53f099249228ee009782195effa5d52767c25d2f9c7ac38cfcae4c1b3e073d0dcda7e8de29df752a7c2f161488a3bd51e3332f3f26c360f392a3681cb1def5f740efed221a13b1217da4b43aefe66b49584189aae2f572aa609f11a2bd8468e6bc67f2ff29755092cef130fa856d3962d99e52eff283967a7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h494ca1f32d9868502429251f4f33b9e9d4ad1f02f3714b5c2eecf62fc8ea49a1898bfb06996fd06ef8b0bf9da039389cc2d61496fb36908fe6ebf432e6b0e8a2675d39b0ede6746ac717f37464c5a82acfecfda457566aacbac508e57025b14938e6718f1c2e5af6b803d4962150c71bff329ac32437e0dde214692fa750672b29807f61e1da17e44f0986687c4dcdaaac6d194675847ea9b7800981e1cd7a562893cc53f1cf523e88b93df9fd63b1782095a68f5a4ad112baff9454c7676c89da718ed26fdfaf0fdb7e5e2b02d043c72b9e605acfe1f78cc1a1e31d6e544cdb94bdb61ad9490d02046433f0214b2a3106b793a2f54de525e377e1c06f754a0e05acfff63902a57af38088640eaa44e4c4028922a3431fd37edb37703d8c0da266cab174c21a47b971f2a03ae79cda1c488406aebb6612de7ff27e15da865ad9b02076cb0c0342d857895fb8d854dc42bb2db2343de5a17d67ddd34c828a97de2506bb5d961d7719e98e6c7c6335199039eb727649bbd8c1f8afbf01ccbcf482a3e1cb8b71f4f4f0818c094fa15daf0c336a732dd95705395918f4343761c71576688694bada8cb1368bedb7609a3d5b9bf26a2740f2e3e9bc422c46197499298671ea6c143ccffdd32405e2ccf88b5c5beeefca1310cf18ac321560941157a196a42b89b28125debdcb1e5c108c4369d80260aecffc1857ba8d4ef899d25e929324563725fe33eae8f5786ceed75cdfc23af96f66c2bbdf17f583ca2c68cf12b49a381829cf73654b934bea553f8385f109d564613a94b14cd50e1363ed0d8e577b26df5a3227512eed7806d7d6f5824d97d3c2a56b74af4bc36889277ff5507ac8718237ca8aa0f453da97e5a157e2c5418d40ae2feb84c57d81290c5f8e68e67f96da7b11996d2d413e8c781b1acf1abe46092e17f0d312dfc55f959a8a6ee5b00c5800a713bf998251133859bcb60c3ba4a2f676f9c736ac2361f85df0a362fe33a3551c2cc06633911b2df027cc32204ac8983466a0e7cc99c3ec54bf5f667853d39bfce87ce13ce3e2612b1adcbe7117e44323b651a05b67eeab72c4db55b6bf5304ba463b70e707cd9cb85abcfef2e95dd91265c8fdba5c99d87f8169b069bb6455d82081133969dccc31508696afe7761aadcfad5af9156b810915925cc0e59a7ab28fbff0833c6f3c4ac147ba8a5b3d08bf6910912a933a48ee9a86fe482635b6f38c320ce44398602cfca68b25446f9b33303b62d28d839e152cdf757f5404060d7bd05df074d64574887cf0568ed3620253a5e727c77f38b79996c56cb9dc890b90dece9c71bffa208f4ac442a86134dca8bf5904bcaea11e0dc6db0c7ddc7739556d7162382b5950fef6551100eaedf718a4cad6b6659469e5acf3174ca76e7a0b28127d7304d7bdfb6cbed85b7b83a35a8b71ba1e56c8ef1678d2e440ababbdfcea0a60cc4fdc295a2d75757c97597247d84d5a4e40d693a94baddafe8562b495ecbaee56d15a5af550ce7415ed7406d81fecc40afd0c18b92a0040dcd9007f99f3d7d544456f9240e6d6e3d3fcd9e6cfd567df258cc44c6ac80180cd9a2704f5502b7b549db45719b1f5cbb4b981edc987bc23d54576510a71f27a7ee50e7292a286ec3c75c0e58830059d8d26c39edcf8443a6f81231f055083f7f3ad9d60cf5fec8952297c19c91e0f588e4c0f2681e7aa68941de6db62626d7f309a4532be217840adeec8b9d08720fd03b8d285d4b9fa2499b734e143dce50836b5b43db3c653deac8e7a105ec6acc063f234c264aa435329a34758b6233a91790cf7ba6f4a7dea2907738227f3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'ha4d4668180d06793a682b02a6ccdff39b94909ee357a15c86a1c636dbe179fc673c95f0fe1c5b02ab8f1d10dce3ff2b2506ac6d15a776a27f05d6f8b197e261a4370d9bc3a477a5f4fd24894244941870ded9dc4691b6294aeb46c2ebc7fbc89e924d378c3ebaf448396c03e1755c8b95a4c8e31301b8e1f194e3eb1bea137f63bbd57303aa7ad084ebde72faea4186d7210a0dfe10b94d6cba0102775ba5f3d7596560c5370e70451f750577d1e0248987cfd702e563b8e2915bca646b133a6a9ee8eab1f5e835b10efc4e0bf50a41877d448bf08043472af7f0fd7abc9e9101d56a7af0bcbb30a326a1cf2735981f7ee3d480b7b6055afe31d3e651d9f3645595027e5259b15dd23303ee7079ac0277ef85f5b581578596e06b533f8b385b2113ea8dc2b973623f0843788e3ef147af28d70fedf1b4933bd598490d6759be9a6091a08bd3c77d8a8879b7ee066c4bd49572217c87a816c9a08d4fbf6abf73a7f79efde9ea0506b817e3a3de820dbd9add6f86af7c823207cae23c707d393752feeb3ec9a24967ac7f369665616302ec11ad81be1501fec594b8f284b2690e7dbcc12a81a2a38df038fa2b09066a3d850726c910c0a3351ad24695d20b6d7d997cf0e630cbe8cc6b68c2070b120ea487cedabd5e2ca2f10ed0269791fe60fbbe0592077503590ae747c5fdbf2d5f36537d1d2d58018b9dec801f355c60b982963edbfc1282981f6c162b2b8dd57a7a154634cf6a27da3f7be305abaf89967557ee77208acd89cd6160e640cd9118bbf16b9eeacbe130d74494c20c3c52e5134de85654b22e17459f2273595abbd3d1919be097e7b66d2305b86146feec870a9ef6d6e2e622f98761ed40caa5b2284a509830e6985c942fbe755cede1af6f2a1a158c4032a2df8c1600cb0354170b7338ea2d6237b5fb36a9b4144ddc9931bc896280210e2fe43caaec536c9b38f1a1c75fc69c5482ecea479e827640af905d8178119a653cd21f28cb31a5114cf97de2a664e158b40b58be2787eb4879fe5da3e6ad4f68ab3d850cf355ac86c101b1735b87dd96ad8406f7a4a606a231670abef034e1ae805aa930df1dcf55d444d42a9d52b76f853586369b4e092877f05699ece08df5708816f322a11e6ff88272a9d8d9b5c944ca2f02f383e3220706bdaf3fc01da76bc7be8c770fddbbca4bacd6b22c920a065d178894a517bea030bb6e2f33a5d2b7034cf40bed71878047e605f59ecc72d376ce3917c2e3de9b22f1f1083cf7826094ee4564e3690e8daa1c729e0a2d37be77077a9b786f065366072432705fc3a00b3c83a359038acbc4cadc881436f4ee4288b79492b638115ec91e5bb0eef4721cd2620fd221781b65c38db1772aafe47a5597e59d2076104b2cc1625a6a8644b580cfb9c786a0644cede93f4c20aa10391d670a845cbc1bee9282181275642ed073916fecd6090a275583b64826e0a3833b913e69e182b661eee9cc15b5dcb1caaeb6151620f004c22c761ba6b6d713c9729c4b7de7933fc514bbb5411ecb4e73573e1b506d720e5e35b2c4af2ec4930235b2a36f2337b0e63cf1ed323831a34938c2e08cb06b27bdbc89a9a438c80b40bd1ba937ee946cb629bb255cfb321f7b4f0ef2f6ab22f45bb57c7dbb2d049726b1723b144d6491c6da5239d67f5b91431469c89233b57958cb8c5e5e36727268e4d5428d3a37571bc057e690067a39fbeb27bd6063bd75829e505542d5c2a69cf8fefe6ee6b4881a3bf81027fdfa3e2f932b8c15a0fb7deac15bc1bca893f2b9e6d010e03290adb5d0a13d3f78aa095fe4d172845d1689e69e3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h6ee38e79f20772235298069fdbceecdcb52887e0632cfd524fb5bd1278be469095f166d27ad7771802e218312e6ece55496ea761fa5f975221dcde662fa3071f2497a76ddc88f05efbd648c2414a5521e30097dd9c1bb710c816abcfbbc4f34ad0f8e89004955d55c059309d2f038d899e13cc027e0d3db0fe3abc8b7948df86985437fd2512102009f57322a6ef4964928ae4a766dd6076c8e09a717b34410fe8a5dab0bc0d6f536ae063c832ee7d66f424f50694de690c3720992c02fc1b13e65327a573288380295ba714ad73839585857769d9a44c083e9c7892a8be60231bd9e3c348f296f31a9b3f87f50df46b6493c5108d6ccd7b1a642c4a5ad51a0d6bd2b1f4599dfc45140e7e6e0c901b2278b2285369f8b5d5116454da58977b1694d61aa60b09669ed76e79580896e3651b6422aa2945142b5afaa5bd32a9620b189e1de9640f0dbbcd2870f6e208454f48d6fb03ab55423ae7a291c0bb5277bea95eccc803853a949d15ff94d8db9f638ba1c2054850e8cc4b2a621f2288ff72cca6a79e15a5e5b986ae226bdd4f19ef48223399ccee018f71ee9e29924f166d04e1fc65d5453948286acebb21b24b7f1547c3cb409483e81cb3d681e22d12a39db82f9ff1fbafda53587bb33ba3a38bd89c04ae1298e403b541d3beb5a1a28537d2fe629020a1db94786d0a5772a603b13b990e63a2892cc7411cb40ef64a405614b0cc3cc849132a3a2e10abdf43a8662bc88e803878f64661492715e1642f0e7433efc63b5a4f070dbaeb0c1210a81e89fc5e07c1d2418b423d614d1834523d85a1738464a7375e1500219e2a097604e720e80069e12e5b4e9fb123f04175c08802c18180ff4041cfc8fb6fadb2ad93a3d411dc916e39a2b8e1686254588dded589314778bd8f9dd410437013f0cc427ac59ae1f443a81150bc092a57b84fcb1dc8b608f46e93985217ebe411c5dea421b9807859c301a45c5cd1ad1161dc37db3ac989e67ea8a2d5eaf872051c87163aa8926fe6bfd6715f1d8478f2439ba58f590fed9298b514017d12cf6aee1fd9a13ce26d26eac0f8fa49d35c93da87976f32dfdaa9fa2e05d22864e1fc4958ca55f9b2a69d0c1609ff9e5c2545b4253188b43dc5e27b66d449a90872dd5be3657d5f176cf69a7055baee85c2a096373c6c771feac2be20197199d50848ff7ca04627b17ff8e2fc76edeeddee759d1507af86dfea692b7b0ee28d1b0c3203ab30aaf60dc6958ce6f20475dc65bdbc9d0a72a3a811435184f7b1af2abebd14fec49bdfc9f8f113652ad7b292d46af50206aec93f6a323602c582aa2f96bb440415838b194b9d3f04c87bc976a0c5549f27edc79c3ebdabf1d55e4641abfa97f2d9a6cc2bc5b4b4aa4aea032e1afec5ac872f08ba4f87efbd7bbe314ad434c3ae119e8e14ae543a9ab7d9342c529540791b960893bcb38be54ad12dbe7b81f38af37e61ceaf9967115aa15f804789f4436f142495e7cdc92d3446fe3fe4e79e34320e801d35c65563fc647274fbee7d139aad1f20f43308e20545d86215389396010afc0950b91527a5cf99627a383f909ab33860de0dff00b955d5c138ffdb0f78306b7bf31b49013d33ea02464854365dadf642c490a65c27ab6fbf86c079fa292ce0ce0880b9ed8dd16686a40e1290b944fe26ce380c4a455dbd5adb213596cec3945d7976c35b5dfd9057125243a107713e42d7de675b9d84e6ac615ff12957af461e248cd3ee2c771a2d68af57e1577fb84d57abce5b5ffa431f43367b60dde473943c1207c464c831b63715bafcaa0736c5267f49eabf52347f492cf19b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h838deeffaaecc3f2097732161f4c5d7d00a562293bd4e82312a399ca1f0b068f32a46e5a5024c0c53c56d90362749f9e5bc0fef6b039d3b385e75b53ef2fb301d1b1c82fd214ac154e915c58f0c4f889bc26be58bc284f6eaa176b73a23f681c9fab2a6afcc705be95001bbc4c5190a002b29295fcfb356824adb8f0ddb1831ab3038a2c90314e080ace4fb6bf2122f5acaf2afa1f1d5ae371cd93101904d71230dcb2a6041a7cc9c1a6eae57f21b5b27dc749825cf44f68acb4c63fde41cd5f3be7b7cf8411966e21ad953379829381a1424bfa31ea4349002c006698df0c281fb0a8aef79fc2c4ee7c5d637671ab3f20baa8a6b3cb0e4f18488368c124bade52a02cb199826ff1594282387329b9f7087845fc2b459cd36fc38f2a275dbc2d1c419aab4f1de40739ca4a90aa502fb3acede8f485d1848cc451287e3368e723dfff74aa0bd4af80e55d9355c8735bc42b8b76bd8e155c1e5dc187b7d45cb652a4230b63f32f94c50530e4dfa02d2f8c007cbd7561d8c7349565efe2f4e6ab0674cc67f4e1df780c6bdf51dcceef97d30be8eece24b55e1bc10400fc031c3ef3a1be0d12a1ec334f8b009a4146777d051cb80c10ce6f66669d8cf9848b6d09ea4458f78d566cef74917500e8709bad42d91f46947c8ccd68d3d137649644802a04576c1422efab4f092fe6b5f97c53f98a772baba35a28e144e745303c35fc4d05f2a86cc8777f52be8f6daaadc772af37d7396e2bca63498eedaa7b0285ac838f1a0d978fbcf41f239a5788f8191b65116a890e96559eb5db5ae4b2fa3aa695a3aaf238face34be3e8b021583103281e55e7d69284f132efc020127a812e267b6b87f63a81d7c2e51ef1aa91078609d25d3bcc401b06dbeda70c47b913e7cc49fb25c779cba8bc37e6c5a52bcb444681c2d6c5da7403fbb9f36abec352901fd120494b1c6e850e8fc9d36dbb6eed884b8e8ed3f2816701fc8474311169f536b5cee870839d64b15a2571b8670d9b38e4f4f76b676e197fe05670846911bb536c2f074771f09fea06bf97f7b644958e68142421e8236d2367073dfe69791a5f4d650bc20b92f250b4c2ee4d66daad0d41c3f9ff6230368dc48a33b0702cf9359fa3a3d836600b7c938c4b8d70fba1199d862ea0ca346391da3d80527fca8d29eaa89f718e014ee26118788a0985aa3742598a421fc83d43a3cd804efcbeeaf13dcc5b42f3507f64c48de6d854af51bfa37158b2881f9835956f1beff867fb11f44b0f7ba6f20d87dd61ca8bcf3acd20fc7b19a5dee81341bfbcdd46b44311edba190a31607202cc5cbe8f6d51f15ff5b65ae1e591afa9b053e5f9e6fa9419f470be4db101a01cca8e26a3d452c1e80dc99eee31dabdd82f48b74a069c0a8a1c04ebc5a90fbe059be2915dd7f2b1f96154c19e39dcc5f4536309f9b7c15745816b37309898fc3056a042adfe1538f6a1724e76a491fc32f6a5a7a237b2b6cfb6e6f0980b2d83a7eadd2ceb4c02c108b90928d1968a0bfbeb8b84d210b9e41b837e3f16de7b171ad7c431ee03192e3dc07269f8f7cd625fd6a44dc7eaa9ea27e7be23d28ee2367fe208c37a203cf3254151316efdaf1b13a70356d4b213cc8ceb518ccf36e74b78e098d39436a18e5cc38e4f136385a3ae42221bc7f54674fb35b5c9bcd25ce4c9157836df4ae48bee489c97c2389cab98b931b1b9b58e27d05e792a64fc6798c01262a1cc7f10b8e0da3d274959f3993c0ecbce78cdf794af29317e6a650106dd722731eea67d138cf162c1e6e160a06a1d7684f3bebcfb1e8994002fc794a95868cfe8cd4da0f3ba59;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8b6e04e959dee80285282e614a55bb612dab877ac48675a60b5c14de61e0e51be2c06cba50ffe49c0189986009988ec2d3f5781e6c4ba2f767cabdb9a8d18724261f4184d21a1de83c6b3d36e062ff914d2de7e828d52c556f3b6b7863010fbefb8085ef5ec862d299a7385959a9fcf4954b075e09174a187803021dff62b3626fc3bc31e4522e30c3b6e611509b3c8b6f5a20544c86642d18d941964adfc03cb83d08bfedddba4689dfe7104d8b0515e69cc848839f011008c95226e0f5c18055d94699ceb4de84260eaa58a88b1445caed6c4c2c17cd33f448f804a64b6045bac8b42bc5306ecd828c966e73efcc2732beb6423049bceb691be62d2bb8c7e85da8ba5a66bb61a8c886443158f63606cfba6cd6f7f4394bcf3cf3905faff3e63ebb86a4ab12ac34489aa79cd217baed32702a3701ca5c64c5904b694e32393a4efc709dc55b0bc2c766f26265fd4445eae3ec521fe0f1db0250fe8160199808cd8ed7fb5f504e26498453ee1016be4430291c0dc58e2fbfbfc06d233cc74e5abd912499eb2c03d4d286069c86f823ffef9d488b81a4496a97448251615e1b06096d1cbb6cb2a6a628bd9a14ee41188aa993741e1f3a7127dfc36ca0f460c898950da9c8924cebb640efc2c8c2ef45f8b7967262f6985e9ff0709a56ea1d319a26df3bf865ffb482457d651bc43714a34eb7e6066bdc854483fac41dcc0e8ecaa157f08845a8593a5361079146e3b9c8aaeca3969cdc65aa284a7aa6884d2e382a33ae55dc9f77d061725b21e2f3886ea2a64d49eab0ec912102688b04e66ed3ac295fbe40b6ffeb0f21dc0b40435db2a72e5780c17a68c7faa6e558464eb60a1c1b17dfe32463276ebb240fc7e4fb0292f04b30aca1a36179d2370afdc44e9ffc6ea89f5b9a9ddd2073910017c7aa030648772bdceb307f4073028bdd096d41d157becb636974223e31d862567a35749109c6574ec434303c328f4811b19409324f4fb8494d046ea58660440e7691b3c1ef70fc1e07e5439538cf2ee967233f3968574eb16593669dcbaa7bdaa2b001bbdbb37bf3886ab741483f8ec2e206a225cc97db50aaa7aa8437ce16e6a149e25fbe58deb8d40e310041f10b0a288138c322ba8699d753ed7bb775f217cfbd8b5ab511ca8e66fef86666838183cfddc324039afe8fd6ea1f6b46e5e1b3050f63536a07c66884429f47b04098df92176625661ad8b5215dcf09776906e33eef06746f122893b425685f3c0338219b24d51131753ac79e199df34fc518524b74a12e7d669484e3716e6019c02a9d712fbca346a8de52986ab62b3c0cef7a5193241eaddc6e1493716a165d757f61134313a103e3c9dd47650d259560e2ca9e4e90fe6088fc2a2c280bfea72b910996bd5b5b76ba904d39ee58c7030771b80aa2c8fd9f1fc89b7d339231e87cc0621d41095c0880b3c1129de61cb00fb5b6bb1fe658154935e66be87fe9894c3ac3fc106c21ba42622328da9f1cae101bab3555fe84a62a93b6fa2707e4f13c6dd07c8eae538fe849613c5e5196e4b31077335a30495bccccbc18552109a4f2890fdd0d830d438cb8c7fbc7e6d8c71278f515fcdfe23f0d3d709084d90b521f05ba5947aecef6bdbcea0d26b267e6a828600b235f4d7466f9ace6a615ef51b30cfedd9ac96b12ba57b90b320c73f7d69ea41842ca29246d5cc2f2ea033974929cb3a9dbc4854723b91512f7f751ce5d6d93ee3ff2ef5c43acd8d28917ccf7b1785b658e452aa8f9c894b2bd1c09807fa8e70be2529f4af3ea604011f723a1039787e0a4da2dff5c87f18748c77d38edd3f2c2b290;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h9487612eb5b09e14fbde91907ab3e4cf8667b4c80cf95cfc51cea5c97591b6e3aeb23d9cee13205ab710048a4af85ae1dad4659f275361bc7ec7bf2a44234286e88a2be1463b53bd1aacc75373583a7cd2cbb0dc4621c4c5be1771aa698dc42abeeef5b7dd084a8892a4ab3311cb7aa76de10e123f2a2bc5ea1d7333a996cae3bd65a6029cc3c13e4277776fdb3d2d1049c265632afc7b52686672ccb9268dbc4c1f0897d7621cce779d7653e743f573c9528a6a1b729819fb01b0ed2af0503aa6d1633ab3e8a811f2704f6aba9b44beb586ec560f9faa4a7b227722f42b0a810d243f0f7c6aa8f228d392c63e4abb507031d02482b01f0965997c697a55a6156ebb15782196a9162f52a6886a01510bb770a9de2f65e9c2950a48c769bfe474554122d90268e8a376b19517c60078d62ad90e4741f504552f42f2e8170d89325ecf30b20a4ef1af15833288d96eee2ac07c4f4432bc9a7ab90dee1e6afbf76c123579480c3a45239b0b22e4746c1aae6f834b44e9dfb02944cd899b9597f53caf160c85d208dcb6cba69e58124da8017c6832cbcc2762e87a6e5e77a41ff3bd9a1a33922ee0eeb02595a8d17757fe45a5c4eb63688005d294436a3347f24ff5182c70eb8dd2746950d99b09181af0b121b57eb5f2e95039c6998b5c91e4815d2fe5b11f417bdac74300ffe217495a9a4d05107d3f65009c3ae3fdccf4b0bb33ae04221575b4782409c6e21e0630ef94a573f23927498d2dcd6b1b733f0edfd718f03d1f11d54d3192f00eb9416df76ba5a1e98a10cd2c025fc596a233128fb9d0dcacf52e50d64eef7530a8970c8a2456fd7dbe6814efa44d0f0fdbe2080a982ace73bd4dad3e6fde614a53184d128d1b436b1c1fb92e7ed4f7f59c3d30855bcadb31586ad5e54add2581a8e95bf9ee30ea94d5f6413e62252e746792b7340199a70cf0bd417610060e4e81ad055d6da58d2be22a245a265a513c002290f794ead54e5ddca1720cd476e7c842a15028abf6f7231bb075222edd1c8d26c7858122e3cba6eb69cfb3769b8f8a97d981fb40b75f5bac3c64226d91cf72a7ee49419bd59d7f195fd109f18792fae0fdd95b811b2b510b5764874b53d47644925293f19cdeaf6477eda522dcfaacb59fd971b10ec61c0d45a2813920b9e8e9db4f8d9caf88d02b5176f84981e8a0f2f2cc9e0398ca24a3d5ae192fc80f47b963c035fb8ecdae9d4217a77d6a009373174577f2268d0e0cadd4c46df06d4d92c4f7d7ebb3a9d92f8a4c945e55f0c059015af74597e6fb2ede27538915b8b950dfdf46aa54c740dddd3fb9b1c4f26fa38a5fdd28e1a96bbf6fd321e5fc9338e51e9a0ff5616937d9e3b7d27343da0f0e605cbf5638de752e2a7927e813419daf4c57c28d26295c9044adc22230905f4b6fb4d933cb3e28d14781ce3b4fcfa6b137ff1435a6e375e2bdde592419ac7f55fcab68f40620cc32e30b59bad78b26f47755a49b98bc59ff5e71083a3ddbf1ffe75dddae874270f4378cfb60b45fd2e17473dfe628c07c38317eaa8e926cfbe2fcfd993fa73c6491687549ba1567671ea4f8d57d2088aa4519aacd9e400f4981d01329f9c1ad10dcf77a1b6fc1357b0925c1a1fe4689a642dd2090fddb1f43f1a24e76558479687693bbe57259a969f923047e83a3e50a5d1cd5798570d356fe999ae9fc0e69ff8e7685127cf63eb2c096473036c044582dbc29261535baf3d8e8a0a857c0e5e47f982c6b6969246842701947291fb741ac929f10dddcaff069dd5919276d009a2660f6dd112e67f8d8345d8b4e7638e2bc5b8536ad8c9fd37bf01b32;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h910e6c281f234f45cc11ce644a5f8e00f7d8127dff3c5fdc464e01361ff87a68b35bb6fbba6ea26b473a6d25fb298ab6dd90150b63b6c84c2c2cb786819e0a37cf793f4e19b499e599ddbc1d817ea8517d09a9eab58d243a7c8087b718fdedf186254aa7d07ee7470c1679af5c4e2cd68b8d9f4cc20af7949a3ae075982a5b9c0835bfb6445e62f396c03e201eec1f0926a34669038fcfa05a66e913a761659be26b94a57aba5a2e0665c577d9c8a3e968f3051691cbafb0247186fd12a0458763c3b18232e5f0bc654118f7fe92a8d8ce7d6e3f2fb0b161c3cc78d1993d6d592a6d6904d156336634c8c3ee339c9c5cb480c307cf6b00008a47a5586d10c906395c52c0bcedc35300069a31d3728683fd289c9dfb8e6a2e9c71f1f1c0bba2c93050e3427af1b26bcb1fe11272afd83dddc996f29fa481b7c5087773bc47a86b3a03f68afb911c2324dbaa5b3eabdd60ee9c2492e65ff373b216452e7cf7859333ab9f616a1561e183cf52ea9fd1b14c0727ed3ef1ff7ad06542d3cef1fb43e8ba4812b6b5e800671f6e45db3698ef92c85c374199bd3f18da51a9b8a43eb811d6f4af8c895a959754543bfe9eaa902c20954c68a30898c90d7cb268cfe288657d5fec1d32b3d0215fefc7bfd6e7f48f70fd58f7f7eb7a57587aff1024fba0f94767759816863b080a4500e8817050618865d4cc48828de2b085082b7af5da04968d3856cb2ce18d745ee1a4e8d0be030ef45a0a3580272b3b397999de742084a04363f1bf5175898c272259b03116d6640fa92ca477c54e49ed6024d8d513ba81d626cd7d37d327f2c896f2705e301b6308e08a23a31c9b97f3cad5c41c2abf2e8261539b91ae97a036cfa675565393ad8656f2e8e2771e06ee05ab186ac120015d941f72ddb16d4158651ce7035e9f4ee8035d33351bb8c2dd585c23017562cde8cde8f8c6e08fda479b24e6c6939bb621a350505d3729838d3f0a87a03a25dd49e666fe5757952bf3ef38dfe758e94d7a70c1af0ef16b3ed8095079700b06a3671ce022ddac5a9cb61b9fd794590ad030197710fa8a053a21201c49507a5f94214f420bdc8b6cd0d09eb547e3cc4a16a3f62c5e83fc0c12ad018fa21978648ebbe58bf6afb633e0640936570f399e552612a3171fab85888975eea511427c641f428ce6c3dfc05454b6c676792309cd8bdb4bded2b28edb640b158b8fc1e6dfc746282fe819796dc76b532a1872022d5a08fd6ebcd7aae90591d8a2346c10051f3678ddfc2d2da3d3d9702659ed31398930c180241e5ebb3a35971fddac32986dcd8b1d9b9e7ef5a9b4d1c69e19d5144ee62ade78e336bdccc3893062bdeee8e8bab66ad7ec72597a6b1465dc58643f9cbd118eee98788bfa715b9a62ed2971fc416514fb209fdb7a0000f368f4e500ffa0005030acb738a2ff3d99520cc860c4b0726190a22c71ce76a4af8fb5db15e85ddabdcde7dbd643d2ee2f9361fdbcbef9a40fb1933490e9d6c8b7cd047edaa710cce9236c2edc0d26591faa80be6ae8d427df4f4efffb6e8d655e36e0863702b157bb84f979e92991717d9ef53e9f7acb0227579138368603f83169feab6dc0b70d75306c041a62c0ca88b75bd15ea2a7454036df9bcdd0493ea18e0e7200a92792cb2e9437aec7f3fffcf230335280db1e8cfe966091a497b9c27a12f3061fd513007262571dade683c1b18f38f8679d6a129ee46545462490f9fd28ee1f57d750ce0961c4e5c1a2b6d1a1919473189c04156cb19e4cb418fcd014b6fb0c7abe8f9fffa7aca0bc7146533690f08c205aafd1edc238d82fff4844c702ce;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hc8248dc3ac4d298a89c7e1880e37a454e8a10d31e5efb5270dac5f92efddd6ca83cbbb3214d9e931f15ef7a69444884549ddc2ef754cefcdeec061c4507397f0a82dbf2f4ad3c1b00ff26adc6e66d7618e257a0d2c4dec1a6d1cb7fd5d98530e649774a47f3f872980ce274b1afb5371a58f2aff18260318ab44d864c38456f0d461b140de691623c3827c7a49a28681dac77cc27367f3e8aab722036e6a50f0de0cd6fede5633b1c14aa49066605c7be4c6aeeb42ecf6f191542888f06d2cd0d8fd30da075772ef40c22da4d3763d8c3ff136dc7a25716410282680c8e849daf7fdd8db871bcf1c3bae9d3b8575c68056c236aae7b0d6f8e90e1c6e3b8183ff7110b4f690049d05cf9655d28ce7542e419f9f21f41d90cb1e4dc7df4eba141ca2c6fc70313997ad920d833bc62a99b45846ef29a92475b7ed3de843f35448bbda4f7e04ab7e8d35bc82ca9e86307fa17928fc7d36e4fad66bf8049f1f7701e40dd2e4f7a0eaefc507c7ed2622fc857092dc07c6c965ac47ab270c6e3991eb4151a494ce04813ef0ba37bd2b24344f4df9944e105fde96b455109ead5eeb3cd84c2354f026e744b35c44824d2e917494143f98333ecf8d72871e86991e514911ae77c93abbaa049df55d66e7480ab761b4d66840cc3230919e8d0ad8b87a735c55805d588716fb16aadd48bc667d896780b2f6d55b84a275306a9635191883f85591232f39bc6a8f9bf45a9b6fde27991217f8d80ba472c8228cd2aaac8e54a0d558b9a5701d4a5cfd8749534f13817de109b2623944e4dca82343b9bba2ff0f027739fda5b289beae874c089fdbea49956ac5f15af76b99a9c38874ed374d5edafa5d37d86e0cfee9dfea6eb06b4ae3008d59527196c52957395dac0aee70daac39a6312da0b037f56e0cc6335840a6a0ff47ad7d864c358c35ea0b19895f173096b7d9142d23853ef3095da0522d6b5eee0b4ac39dd9c2d89b4cdc844fc644181272a5cd7e1e69804bc59503255f099299850063e12417a0cf98c965c2c13b00fc995c3f8ba815ee44c8d1e289bbb145f2c15a20435d98c006512aa3413bc8f2160b62a668f4d3dd3d7f74dc025e586ed4a5153dd25f0886cf96f39c53bf638b329c777cbeeb32021d7c67ac101eb1081dc77e179b1b033b7a1f9a35ab7347d9521a4d525fbd5eba9a17f47aa8b361097b50ee2a0b0ba2a0289f8491f84ca13b67a901024646dd4e746b014aa9440f52887dbd5cea61c3a7bda3c129d875ff886574f3cd943c0dd03145e20b7545b65ce13dd733d2d50e8fc685cd38e0649c5e87c41e806bd19a1fc57f647c571b3c1594b323d3f3c346af193e316af1a30e921eacaeb783d23ce15325d30ac61374401b6ab426497a3a7c652708e179352efbfc63e138e002d8f00eb38ab66ad47acd2eaadbf951f6787ae61df8d87b303eafa5d5c283f717b93d0bd7bbd5e8bb0a5a520370ba9e2377987fb5ee5539a752f63342d37d13d34c5dcfe8458f376e84556e10bb7e2d9647aecd36716b80d5aa1f292835a5801e687a7e00aaba5366de0d9ff68aa92ec8bb4db2763bb11f5b0204294daacf7abb7eb9c752ed5d2614e3d03a130e9c3330565e2695702fcd0f2773673cb401602b1377accfbda8c8367ff280a48ea688432f5c5689cad1e1ea35a1fc5d69fa3e105274fc4b12e0f4b2dece8246156a8164927bb6e75df66d4b5fa279331b5679a2d722e5a4c5de9c37efb005c79eff7f01647c7e9bd86085d9e257c4c72eb40559814fca2e960f36679557f8d40f0a68c7444c562c319d74fd1ce86ba7aa80c236db88d650d888727776;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h484fd1416568f5c348764db7825c9d0b346ff041787599ccb30c69df8d857ae4539b4628da46f8f821ff572c06e7bacb9ca13f91791f565d6b5d73ab9fbe7d9dbf1c17740ce138ac5a5ad6293fd57ae7b686c8cc9c189b721f20e31db637d23c889553474d547dcb527792c39bfb791da30a6174e987db6186f3a348ed83db360c09e20ea7fc91340a14b1ac98f5cfd0d743de461dfd8f31a19875a5a65c5727005fbbd11f636f83a58cea296a99999bbcc02e3c7b855d9b7a941a02622cbf4dce3ff5b70d7abbf14590a2870e7aeca989b69a6e1b1040ba3cbe088ee69d270be8bb8b02a0498b7d6e2e346d5f39d460228840266ad95ac43c92470599b4b3c7edd9f6187b42d6bc9e5359eab2a926c9a0aa515bfd65ddbe6884ec5ed07e6ba10065801c750a9bff4f1794e3e1c6e2f37c5f6027cf9f6be15821020c627831af2acccb6aa45f1d41e2977a309401b2089979218959f99e79b9db694d0e78a75fe307997c4b09c445f8d74beed943c6a09c1dbaea8d63886c0c997edd595f58eb796e5dd359c5968ac39ef35a9b6909a83708771961034b36e5607b4b78f46c22309ee2f6ddfa943a9e467446ec53c6f8444f1df9ee1072a41b51b0b1c945b907b987eeb8bd42fe8b8f3b5217962d5e8ea03f82ef2008012f33b8ac2348c312a7c2c5bf79f4b12dc4fe909db3b1820b3fa797177bb27732d9f610e57f6b89dba10e12f3e33e4f99f6a5f5da124ca9a19c79f8675da6f8602422facfd6bade00ce7c7f1a893a1e6b914d10929e252197d64ce184f865462279763b95e55f4cea47cb7c615a57a684b010e9cdcc89d8a9bfd90dbaa24a2d9720fe55e23cac227ccfff65c9b00c368ca935bac72cb7ff47c34e02344aa5668fcdf2a8ff7e7910119d00d058d33b41c7d683e8ab1f30e2fd937c8aba8fea53c8bd98e81b687cc5d96c2897e13dafc96927357dca570aaad0dcc36e1c8fda854e79fbbe0fdcfb8744a67e4d39cf6f6f607c9576d97c96c190c1c6b79e7aded3b87f5a22bcb3291c82b2dcc7517c15e15475fa20d5efaff7bc98f44c17dd11182c14d0e3bc58c414924d0a5a90fd3e7f9e1a802ecfe0a2d171b45c481fe5f85450de9a0c59ae23fc01b47341a49909b0bf0d67d185c9a57b2c6287ebab55a9de89f6b347b8637c1a76be14445e9276a66910bd67f5ba1c86cca940123a85484bb4fa9fd30f2ffd92da0aa5585d4af5ca699561b6d3cccb83a13ddc939e0ac4c8361b3ab21ab669a419f64b1d8d36f782e47ae4841e5d3b476882fefe3cefde9e247f3115c9aca457f9fcf925d84bde101271488221545d098e761fdf7aa07a8afb8a91965984aea8c77aa5520e4c336097f8bd0c3dee098480415e6e733261e625248bd97f2d5b4bf3b0351ad34d7dbf523fe7655bb6c4b84bbe175b515af903c25748bb62a84b9f0b14af67a22c336409818e58e945a7591bf4d6836a1e684ae7ac0a1d83c368d3f3289bc497079995780c94be97d3e0b4df24231c50a6a62c52371da607c6858f5da417ee3a116eb6903f03156ac176394872e4aafb58f244b546aa1ce6792cf246cc9b64ea52b2ad05643e7020b73da30dc510690626ae7fc67850bad4e5580f5752cdf671c205c31b650686d8bbc653b26bb9ea4bc185b42226111dd6932697ae8fd118ac40df5b6ed18ac942619dfc1196728f8930c1d6fabf7e0e8a7aefbf648bfcdec9b2b1939dc1c482cc814e72e9ba4dacc3b10f5ed1fbf859c7c51a3ac2b4c12d50ed33e33824e0421c95d17f72214d802af84760c74cf89db60e84ab740c09f262daa3278b792de406af3473e972;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h11e47a2a3e08aed67bf135c173142fe6bc1f60c67b04e5f2e82a742b4ddad7719f2f50817eb218174143b6028c58e75ceb1b5ae06ac28e527516b34e7bb37bbe73b4dbc83a0c1b072a5485033f3de0f2c3a13cdd5949635d98b7708d9fe8f5042bd03c4ea9d970dc19922b62f76f5bf341df013208369e9449e74f81c14ed4d8bc3beef0f925736d2bfbd7a799d72bc755ee3309e64fb2ab9e73b806647f09f29567c295e4b2d3574a7a072cfcb95c237a83fc6e9c97beaeb8eea60be9e6c6a577da8a05cbd0b15d1d5c391157f83d56195a526a13df5fe3299511aaa8c310d34103a4f15b86d883ae2e2365e96e9055dbe3150e4b14086d891aa908507fbdac20829d5b8f0f6237a29562fa146a6cac8a6638b548c33f6d2c610cda310907a08563bba347953b9239fc6844cf02f8197a44c3f1c643c435acbe03b854caf6ca45e06f22fa4feaa10356fff2f1b62529951071323e73af6bcf79f55398e49b9554a09fcfac62ab38350a42e236aec23c934847fd1ea4da67b7e649e44e0487b4e2e451187c37519a71202998eb3a018ab1991c664a2e49a405ea39cfe2832e2e56f12ae400891589596c42e3e595a41c68e53850bfe6cd706e94631f70fc2d821e67b6ea1a7c333c9e70cb5ca2fa16a8e2453ffaa29f01ecb64d1df4d28b90b39389c293ec3876d69684f5e475231dd7939a63c7f2a528b608eca21df6ac1d4beebf482284b59776843b7b4c70a1e9015de3238ec9228b360dc55ac2fb5047b334bbeff53204912b5c7c75fb8d539368f1b0467e9f5b0f7f35bad46b1ac97d6533a418ddbdc9b69191bd07234f891bff7f6d3d4fae03f536aa2da872208443606246ae73b09eb9816ba294bdabd679fd8cbcfd4a408f62e6e35e87ceb6a6cd6b72484c1de66682cf197c8f771adb0182498dff452dca212852e894a6ac7ecab7bbfe0c4419041b7289e991e88e017c3cd96887d3bfb2450dd60eb3d7c44c93f8e4345e5f6f11394af8fca168a7ff1ed553d68edb1e2dc3fbe9be34a5cd17327b07345d54cfa121094f2654b3306c7e31ff09ac47d4a1fbe738e0c9c60c252cfc0ffbb7534a5412f59c3a74af55d8d23259a5653a3a029c3c79ede676fa55bac1b82d5f1729fe02ff66cc00eb79a79d3ac3f3b5db81adecab26366c6a985d1054902fb9bb2b888173dffc27b8bf2c4f604d0ad4273897fb426e13a4e43bf616e9869310f8c5864954ab8ee410c4abe648be7c4d405ecc261723613aeec4f921620e9ec13191350bfe6a3ffa3f7e63102b4c416439b172896870a2afa73b945798ccdfebfff543dc3a2d925ef12a6b9e0994705634974e0a25f3d14de1e061f017f423c777667efb0e67f7d3c131a30d0666f967cc74aaea7088808357baddced6e9c5ac6dc2a77fda0978b831adcabbeaca8e56f7e7a5e3a5f79bfb1128be2aeef674349515ddc9f7ceccf453ad6c9e6d28d0658e50b4e95c6265fab680ec91bac5b2ec5b491301c5dea6539d3bd08c131d2a70af76883c284e3bcbc879714374bae127312c33d7ffa3e7a219dacd6e3792822123825c3265c59b9bc1da71e4c68b4d1bb591c08ad9a807e48658f0a37c41f93f9f0a32d467e00c98a26ad0c5839dd7bbced51782f581f23553b786f8047aed8270e42f2e8872c447a26a7add5961db533f8cefff65f165f8d2b6dffffb5ba557db662fde6b4c48d6e0eb36acaa6db45e884df2a85c14da2764a8600db6e5108e8a62af7411c25af1b1675863e89d1c6709ceeb5c64765d2f83612ffd37067332c301f89d7f067542d50e35a4e29dbeb82cc1681a9fbd0556d33f21086b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h83c5984b4c9842fbb76702fe664c790bd27c5f0f8ec019703ccceb3f7b43b1476a6a3ad196d20b1bb47c97bce4c0dc3b59abf7d92ffc09118311ea1917912dc1c45b0bf1491c784f95b339c7e8787fad4183a26562ad8eb8da344c204366e616616d134519554b5ca4eefd6c659f208b564195b8e374bd7d5092a0d53fa5d0366e2d11bd6bcabbee06797adb260afdd9a26b96df52b3a0044f0dc0ab4b4527579d78cd6c73c2434ceb388194a7fd14b6a77a81e1ad9aab4337ff7e79448bd7b7d0cacf0a8daffcf7dd1eee4b4fbe70b8c773b96c8591f783e93380c956e80508fde604a219e33e9dce22d5a0754f7b884bb352d95938f33bd96b25bb7bdc5ed6b576dde10adb6d0b441aa164b123e0bc0666d2f16f62822e0a81f6f4d178ab67fefa783fcd6200daa2793dac1af66e31257aedb067db6c0bd05996b88f4e4d13e7b5ea4620a94393c4a45dc81f8ed906bc6c2b5c4e1b6da66c312ea3bbe81b450cb0eb3fcbac8d4b0e94de9fd090a0ba3040ebd6fa820a056de3bff652ee0dc09539afcd82764b9172abf5efef0b7bd492f9419d3776b4eda4a1fe6169b512c6e5a90f8123cb47f7ef9ae13d2d57ed0b3a3ef23f3ea66fe9423bfb2cb08cbba3340e93820492ab2bcc1f634bf30ab4d88b8947f78935f6147d84d72cd2db0346a7a1e7d2c34dd5596e4f723e23c6139fc3ab1418743d57b93b25d4b52b536aa947b3b82ff5b2dc2e080cdf325b6bed9fcd303bfed19690b569db6ebb3305ec45e4f61f7ef9e6cce64faa640d76ed03ec1790f9329898a987099e3c6b1c1a73fd08f1e7daa73b9434afc9ecc3793fff4bc0ab6b51dc5abe3c58d9f12c1de3e6a32a2d8f66e702a6d77030ed9536f15764aab0d0305ffd3d869f7d25bbe635a23dd09f2a6d562d52c514e46e7754cdb38cc24f0dc7f329b458c8a1c2cbc0aba697a7407b8646e6e6aeee5d6fefad8dbcdfc40cbe9d82aea74014aacdee8850dcc8f9e09cfa1ef242d0f9003a39c5dd2631f3deed028a069b2d4170fc341215125e1657b552732a60c5689116267179a9cd4dd1f9d75e51c4b1cc7eb56c9d68e1028b6f9792b13ef253d6a38a672d552107806674aaad2366c12c314fb77b1646c0ad8e9bba081fb599fdf18cc751355281d02094a3191b182651b190fd14edb0d0a93fc5d051135c242e71369cb4969ae0378128e6ac891947cc078698a555f1b00118e5c12150707591abc3bfb2ed1096d6adb925aa71d07f25e8a2db57ee185fe1b4bfee04a1771ebe8cfd02d5b0ba1a65d965c42be9c9c442443eb00e14766c4c358e77612f87f5e41883014a54e23ea9937e9c4b3a57435e71684a9c67cff9500f267257ceee89fe9c00a45ee7641d8f36e67b235ff813a32996f0103692e57951f779fc197acaa4f1dbd15781c6b730a58a31b99133d216db5c3af8e3cc1c0c3a14b204345b7b466c6469038c4834c651f7065817558b78b1a7d9fa750ae592159e0d3e985df7a9ac4ab8ceb6ac5b257bbf5c06a65e039e82df39b2aaa916e9f5028efbd6663393fe3cd5257e64140022b8bed60c8a5e7aa49dcf00294f3c4cd0c6351f344a79e08a61cb7495967e960fe11cae1628068872f5419d0f2bd34e9d124f2602b7d7112d016864e33c234df2d7a9b58d5b106b48af0cf58ebbaf07d4a926a267a55ac4863ad77f6ca567634120c1dea1d5b0af55ac452904bb3835537998461c7c3b416f025a7360f1cc0b5602fc20d9c281447a5e6d1d39ab7e49ff022c9c734fade98f0a9e491f93a4466fa26b48893804ce071828c352aa24f374aac7bded3604b33d754c864d96ea;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2ab0476a1c2231f221200d00a2af7cee27282241c9d86ac6a9c7a458ac4bac5a85247c298d22c7f44fe782b6442ec46c2aad137f013e6c6a84227b8b3be0645ac8c47a5e4b232efff328cc6f13621e1ab49bb7036e9da5c359810e97c04feb5992b6c6b980dd3a8a960504bc7f98298c8c7b171327b55c09df998b3d2d3f2aed066e1efe3c8a6bb47c437bc80d4a105caa4cb3b7f7a5d8c10fb37bbde9a9f70ab285f69c7bf0b50c047af79520cbdd50adebb90f6223c796caea4e89fe6cd4d8a0f5e9debef14e072451abcdfd662c8faca9532483a524d3164bd0b9c50f94c8d4fb7743f4a3e35943267ab8b5a8414baabfb5ab9fead74a1716946dc070fd614c6e407ed9efddb9b08b5010c031f0f280b8442efc0a03cee966d84ca1d7514495684779c6d98b481e60cd2b74c500d42b5ff8beaeabf66ef81893c0477d060615705d4a0c78121133c1dc9ebdc6164d2ac59f2bbd329490fbe80e2bf4e22cc07221c2094577ae86da19e21b67691e1db2420e93a819fb1e94db83b584fb0987c344fc3873a7ce426f1089e6dfb2080a0d63b4f1cb03bc0ed8675e5dec5a23f976202fae14dc2b9c1bd22dda14f23485df8404d419bad1cfb48c407264e94dbecd0dcbf11d7b80bd2f937cd853f40a6e05d6dca9053d578b0c3ac999a44f19891e202e578fdd398c32529e7dea00727dd2639643ccb259eb4cac4aa75bb2299deafd0d882f9f281709940483b301b6178a4cbbee97ea44af8eea730e06250ee0a846e6aa080f641980609b88bd0a36f7de76dad1b9e61e6d61d8176b13bf1687106a930f62808c6e0c9e61b32ac8bd7fe0d25876f2af4b59aaedb096852d1db6d6c43b5770e4704bc23c1a3f47ac583d61de31f9a3fa4ae1ca570cd46420faffb179bee0c0e1ec278e9d73777251373e072bf93b92461d0df806376519d4ca70037caf6604e88996fda23383e6416eb0486340b70f84b6e9dbe307c65f9d795152ea4d83ffcc689b8e34373054bae5e219242dbc3c471f6a19301d4497758648e170901b48a481bc19c1384031c002b650732158caf40a92564432b27fba240b57dae889e47fbd51fde0b95a2c263884a8a571a94542f2450cb6f766a7af74e19863b258da0e6f91735b0126bfcc356729fc89377b7ff0e8170083d909f2c49e09f45ef3d9ab6d0bf31471476fd618757afbd9010d0db379c7d2fb46aeeddc498b95e7707b83af5d0732c663a71762a04a7214d6751877b1a2710aa0baf45f20b07c061160dcab0a6d4ee6b7f0bcbec6f647232fdb971c016b79e4a1edc891e0c6077f418e0df857a050084df0b67e30ba382d1263373d889e3b112eb4d150578302e74ff86fdbc7cbd3502526295def2c911204c49852213fd6e60a194f0ee86a6df215f9b56b831f707d44b0fab357b51a5d3f1e53a6e70fb31012050a48e1bc4a51ec7493b5b342b8b58d38abe9669642e7496a2dec582faf3800afceac40a7d9994fd4bb5f3a6ba06b91e90ad8888ef8ad2900a94bf3410541906ce869028687ad63f635faee6e8bddea6848e171644f99f7e9ac275c3c97dcfcfb9e55641e3f5c5e17373510c39088328659493bce6eabd20f3c06d87a6e2f68986079db434af9c9296800567a61e8ce023074f440594a603e5088e5c5fb88193561fecfd56fd5f3711dc5ffd202e1273d8bd15a20c76a8cb8b80297f416117cce0f4b244f0036cb909d18c39bcd0c3b5fe1bd5d9dfd3f3b9cc1d38722db78a72797194d0193c0ac6f2459fcfb297721d20f30b139f5b55f66ffc572635f4a4e8d98fbfb4cfc829645c56c8811e7c83da1bd00b4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h7b63c5a3e0d672cf7e004982107b1a69ff258b43296ae38ae122d45b82854cc3b8a7031a77e1464105bac9b6b1d419cec9d6f6dea37bc08d624eca3b19d7a797e8bc6fc5544dac19724186e8957c9e911ccb6fef9f6c54072218646ab378190684f5f718e4de3b93af60815e9dc60e02928ba4bf9e45cf1088bc2f1723256cda0ee46a3cdbedaf519c22d4cd2185a1791d6e12cbee8766a6c80cdbc26cecff9a55606e1cca2a2d1c58bb4c4b11248cb029028a5995b56fe6bc3311d766c584efc737cdb452102912b7e8c2ad4e1bf4d7aac8c17e3029e5814fee773e310f9b18bc73ef82c8580f6325750eafcb957b4d6e2e25454f3245ce522566f7e78b06530ca6b61785940db110c22fb4d241ca287054c0ebef83c1b64ccf653415ea1bf62c9cbc7d9b54c3ca5e458c2859f2dc1e66c5f8cad12d05edf09db46b4a4e161a5c019dc4e3cb771e6f38c97606cdf8ee25de229e86bbc9fa2f9d558e9ee33ec90f52dcfb396a47340ecb19afde2d900f14bb51db86ab4920c5abed4d900722f8e5380d1fefd9505c19d1b283b4c09b6158e19cd08fecee1e26a3de0207a7b407a3157c80f8405acec2136b3baf55a9c5bcf48206e07e8027bdebbd151447abe27b72b83bb39fb0fc95c13be870cc42b9fb0e31ba5603c17a65632d794fcaa6acc6fab5e76eb8a3bfdeebaf5815dc32d4a55f89d4c571f513ab3713b9a4594a1cfff2188cf969f04b1480007da62d4cffe165c922b1fb312299a9280645c3cc212133121cb40980ce9597c5fbcd28d86d9afed24848b0e23bb47c675a343ebb2167080d493bf463946eeaac7b1b107053c349a28b41246b105d8fb3e18feeb34bcd374349d00dcda99c1903ab6c4194b2a1cab4219b9ac952dccbb16eb56a55429ea43b8bd086a609c0a24dea6a9623b5de6badc5014739d41bb21b079eb885e3dfe49adc1b2a0ba1630a13491033788ae3d44d3c803d7db6d0bd38997527fd7d4a0a95fa35a9f1ec9c8ec68af55e39d0d753b38e3c16388108309a2e82f45427f731a6c46cf06110144d0e1cb16bb58ade026a481c9ec46a4f4570da48c9a5f18e13138d566cb97dcb33dc775d65349b2cd7ccaacb03673aa216f429b11c02c834826cb853b5139b144ecf679d8951fabde120a86b7cd88365232e59b0b9ff7bea3b00582477215cf0fcc424fa1f36e269da4c57104fbdd4d92346ea81b978628345738a4073fbcce294f68ca64109ba60f25602c4add074a602aeb7d12ede02b89afcc5fe4fdb1562715ddc72bbe4c6543269a388411d456896cb07c0b0aeda7a099788516d5f44d8f8fd2e88ec7f25171a826d974f70291b7611b4d63f6d6c5a978beb1590d2e185d7598487cd5d65fa8e093052d11bddfb987a0ec54f21cbe128f7d1dcf18e0d66a4cecd00bd21285ff140bc71abe86cf035aae5ce1f4b84d65a82633d0afc7cda4b366449e3167109addaa0b9c32b8b0e5d62857bc36a3670966b9b54038be48cb9281a0efde7c1ce7d2cf5a188b034d7961f29e0b98b9abe90c46058fbc964618e4c3c378cf4a649d323c4e80699c1fc974393b3f4932264e92edf7a7cb1c1120919531880fc2ed85e843ce3dda9a20f817c1c35a132de523fba76688c42c52542d3c8117af3b845131a54ac57d8bd3402e03d755e281ee2afcef8f811401a27619b31b317de6311df23704bf501903b638a454594859b0b4dbeff5db4965a4c56f4113d5a823d8e335777934f66e0260307f3643d133916a320eb2a1aa0059268769ea142db68fa5fa2f643fa47db231111ed7a07abd8243cf1975ee1af88dd25e61ac748bff4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h7148d957df138a437f97af635bc8ea7c8519eab0966686d1296db2190e32ba3f6c028b89da08e8d0102d0fd086ce395d6258282ef050ff1ead9036f2b5623e622e913c0ca924e8c3265a762f293d0636b2d875d739cb2ca7605499bee2b13077fa199a8be285664152c61cec79af8c6fbea3453e9a235e024867339c0ce83bd4b072fc455065cb2cfeb8643f0e3deb2ea27a2a8b6825882ed2eb36d4b1306bbbe36608e790c4509ce1f4fc02c1e8cb3663a6e75281a2d8c623c7295298bdcd98eab1d5df3b9aad83118271c7dded2796c8c9549daa6d3657b8c37829357d94491cc9ac134c41033917285e1ab2dd70629e8b860854821feee005d3b9e3a2d72333f11bdb1031079c165fdc196f6088b52f41e010d19162e13ca0ba77fb3d4b7877559304b88f6dff52b74139818592f14859006cde1973a9152817d83709ff92fadfb48a8307d7a196cfd63853356384f1a2fffaf462f6c0a02bff26ff6c486ae4d643b9e5af06d91713d0bb7b482622097c03933e12d09b2d7d999a7ea49608e6ce2a0740e781ef3f99d10ce2226ba3a3ac4b5f8e15546ba96449617a6d363f9ff4540cc9da79770ba2253eb8065c33f2d79d2a1fda16b3acb2be19964d638d4840e85658986ea57d793e48d0d8b775753c0c1a7f6d4b1b7f8170579a9d64ba4520d128494221404c2e5d32da6e4a0bd2637f8b6a26726b8ca1c5460bebaca6f5eec6a40b85c3d0322270baa8bca3161f2eeb9bd6afc0a4422484cc54c7e9a5a241e2c1c2ac96e2733decc9a4eae6758059340b7d78613944969ab5d446b13d4d1362b4df981f7a5fec574f95f08c8c93c7af12a4254a256d681ce1a443d07fd2d3a19bf67ae703323cafe9007bcb30ff9900a56eb9bdbcd476063189b490d8bd5518c1705326ff60a652e3c069765348118e0d05f81347e1e97057e50be4b2f32e828fef8e92e82fcb2d9c61d4d3a04ac327a7ac8f20422c3f359b9f0be38cd2b1aed0f69c0831b127f0fabc458b47d314ccc4b9edee7e6a67601b23384094b3a5664f97c546a9dd17c451a48384919443218becd0d591797662b47e374276dba04648781890041766a3838561516e212104a02a647734f54e816244b3a9174b49dffc2f04be7906bccf314b24e382297af71c3e6a8a942dbf3a7ba25c0d5c7d1c39d58042162ea552ce70e8c31681449e0335e322f55a540af9d1762cd79ae7dded485fb8d9e1f41328a69b2548ee8caabd2603dba98dc9e5ca7cb709244de73314724a75ee3ba76835e65567d421b1ce946e88a960ef02230cf025bad0df106605e7f7e852ae3f024e61190f710142c825dc90c8895488adb71cfc8fb462fe96a17db88e049d013a93bcdd2bfda9aca609763f5853562e41453b4742ac651ae35fc83d4cd6b452efcc785770f8f15442056316f258a5c19cf5001dd19f5627bb23c0fe2650275b81ae423b270b81e9abdf426daa06164e2a58d2d7f1bdfeb5270609b18ae8369a59988b3f7220b0ebb8b68b9df92b99945e16e54de05f18f62fb4379f13eecf85432eb5a543d55832a2eb3fd857fe974f0b77254988f4d337ed39a0804775bdaed109e45ca5bab38f542c1842d8667e75e6e217f6b45e85390f82e129f67c8b84afcb72361ba03506668a612526bb3e21055b724930053d34e3f571bca2fd0fb17dad92c824c39eeea3bfe4317c89e31038dbe654ca2e1c35a25922426e7e6247918b7abb412a706fc26ec58a88432c32c5e786d05d24fdc577f3fd63fdd1833407217bf3a7123d2423c327a19333ac32fe64bd69d64b91c51e89887eb785dea4e0929908703ece;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h9b9a549f5413909c49175d215ded819b3c19ac2770bdcc9078d7a86cb56f4795f561864ae8d466d2855a278e2bbe15403a94bd56cbd1b88e094ce86289be50bb92a5e02711c4d79036fbd9e3b51643f7e718a2eff9bd0651be2d9cac21e9c0798976c0a2186b54b9d3959aba84c6a23bea30b8d516b31715275703cbf7d63cf000cdb43aeb4c49d80c86744ad7b97ccb3ab58e50d679d3da8a14809fee2e36a77b48ffbb837c948174229837324c9e478bf3c2ffbdebe86b335d1dff36bcb14f2d2d18d8f7ba8d0c79e789e30256bd1738e3b20b47cc72d9fb4c14de2fef8fc63b9da175fddda7d9dd5f39a5e15c807bfd12513efe6c3c80f8816ea52d215ebbffe99c001616fc7847724281a07faad80198e426b52aaf974fd935940f3dc63fe002d1b1ae17dee5487e566a677e407df5a545818d278eceab3bd7ad530c7fd5c42644f477f96b06299a7e1494f22eda9e03be8a5f640e396d0843105d66cb266fbb20ec9f4fb021ea4fe66499780bc0396a57e2af56d0e77e60212081996f01060d1fa4b01f562014e066ea855647fa3586bbe51f79a6b759c96b38969141014c5d2e8d33a75a4013ef6f5d3ff4f907c3add8da94287706c0a9aef3f2574b7d446ea9c1344a8eadadb2f60d81331117f05ab654deada202f4bdf21d54de58270504a1661f94e779d8bf59381adc6cf393639b0d8ea93d8ac2836cec630f34aada984096e4276c0f69c21b953903682cebee15ea90ea77068f2287f3ec199c5da9fb15f0956bf00bd31653712836b2b6a07ee2ce2dfb97a126c25eec2c3fa8e790e90fa5cb51c54f8afb4ba178f997447ccdeb94d045b421406103556ef022620cb305c1ad86299cc83d7b7177c71321d812aed65b5f2bbcddfc09d8aa644332382a8e4872a9633f01e973d568c3c9cb29c6a70bc776c6842dc3c6a8a30bc20248497b896884e14cf1f08b3e5ea127fef6440185b2c7d7f33cee71b5053669da60d920319217f02889155ff8243443419dd55195e943fa4b2ab0bfd37719e99c19e1d67ea625b12a3d24e72dc73e1f7cdd63a5f0612e273f5d5916ad372fc02a8ed285fc77729a74c7515a516b7219d78ee9e31df8b2bec3cc97f8bb8a20a15c367a98603036dbca4ecf3756349b1bb173b895680697037c2263103a86f12d88e2545baa39c3d4198318da722019acd13b8df14c333c5050eed9abc7922e5390bf8bdf6e1541298444e7cf718ac51b6868fa34350778561db79425eaf7a26d8e0ef1b1c857b135ad453c2679fb0c7d93be1e881483c7c38ee1109f48717cb4b26fe4971e31f10cd9763f95f4f47765b10f7bda5b6d11f4dfe3654db0081c44a0b4a84bb9936fd5eb4cc0ea1f62014e8e75544c497879de349368ac0df7d7bc7d57c39e86e50d277d7dbd80b729c36261b0c413b4bcc4f74d900ad356960d00e3923ee1b42ff89e144fa295f602b66c367ca0b2fc2931467b83b135ff8396b226bdad1573eb82cce849879be6386948f11114bcd0819d7806be54e3afdd7ead15e274c320edb929dd9c2f74b43919b723aa9b6eadfd55a735cd5037f18e328032038f3b73e865a4ab592d5df6797705af0f666766af59df85c9afb2560d019f34680a60c202c69a82adac30b717d92c446e0d8b031395cc98b3fa8db1a47258484e39d76282e5200460cdd0fe668a33904c636db26187638e9d0a8abfec782efbc8899520544d2329a1538017a25ea3617ee8e87b17b4e5eb2cc42cb09d50aa028a624f6d97d921cf274414daeb72f7fa309930eda863044d5729a79289dbaddca79206c1f46c322c7c9db4f6bd866a0b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h59cf6ec7e2879b9c07e987307dd2def6dfa439d7c7a9dfdc83dd1b1bf82d081f0bdf488ff9c589a015e236c7535627942b04a69619898fea4398010adc0478260fabf60c1be283e5458b627d9ae5320460a07a5ac3672a9f2b925b15f803adcc326bfc4462e72ae4a8cdf10f08027ed8133088157a102cabdab6a26bd0eac2d78d3fe0877e08ac2634f52013fd4b67960dd2cfbf69bf3aa51b7b92917147962ddf613fb9364bdfaeaee0d22b25fc52fa7195664313a4c62e57af004d2ad7c3ca1104aba17d194dac34835295f3a72dc75f59dbc22bc89e1b1c596b4fc672c66b5d1f889bd545580e3919323710709fcb4f2a535bb5d1c46a3a8e330715f74bbb874419f29dd119820e228dca65c5cdfa9132da10bf6291b3540dfcfbc3b2369307cc821c4033892021ebed8bd033c2c1885f7d90b9a8bd3c935ea93669a2c739be361901040ed3f6ebdcace75a3d409c0beeda1280ba310aadfff3cea6b690db2be63c792458aa26bdfbb4f1f3e30f7db472ac2e84a577fb31471b1282e599a949e592eb914f202555bee78708c319ec22d57fbf0c0ba0b2d5864bab49ff433fb9f44f76e42c3787ffa2e3fe2c7c09dc6a6350d9c6ead81fdb887e5ec4b342f6b73ab261304faf929e1718fe32afb5043cd8199560c493656ad6411716c0b31023fb35aa0406d060e9e134f1f8c848909a523657f80cd8efd04f741f4f01360fbb8c2a28baf17b50e554631665ed5e43f8a145c03048ea20dce1ea602e69f0638da3ac652a92311c534cb2c485c6f1fd37b997bc1a02f7f1fe7ac9ddb10f425cb9fa42564bca578b00639ff98e3838eef2b8396d503f1d6c0b845366ff05d8f945e234e8d10803a58ee6f7143f0ff18342e7d02b98804da987cd5b41a1251ad5a2870ce71c939e9dae9457499dd87be5967d0d6cbcab2cdbf7841cfd073edd298264c8492b53f6ab0a7dddd19d4edcb393374c8ec36ef1bce432dffb6fafe346356f8a74e7143c6d98c48cbdf80e201f4be59e092f27312c4d2997050f836f34e0d80ef1a7881a3703d19f7e0d3a76f62967283eea209263d878a2c077658291efb4dc8e456d65fc08669816ced6c14f08ff832723c3f0377bf9e4b5e192b88c4f204c31b24b1655af5f55bfb4d208edfef6c6f1d7da5f5d91c971ac8086782b92d15d160055d5db2cb3a6eb3336c95bab594a0d21caad2f6e5d5c46fe37729e82773e9d5831fcdec4d1f9287efe595dee2841d559f233bc7c4652020d490b4f414206dfbc2d8ad405987a11421575b2075787e506b74e20c8b77fca2780a0663385236b2957defb3482dd736b73a309d3a06021a713825c569407863993ef61139380e7782905e14893a75d0ad4af89966b3755d13169914c3584974388aec694d6838c2232be967651d13ecbf95f8d3d7a784dec8d1cd8c9f6f6cc65cc76c4bdc5b0c7df500020408dc2cc16e1e35f6232e9676339445cf55c0da9c44cc634e00c2435c2760331e927a91a8d9ba7ef2e40cdc55d3d9809567229e0939b9c28e361e1c1d609d7903a34ea91789014000c445cd139ba9fe7e7c0a7cd2a28deb52cc885835170856fac57b8f167338cc6c4d9b26f946346d3faad7b50af61915600cca7f63281a4fe7410e6315f29d02a4c4c3d0e9ed1f9d36e9fd6e8ba536534328634ad1eaf82ec2cca1858d55d2a6ebd6f1cde001a005e3fa62018427da0d8fb62690c6d70f98f1bd2e8f343892891bd3aee17b642f6c41497423d239fd0e232d7d403f8ebaf9e3a3c1eb50b6ab97b6a71912915ed0ceb25dda36ce32f1913b49586ea671c9e49cfe8c8683a72d23c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'he0a7e24962d85bd6adff86d07e4e6b6e3ac56745a357a3dc07a2dfbb257e240a22b67aedec891e9e3aa394c416568af4534c72ad81e8ef4181b3bef02891c7f00aab17029263be313471e43b54d1b082f36f2afe615d505550ba3340147bbc41d6305857a991a283983a9b7d38fcca2eac4614d00fa17194ac95d178d77b1a1be2d3192ce2ab6336b85be590229272984c5814d1a866e8e62836d43184bb51e6ca898a5721c9fec99b099f5959d686f66cda9ba249a93e3d3c3737ce25da877237628a7ab6e1628f180b6050c2e42dbadd4fe0e69aa8cf870ad85851550b43cc10a6a5f96c51adec95a5c644a2987e84161338c5e2cd3d26c017f6e7f33b44ef0e08498344bd621639390b6e9056b1b9a55f81d251d4514a227b48d154169a88d39c861e5a07ff3b577bce8370091ec11e2ca3b42895d5bc394182a40aa09eff8e96eb0bef5b8a2684b1b3ff001773296436f87b3be97f44e7dfb0e36aa7d7e7c0a213d45bd443ad24cf09e7cde652636dc59a61a2a9d4952ee5ed4d39b6cd28ea3de2a8a65bb506f50079f3447970c655d553a1033bea10c3a958296d82228b99c513fcfe4d312e0ebb1117167c69b53bbc40bd3c2ca225930a9f933570ba5af43f680a30a25b251ca1755c21855009766acbf468810a558ea5a6ddf31fcdc59cfd6b21003e58f97026efb6e85e31ee58622238b675cf61d23602963e02d29bf8423e0db99327f163531d675cef806a6de06a91f3bad5033b66d2b4e022e57508b0043d78dd4fb870a7d356075fd3f0a8b1804d3f79473d87ebb671efeb3bd29ed2d243e8a7c430a47058de2eea74eff59d46bde8a7f448e1575eac8984065f11daaab0709259f2b5e0ac7f4d5c266f6cf75e60ebdec343cad5064617af65040c3b403699e649851a1a83ecee5b87d844e5a7c7c5bfcc146ac723f3fbac856442bef9aaddf55c7e15946cfac4968b8cc7360be197cb5face78e37b30fc47320c76276a7aa2e2d5a4839b5a5e41cc164b5bd2398ffaa7c6011063ee4501fdc8c1c29fe5cf81e3c12a3bacfcc29ecd56756629b78ca334812890b819f7e4374e9b890c0f35823b57f4ae9e2b3db5980fbd78583c7a3612ae3a10aa6f045f7d365902e82ad8bd773a7435419456f062622b28e7b1cbc43f41527a893c8d63d97882bf419890637133bde02ea4008b2889ee119d11c9f151de80578f51f8d8e25a3932563c23c1385842653811f88d990f89b66ad99f17bfe84800993709fd8a1ec6ae9c007e2fea1e7e7f42450b79573f943f76508607eb87bb7c74d206b27edcc9718472c06be8116ff0da276d823c7c24c1b964367054208e0c88ff92f9b8a14048c035ab480a72e7275709bd7f924cbf85cb12e604679ac848eb11442602239dee14e1f012476492b33449df41d9cdcdbb52d138a20012a53e68e874e0500e59d1f2b4a253498aff54b8c913a91943fe174856c58bcaba575cc806666729032b68fd7211cb75609d4626339da9b7127c1e0c024dd49689dd753bbe223d2e9d691682f467daca23b82df8eeb893f1d699943d32253ef319e160630c29b9756b7be0ff48e1d3147f22af76a84ba366592aebe4c573db66e34f7181018456c80f7af82e91c01f653356ca02c4e23c48b1022642bedc36ba54160c60f3dbb0cbcef66b1ed3cec0393a7de3663cc72354f2b72f57c6e9a8037132a6bceb1b987044679196f51be1615d3e7da77dc43b5e3a1228d4fd5a39936868d3ad1153c2f6b189c3bde4eef93b79427d71af65e37e357bfefefc628e3e09dc23624d73b33f190249e4766a27701bb7ebbee020ee3f4fb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h4ae616219719a56dc4376955196b270bba720771a615bb3affd21ef04e52306c5774e5f592feaf5b44153668c2119122ed8aa15dfffc41a1e565cb553ff2c305b258e91da669d1617e756fc58e08a012423d12b3ea77457233bac90960e2251070edf443e2282c1e0c801c684f02a60a02fa2791a06f258adb961ba72a2b505bf6a98b10232778ee17a93badaaab0c2802ebdb5dc533eccb1120ab30bbccc8a9085dc6e0d17ce1921b58f22e4f04eb4d1c4240fbe29063b16d55d37f71ed45aad263a6eebb1b672cee6bde98768fdf26a35aa2024755c1b9b485f64b9b12a44f0faaca7a23207fe8288b876235cfd602570b66c9ec0d1b31d0901efebe4b0d88e4d239a93275ff1d9a5305a88f53f265a6b739cf54ec8829a8c8b0757363f56e05d44631695cfa6ee3a3d5549cab36671af097bcd9c96125467c11ebb894c0a7326c21ab47383a09c73ee2ea070f1ad773f8428d9b454383bdbee2013704e51117ce83be41fd2b86171f9e2070a25a383dd729888f9101e8d510de59c4c5a50fb7ddd7474c5ee4a723c2d59f3e8b2e457d2e884a6b026a09145a783538371eaf51bff3e845b12f32fc1635853b4de5e7531f31aca0327a0d381081edf858ceea367f7d7aef006700188c1b84c28b2e3e2ee194d2aef230adea02c46751f8c156113758a77085ffc2f6cfe888a3f4ea1f1cfcbf26e344ba13e071de7ce0c6fb3ae93b968ba5a0eb6d523393992112f5d9d76ca9db62be974ef91f8cb6a429846f6d8de18ab505342b3a38c39b20009659239d9dcf50b4ebc34d1cdfe2b3af041b67205f59ecc39af3412f9f6909ba0bb5d37b4a63636978a7f43dbb427fe2d3ac848f7ca85220389c24752662fffafa235fc3da424e797b37c66188dfab7feccacd04706357dcfd2ed22d0f5a2dffd4856c6614d2485ea46f135dd8e3ff94621a741b82eefcbff9e56dc35814e68c4349912a3e519b2931f0cad27ed2fa18650fd8c4fe62c13fe50cd284478e716fefdde54e775e96aff29559cce78495ea7203d3226950fb08a32f292765f0b5ed42c22975da45f87718df05f978e6ff96f788a1c19cb68798cd5a761a60ccff83a4f1cd95533ac3cf4f0136f92b65a6a78a54fff624fdb466181db1623171403a1eab19e8143699ad7437aab8fbfef57b9caeea5d183a20ab92af459eb79fa38b6697940208eb8a00c4ce7c46c0a6beba27cd7602950907eaaf29c6df4a1be1ba948b37eb9ba4109a2356dcd6aaebc399c375404ceb97d03daf7ad8486410aaaadcafb9db7f788d21251eebad9a26b72de970c71e2e493a326fa65b6e6b072484c054ec447a95e5a97db2c78737d453e284822bbb8cb1b6e24125707227f3b1e7fde8f2e93e0cabdacf4130a64e9c9f4f4f3a91e2e5e2bf6b9c33df6d5bc694d804b9bbb20c6fed74af64e275cc6c346d33456aa12962390427162a86ed1fd56a7ec9e7861239661107690d31b60a357ef8a43d0987aaf2964dd9c418a9eee53671fa97543be3dfcc6633f732e6eaf801c5059b636da63151210d71af1e25656981194c4dd1737e1ee07499803a18bdb3e35912cd1d3dfe7442350b097617a346b8a6e279a5187fb0e5535dcbc6ddafa6c15bff906ea80906ea2b1d7d0f192f551188363a007fca1e12582c854903e645bc81b60cb003c49ce340938490fe4d635e2f02cc012ec2971e7b35aa232fadc6f1b8af5b01bc975274d151284a6d7556c7b80ced9aa3308368271607f07c045bfd00026c0249aa4de5434516391e1eb651183ebbc9749f6b069226dcd6230d529e8f89d8eefd77c24a2fef5fd99caa963bd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h83710f7c04f573a471c3d20d48f98e1ac36933cad22c275161262b4168f0e101ca9dde7781c260968fdf2ca2c1aef3854196d230473a20d7a7887376b42bddccf2547a907050c9208be942dde3c1ffcb6c8a09299f390bafbab7c050c1021baf1ceb4c1d52fdbee2b1c943ea23518b17f52348eb844c34729692b55fc8ad3c53e5baae908c1634735800dc01768a201c31f0a38273ce6afbbd0caa9e13bda5e1001e3510a286b875924bb2524070496b5e924f4a3990b7f83a37181ccddebe167731362b7a50d9214dd7d1632a0b335471075943a4654df9a7ed1a8900efd5750eae3a64edc11b8ab65431dd37da10967ab8a0aca5ebae7ef5c5783054ee0cc73ac92afb6bc0fce5ee20e14db0e17e848da183e62b7931530c226ac6832c69d13dc6bc506bff3d0d9994c42abf805671eb76fd2738b28ed5ed0e5ea6943fc24ae6cbb6296366bf64492a2c5fbf2f085d1c5562386463b41ff8a296b6a54f9c7f63ec874cdaadcb05b7286a0406f50b439a1ab6df7c30ae0d368757c251a693f0f7d2365941dcf176247717838b36b74dd30215154ec913d883efe9e278900bdebb2426a7eedb2d90538d5d8336566228e54b15ccce60d763f3b55e80c1a3932e04c3fce36c68a4c607199bd253a4695585ee2e0ad436621def1020af554586c875b4c5e5f47a84e4766e79371e69099f25bd93daa33cff08064e439c9004024194bef597a851a0774b998e5f83ff218b1565252d561e5c6ab6533e1f2f07f472dec5882bda14964241b25e66946ed0aacd9a720e199690a7769abbe023eaa18aef606131d306563899871e8e0f5cc2b5838d240a1335e90d68884d0ac6680a2d451393d2917a02265fe66a0ed6e57f3bdc88b74a28d40d44f1df71a1708c0b5c02b9654aed85224732719a8be7b5f8ab4e7bc85012ad65756f601526c810686a906f0c41bba907ad25af14907c2375ee59ec3cb3fa6e280460307e45e24f6ce8c94cd8af18901d0f9310f2170204ac27200d4216dc85c1e345baa9ad596d467e0c3ac1fa66d2acc0421d08a7c2fb7bc8fc2d5ae9839491eea8496375d071d36b73424eca4e45fd1cd7ec453d98d8a754e572a4a56e070a650cfbd8b15412f42641716c53ca2db39cc7f0eff51c3a3200afe480ba436fd6ab604fed01201fbfc4081b4d4a45b8c7ffab9583e182170c25949dee7efe3dc143cf6a69ce1b6630032fc1d8a15457aea60195ec278ee373ffdf0822021f6728e00e3e4de2f061919f72e9b55238c79ef4b18669cc34c801affd7eb3a9f48eefcefe3d21c982a0e9074724bd30463b8635d9a63e0f7738d29f92c9e62a095b0376ae32bbb6bafd02abb8da570783730de754a60512ce74beb768eded2b9ae28cf43855b610f7a8e62fefdae355941f8fbf5dc0c22dafedc48bc549049d8bf9e31b491144aa2bf9b1d8244b28b8cb730124c2819c17765799770fe69587c62f47553ae3cc07d0a8480b6ab9ce1d09cdcb6a560e79d526ef4957893fd70b7a5f05f05a5342869e626b71d5ea44247ee6be3d0a2d4b3b8f8dc87b6e281b9005bb615893c0a6ecc2ac434d8ba1f2bb1b9a653a6481c09ec331672f3632bd1ccf19e7519f9719f08571e45f0e5a7d2915301b39a12e12e840c111dca7a4c14737dd89406fc084ab8e0ae5ebad4577f2c17a0254cf14ba296763a72848686c60f5133bcc7255d11e48f13609816ff38ae88839d3fd2c09182d3fba9eed3a18e196fa91bfbe499141521defda7e30cbe1aac6607d08d9a48266e4ddcfc50046f8ee77c44a97cb8f481688b12e6b21d15979347b2aa8dd8be40476f151;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h11f78e5fd87f35e24f3d9d83083a863aa059987e9b2bcb48e85a71d7a6d1527f100eb69d573c2a0e824e4ad4502fbb3df492ec636527c69d00ce238962c622b3b76898a9f93a8ee431215e8bd2b340c98aa41d8d3804e0da5daeda7fe6d1e9878d78c75b5d63c03dd052543bb2742b4c22f24ed842cbb40ba69f77a7dd9febde11c7c83cb6b45f13b590e4cb84a2c07aead883ae803846ff01328e5671d0afd99132fb9210caf206f6bf30b2f681cce92f3f51ceed81e1f6dadbd2ac9b3af1c1280ed4d2bcf0db70d6a78b398eaed69ab01f030dfb9658e724ce756adf493f1abf33b0f30361094a2cf442d25fdb4b1279a28f9edfd6ad03ca960942a05e6a8665a20a9a6366c44a9ab672fd63dcba4d45db643519846c9b01196aa3d115efc04891b3be8594540128c57a9643013ccab5eae3d1cf3e714e515df46f09eb75cb84d55ad8703b53677d75fc2d1c01c68f92fc27c43232c800c405ccbd046452e6a32cae341b5c6dfeb4f9b3051ffc6e0d5d90437f2a9bd6548a5bb9e82454d1de167e62f824427259d27f8f6e7e7f1a5c2a8059f023d9e0785595e86b3ca93d931fc0de96ba446e3a009e225f9e16cb3fbdb4b8d4c8bfb91b5cd2def9d0716393333e42fbee047e32d9bb74344a742965efe56fa0e2fe5e929027ad6cc602b9608853c9e4a5f74d02308bc9531adde117135901493747e3186e1e1a7645811cedca5d3b35cc284a64ff651eb93bbc36b3f8e9733d079df3240708db81c8aeddadfd4205949e1dc3534651fe6c1c81b8429ca31c0ad595c9c02614d477a95dd7bb7c7869e6515c5c45b28eead20360bcedaf7eb05410fdf97f10d914b0b0a183bb2fca7b223c9b58a77ba54ff693d5389b18bec7054dec38d08634f2292eae60d233fa404c6e3b3b27265516408daabb6b327664dea915823bda7faa3a402dc2af89ab1bb4523e509d6793096be2c95a11d96d46c75647f1131428b13874e44f9cd9320a72f0c7cbbc481761710dcd0e2a7ac62bbbaebef4538186981b203b938ba0a53b4ddc3de30602559614c2b3a6abc75ef796b4fa26b2a249455e08b11353f49d28bfcdb9335d887df8eb7d6c939080c41104c36a88c73d430efd5ff9bc9fa485e9c224bb554d96b3ca873d43610d0fb916c974bfc33474657a8cb35ea9a4bf145818177f724991311acbb3f8650980699eb95ce2c9e4526ae5737fe157ace860ab597fde328a21917a0ae3ce3326106335cc5c71952b5f397267cf53dc35e0a17b0b0245710775471e000d66b48d96cf107faf578624dd94c55cec292d67a7467b09e9e61959e8b91c5d13534ceaf22f8fe28d32111c87e2f48ee8f820d07f0648fb5868b39f5499ee0bbd19646ff9aa2432021ad0d0d557eb1b71080ff214ce45e771b7a5b813954aec06cdb4d6e77e52d5bfd7613ac0df1b0239162ab5ba6ffd28cce6371af379900a4fd06e809f16ec1ce79492b122c0960cb2a855159fbad5d23f071f2a552c1adc3dac396263bd44a3b5c7e5fe8eb55c24c94515de3c0b980e6442fca46487a88742254326dcd91952282d9d6a73e3770b4f08ecedd9f1af9afa152c6e0f9fab6f98a2076b4319452f38764dbeba3c6835ed73c48e481f06bf76839a3f9c1393b12dac1db84392b2720beb9b36ca6b8d0fd22b0192f4e9aaaa70a371f7d30484bd974dc68c1b675b8cc0393f27242a46e30777387dead7718fc0a1bccd95ea64f9e348340003b4ab0d6de5b3ac8cf5db280d147aa8d061ba4cc3cda6c2040ecfec8d6f27064ff91bfe2ab03a8b07ac712e387652ce37b4deb0c6f685b895fedb5bb6d24c9d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h77e36b266a52cf993f52a326db33cf18deb29fba8202f12b3d5f628c5949adccdc8e455020dc6f672837d854b7ef69a3963f44c5c12f93203e68085681ed9e36dfdb49f2a849ca149db12cb18150c6a6bf3954051ca603937755659746738d0ddf2e6fe5a6312c2ce361577b96e0cd05e3cad5aebc3b83ab543bf28f8141847dcfcd240b6a97dbe935ed98171184bda22f757f1c152aa395e25163938d2b08bdebdc52f130883bf3109a8bbb3516718e93185856c04f59d418e6f3ca7c603641de760af17bd5abaae6fdb276da27b121913ad0fb5ca9c52eb432b55fd8534372ded6691950d533f591e4f2d94632ce0afab5e0ec0006732b393855b881f3dc82b751253375a985b59b94cdcb1e5f05d6400dab9f8595fa9239735acf96acce8b33dbd13dc8ee63da3ab9439253158954f14d1d16f3ecd737b5fed0204ae7125ff54ec9159fe398a875e6bbbf85aaf4969664feb9b3932ca29cda83988411b8cc7ec75798f7fcaf0b2e7b642495464f17ff25b663bf91f9f4b50fa8d8e58dd0f3b90a25c350579eef1ba8398c7f2c2de69d3e467a6a0e0b19e83027a5565ce7686d8f0c9e71e70c001327e1fc849f9deb61e7b9e9ff25aab56c6fe95e410c144175935cd404484adfe5f1cad02c8bb993f734f859d8d9c57d3e365d1fc02a77f4f3111c59e1507d96d72fd6428029bbf9df9c4708db274e9e6e66a2749defc668a6243a75435999ea286465601af2bcfc2ea395ddebe9f2518c4ce095c4f5314a8dc9169ce49cd7b5d10a6bbf637544c01c03f5ba48bdfe25a9c223af6b7f6ef88154abc740e0b242dc3fb11b81209840b6d36610ed38d52996a779a8c3d843a7d80970785aa71ea6363991913725954e9d31461b948e6e92394f9756faf6fc38b2bdbfb72600575d26607c3adfc58566e2fd2d4ca9487a24c8efa4a9c2d922f8a895ee68ecb9a2082ac2a3922a1e4ad741f24de7a4be55dba1a30bbb96d0fd017cc579e9cabf268aca8e1955faf84055d8db0f33450db3f7d77b662d515688ed2d7b891a3ef35a6149a837a300be75bddce7b958d2b9b397173be0f60bf2972059ff9d2721043f3c10b282b5f9b3c588e8f864acebd13843537acb7df2822403d0d812fe232eec5fe62b7611b372f14068845d0cdfcaa4e162edf0d148be19514b47c5b4d9f9f8199889e9441c03cb8066e0891113ef6e5a2547a533c71748d0810a442bc5fab1a4800e45882315947e8eb210db6042f6539dc2ef976b78e6ab5e3332c67727bc431eac3618184c35f305915006e0f99a6f1b3510cd5a8a1449179cf5d529ea8ebc988d97c69e14e0bee699b956dbffc956031285b6a2f545f49c0934964d7fc6b9b1377558ee98ee5c72634bf02d47848c62ce1adbf9de6c9e586b2809ea3d8b6a3eb1e87f5f6239e4d6d868c269af6d9306f5c399031385ddb2e28f2a2764294aae669f75e6308650f484a5e9512d44b074c4669a3175616fd0cdb54f14d8930f48d2b8e01d4ac6d1206b3781f0d9af01cd3d4dc6779a93a589f2d2684c6269b6716ac98fd4f0a6209d86ad490a0810350b0e9c7113e4c56b06fcd53eb745f1eaca32b5fb67e835a600507369c423a9dd33a5305917738da6392c38217a8a360b03c30338b8b9c884132a8bbbfc2b45230f12ab8732441f2e0028209d4c93c3853506f396d304d0c44451cffdda7b901be171bcb7c2efea2d2865d017130410f507bce30830547223c3c69fd167ffd15789896ff0a5f85ea3b7b3338e7cbded314ab801ae240c16e1201648119324efc49b3aeeec00e8dfda790d61387a5a1f53c493fc3ac49de620;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3e88c1cd2fcf7470117bd67f9539eb57f59ccc2ae8d22ffde824f53ae51535c81dacefe4f72d8ee655501d13a262ba042669f0483afd33a0a3c9ebd01190c253cbbce1f586ac6e7903273d7c132a1b02634ca2866903682308b4489521216569c8015051a7c637afd6cc2f1ba00eaa2f4755b8759c4837c0b23721078cbcc2758f50f624d81bbadd76483890c7c6241bed538576338146f02925b5271232ed55fbf25a2d3cf31d88d1d8fd7140bca619f1a829676cb3fcf5b0c75c18992c73d9f8b689865cba96f8173c38b96011d1b1df78729df683c1237db82ca43fac99e5b8f900e6454164019344503527cfe607a3938aaebe4de71696b7234f5d0120c2314c6008af39ab2632aba5d324f7a3cdc3ccfb780282d94a168a6a616599b5a06b0dbc1a76896e27849c47afc9e93b21477bb290949150bf04d520e35bf2d58242d68d69969da4515b574f3c4d9094ba050aac57dd1a5a4bac23cab28071fa6710755260e3b54a13cc9d88c775ba918084a404615ef489dd9e783cbc9a871706e6eb3e0505bd7fc103ed0fee8bd196fd0c89cc62ecbfa62149eff9a18c259d3719704a87c14ca2985a5046369385a7072ca8068716f63914796ede167605c3979c6fb6d8c8e81fa99d0bf830279ab75f878aa2a2f1cdec15b83ec8f459b5c953ebd6904ebbb12242925e001c8ccf6ce0ad5ddc59db515fd18d8ac956516fc556a10bcf4d2a6fc4f88cb5a1c90c0cf77c442079b89747912ee9b81472fdf49e3e5a3610599bd138a54e0244c8851fe9c542ecf13f801fe961af8be3c7bbb1d9472510e6e11ac0921be2e579a530ede5d534c309064251dc8da55446304effd3fd3a0371f790f80de076aa51c96f1e051fbb3448137417df7a5efb1598e1a65949ffa68dbe1b15a7da7dc501d5f6245c7daf08d2cfb7ee710f55b0fc889899fd89a1355e85abe0d3a1eae1b5cc23fe5e62524179252f691c7a9155a3038199c6af59b24593c6f29899eccf8935dea284904b1b5f8032a2c15206c54d260f342b9ed34ecd6858955a765e1e165287706cb800c6f79f2e4bbb7e3842ebfa5cff10879a7dbff2ca391c0ce08a26b8667d7a0aa76b3035db0c8d698abd2f429c95abf11adbc9ded024906f3c5bedb0692ecce42b42802ad7096db424888f1782113ab412bfe4143cbe9ed9ea9a22ddf91ba539e558d5f7d43e99f76e03e19e70d6bc1ebc67cc04d9ba633fe68b390993b55aaa4d388957e28fa6636e603dd26458149b2bfb1f145e70ea50867d4ada1e4b761f65fbe0f6ab490fc74c1ada54b4f3d38da5f521363b6d2d6f2f9a00711f2387f4e158b9e08e1134537a889523c7c30a6ba1a3ae90cb45b30bb5b317d40ee099222ed0331700b918916f9300eac5b432e068e2aae2c574b898483afbc4e6282d9d4e7652c9f61250eb3a1f413aff509f838e623025308f4eb3352ff96c2d0748f01784fc9ad75afdf12f83b78c087026d74efa88045542e56cac0d0ef025eef74092684b73fa71ea1a2b7c9a90ec7a8b8f3a5b50ee77883bf08ee2f5f1d97d371038457904a638d0212c8491d65d68c0ebd56bd00ef5398c65dadb4fc3a8870fac780b111a068a42135c10fadf083361d0f8490ec962123a4fd64b1a9cf3647fba13d112d819dd6ad1c4a981b5bd8b47ba584a2c3620753a73668c3825dc8a59302c8f5b62427fa91929efad41a4ad340a675c970440b9f269d6a0f49aa2cd86ee39e350ab445e29d334fe28be5d538f41701b0c3c66f2ba3d3ce235714bd6e13ac88ad1a6f391774503002c1e25c146b1ca3b92c665c27f8fdcaaccecef473593;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h739b55eba334ceea54209a1aa0f2f601ff1f5ef344e5f4bc361813d9a39bb6ee08ffa285ebcc51264fb80bbf9564fab603b0db1e3f4746e74231ad0b5b72e47ac32683722461c187ea4964f2acf50006cab56c69c1da3a1b3d7072892d8c19d151b7f3f5601fa6c91f439bbbfa36b74c580f2f8b5e534f6a27226a02d5221a68ad7edeccc8b8bd44750790016fede852efccfcd7b5fd7b2a5c08b1f1161580c597b6990b879a4f07a0b08c54d4a025ab25951cf22211189bc20555cc040b8eecefb607dc53208bdd4119ce5f3ef6a83b2f668a00a2eb8989e28754b79ebe8e3f523167cd3cda7ca38b43f794cc1b19ba86e95c94c2e827129ff88c3b9084383c39b52eb7932e440770f1d7f8de34eea94fb73ce204f17f4d2e4816e7ac4e89d2702bf50c7926ce01e328b123103010872d68641ead953c6f76541ae16c0988ea6e22dd35df2e40cd3807483682fc1c2ffe41347636f0b89133e810ca8c40c7d0ffbf181ecc00aa8d9345bdc4327805a85aa8bf7406d15bf47694c5a9353a313c900ba937d276c408337b2a68caf8f318742b6ad280e5d0f75287ba2d236dfcf01c4e198fe69aeb0df3266db5f6ec307caf07a82e1948f62d77ae268ed1f52cf232c15e31962c986bb3a6431700da16f971c455be446e00c7293494bba5cbf7444748b4620f6ae8f696c1d729b27ea2088da61575b4063c578c456fae17c59db00b53b65af6194f010abc66a952794efb9427b4774d6f4c227a8f4fe7ece6c5e1f89216f421a429d21834605d18010d252dc7b6d0cf4d15337b61decd4abb27f4f9cbc73e7944934389d11ee93e1f1b5fdbfc59e8611e60761cbd061c9f34faf984ec9b1aad14b8fd1beabc6bd6f1e15a84cfdc496c6c6a5abd40c03aa2a312573711e7b3a8661dd8ca6be33acea45036cca3c9981e520a938de6b6f57dd8c608133148c35b9feb0e55732056eae2bd3d0f17fdb9225bc7c7f75e17d482c44cb1632a77efc2237db68136f07925cd3738b3dfd0d9d0f3582db644984e9b505bfbfa4d63f812f2a64c0600e2b61cc7f843a93d7ec81eead90518942aafb871b30cfc16c4d5fd24e12724594347f74145516c45445ee15a904e041afa6eb8b8d92d9f1fcf676a106193050f2c822d021ee7c609173b003deb9207ae2bf3bd973b473e6ae6c4dbd3c89209cd24a53a6326604550e4c1f066c00456a61de93b93f4bb48c18e5eed945ac7c3b2a5b92ae097ba5e5e80ab97122d1bf40f4effc6d486304290a342cb08c4de733f2a18c533dc4b6e301b6b2178ca65938992d56b933184b0a12f7d49f85f88ef39b06c93d3a857d50269b20abfa1570d6f249fc8f86e05bece5a86bff816e4be1419eab15a67c04dc426801a129d6f8c9830c41d427a7b6a08e74f5fcdaa027407f4451a21ed73cf7e1ab0992c6c8a942222264e8721ef7ebbf8e0ab34c0ed8b0b8920cda7e6efa3e145bf0963e21e6af139a5e0294dcf83dd7e8735f4c8eb2fd26e91a946ea8b779701e20be29daff6de9336455f200a68790fe652e93e0e4172a7de0f8ec446aad01900a3a63cf878254951b4d99376ec21652af5e828728fe4a9c72b3873d47857de00d4da1b24c3c1edb00b13ce4c18a8577d5fef65562a9169d0a2ed4ece3fd27632bb14f873a181c4c7a5df49d046a4b81fc9aed4f2aeec933266ff159ab8160d3d5599292a4a80419da0ffe81471e19ed653406d39ac01cff2944f0bac4cc11cdf0e6073d546a3fe27731bf4c0eb02ccbd73320ebfef30006c076c573f3dfbc688bfeca05822bb9c2b40a4b5118eff90a1622b71e6ae23af34c201d8c7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hcdb2a25bfcbc6a81e01ae72cf231950a065d63cd225cf5f4f9a193745d910f510ef4c52b40e10cc52999ef897d8c1bdbd5e60ec71e098d218361ab739682448987784dd2b9808b2ec31fe0b87fd1f1110060da677916fe8a44de53a9ebf2ffa4ef02601a0825a7d4953ed0e84fe39cbab399eb2bdaecef4b59750a8e4686d461f80fe783389428060b27a65b7d8d880323934d277befb5f699a5439002dbc894b0fbd5e4958ed85cccbf9e64e10c57b69369ac735c596f105c761db76cdf89b76d586e3d4efbdf740c80e7de34925ba9e8eeec66ed4d31e64fd1191aa4bf78364ca91ce48d9576171504d88463a6b70e281ad320f3be0fb7da9fcbbdac92d0897459432d30bcb557c7337291dc191dbc849842d09e7bc73fdc4cef6c3e63d0f6aa66451ea26c8287b0b6f9ee5075d0d69905f3349538797ae08dd5205fa15e06a5488e1f138dfb05d3a14224cb6f62edd0de1007afdc4d5d92ad7623c1c37c1c2576d419c96fc81351617155ebdb231fc17742e021fe99e553b742d60a47141e912dd2301bfbd7bf520cba6d86be00a403557745920b3cb21d2a435a6e2eab60d52cd519428c6bc07664545559af93198534512e857d0a04a0ba10fa90755ee1923fcece1e38bc3c33efbbf4225e56762369070cbca1a1e32cbb2a1d238040290a20286d95f272dfe5150fcece10961c52f61e01b148921002d7c3795db22d7b0e093a06fe8c44a75e9ce5e21e76ba5aa77e287392add7d327c8a3ec291dc6cd9ad996516003cc26c254b3b1defa14376daaed1b194470a2504987d00b7403628f0d62741ac0e6e34a8c59c46b05dc498ab2536243a670a315ff778f26a3c7d51cbb6bb37d5b1b951a27fc0e6d292fd1a809f5feafcf2c746e1df41fa9de25872809b33152c0cfea723f1c345f1f9428da98934342a5b229cbf2d9321a866912e82b4f056a20751b44a34b3bbe2a141951970a50b9c80a3e7aca29c8dda67ab1efc52b80a63f21dcfc3adc5bb5e098052a9bf8b7646b3b7b567025165790736fab913f62cd638a4230f4535cccb913010e2dfa98b63e57a2fe080eef2d764cdb8f533debb8e91fba8483dd4bfe53912c7832e51f02af5bb789f6aee210f20f686303559caa3d9dc6df9aca5ea1be8efbd1738dbb27f509f0abf2bc8ffd89ed77c631109444e8aa3ef7054fa9c255bd6841a2ed7fd27877fb9d6f1126b8c42dbab98851e2ce22e7cb4f83598cc3f0bb6fa8a76f71d0cd9169793209930950c6355e996e4c512f86f51f0e402713cec9c025c726c4109d86916269eb73ae87d86cf2cb090442085549c4034d816627c4afc529b728219a33be7dbd12b160fb40ce46e0bbd11fda1f6a1f58864f4dda0aaa211fbf7b18ba9a630465e0ed45b40010b160d20b07db0a2ed4e3c89f1719640b7c467f2f0d5bc61bccc4e2845c842fed14f11d9cc7c7ee6e36fe14d019515039b8e003429619d35b429f27098ca30374368346074d091af5183e930da84dfdcfda85b7c66e852d7872ae5e53b859f5d699fa58abad515e1ab5d902d5378e2c304b8fd775a71213eafc0939aee6c2f542bf8ed54b5b775425d3900c6408f93119257cba68272ef0231e02be9fa64ef751484da603158c8a0c87d10dc844103b7efbdad4f05223a23089c3fbab985ce1bbef6b0b71b577a3b9993147adbfa3e7c3728f26eba5db67b554eec2e5711a2911c47efb59cb05a3111e551c1aaf4ca756a6b66a670c163f4eedb21d7f567aff467357790d49521f6fd1e2b9b16c4b2354a75bbd263b0e45c6cca4fd64f16463d91a1d3fe13bc564fbd8f305b6b8a6cc27;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hd3217b2c1be860211696f3e64c01e61e7e376d86109171dfb51f512ba3d37323f38005ee7fe33d6d1e4d06ddcb6b977b7bfc604fde6ebe7b593d1075ecc30d7c22b029ecce5f784b43c7caa203a43be4ddc2d28b4e013f1f1744ca61bef7396e515c1cebe43ccd01ae3e486bf835b374b6d2bc1a4e24678cbab995db40c74c61fbeea2c94260a4feb621197b9a18b12f6613c957ae64808a8869997c5818a5e4a7b6f8bf81dd68232a9e9659d915a86f46f6478f8fa063de8ab6e759dc403a1f0f5e1854dc5d3d50f8e20b3e8182ec80e94c4eeb8387d3be014eed26dfae560e8a967d2ecd25505d4362175fe65c75ce8ab380d7a8616c76946bf38df33e3689e4ea25e8117cb0c6e9114daeed5df35a475f1f71da1b1b07dd2f639e109e6b9ed9f70f4e2cd28d30150926e04e68b2b794077b1c7380bade4f2d0c31cadf1d6a36b47828176d8ebca309dd68317840a477b132003f4b44cd8aa427dcd5a47bbac0e00f8d2cad20baaff867998ae5983fb7f1c4a3268ecc454de20d18e510da3335c3f0a463e98ea1e68a3cfc45cd24974639b68081304037d92d5e9413fb9f3f0d2b655325299a8cfd7f9d7432657e7a3bdf911b0ed55c9f2439ddb1f4c59ea86520a135da7055ad51503a3875fb7788a98b22d2bcdbbd506e1b88e26015d9a5c8accd95391473520ec68f9ba39f26e09b0f7b271cab36b3e6acf7353dc2cc258f46f6e5365e3e11e3d933a30b93dbc03bb2cbebfa8bdc7cb2863e4192ad1791106c241d9f978b355b626285e441b866b1b3a7d79d3002c6e07a7f59ddc83a5310fc737b621af8fdfe42a860474be3c0e386e0891c7179d4b51eb99123131c7f3c1758c0f3e2c67e63ee3e1cc3e59e4c22796dd8bda1b30cb4bab533974883b52b31f1632844081ea93bea50db43afc0ab8d35a3031f0d552f8b84c6e01a4e37fada4db945fe0b5b28ffab95be3228363a7ad9541cb258e9a22996daee1ee0b10884ff7a883c52f1e67a6800b55e72a84da895338d142a7b67e7ee3acc4df784c19b2a0e39196d1f18578ea7c3800253d86dcdfff86ea722c85034a6c82172ca93dac0c7ae2516c047bed6ab8220760e26ced4a02d502513ac3a8b557ca8306d1f3e057ef5c46d12d85ce0454e923615dd3540d70a89e2caf81f34c89369f81639d271a1918584fbc9435a0fb2cb943c3e0ad5f5592b74b04ffcbf10ad460e1933114f68b6b053a0a33688a00f7f5d9438639b6d2fa5ea50f26c8a2752bea1c3aedcb8771792cf0e54aae2a6bd89883616d3afbad0cc9a1d451e53f8ae8547c5705ed3ced9db3eb9c1d20202dfc9c2fbaa464f069b61a3bacab2b9e8b96eb26b5f420a159632e55a462398d062c32f54adb9ed119cfe0b14e8a845e5a2b39b313e0eb995c69eee6d6e47b8c796ddd44ee096bcac475babe6337b446182be3e9b3dcdad3696f809dc84dd80fd5e12ed7d9733ab459dd109ca50bb7f5a27c2b98906a692d2bf88a2b3f6869f3a5cc22f79a5192b589beeead6c64abaa5c299871bb596da631b0def2377318ea1c9bfc0d3f3da5d1b05c7c4e73d4281354c90897baa4bfa71fa40120c4e1b8ea7c5cf2a4e05c3f648fce6b26731a0ab71b812460344d714b2a71a9b8cdb76c340f511bffce934c16d8f33c686f25d93697bb7ea320f6f6066a51f75137739bd7c33354d780746917aafd7b620b72dbebe5ca063ffc12a5d387d8732d84d77fd655d35de918266cd3c94c8e05050f7446eedf6bd52eecc1e47b21691ae3c83b6e4c6a46dc8005a2f25a6ad4e823ad4c59786501ce41d6a8317ec54d5aeaf183ef64a2ab96f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h9bf016a8b5ee3c529f2dc04ea4840d85c945f3e8f36c4a6cd8ad8a6b308f9cfc6f480ed1b90a862b5dfe6b4722bbf0d8efa1e730f52cc3b765010b38e845c97bce2b33a22e707b7e570489b82642bc884987070bf34827167d7f6bedf2c604926a84842d750057aa99f4dec06faf7aa5339e3dff072517b2060b430c98377bc16388ad666ab2465c06bb9a0e631bf7fda4bc045ffa2fe950332314e2f3029e0add24bb7d7269b93e47648887e8ddaba8454d25a25b2a640efdec64f37505571429ea24f72fc72b07d49e9f07d3020ec028b5c11a86bd7d81d26cdcb05c2e54b44f7e24b227b37d1591c97c250ff97998b5c907b95c3bd372492f91770b7be910a5634f8af44ce8ed1e60d996a387c94e962b3d0220eca2d5256397aaa26f077d7722bf173936e52810dd04c173e5b1bba6b508f9f1b96d58b6d80bb84213274ae5ecc15528fa7efcd87a1387ace270971516244c64ad1d98c6f0c94117fae1a5e741b361be4c963348f2c8f689db9787b2ebda54f39d426f6a87a430a3e65e3d15b9e926b1d4e1041ee825f3875b36f4d73da33fb60ef6e65c026f800cc167000d9a51aa500eced7c4e5efdf1cbbec1fd2149a2a14e90329dfc4ae3cca6a8bd9244f532744062fee015ccbcc9236efa510525fd90d139723c1883f960a5c905f772ca14629079bc7536bc14dec3a799c84a4c8593dc399ca4921a36e52bf89e44f3af51f4786a15d4708ed0aaa99c53b1e212516482cb24f5690cbf748e3363d7e6aca7414c64e4c003ca04486fa3dde5673f633fb34db10ebc9461a649404a4bc1aff497b86d067eb2cdcc0c2d60a022e358faaafb5ab92076c898488192e4cc4f4cfa3826c96ed367f7c2703e56c85f393aa9f32dfc3a33384189f33621dbbaf9cb74d55b425135c9bdf3adccda13321d5ef970f50d8a160e1cd39c79f2581495faa897c5f19eec984775d3949bae969daff3f74f7bed60f2813af6b6cd77b9befd97a8fd2e96b724d680daea508542d804771689061be6834322a8155e9f5e53d292c7e861ea37ab5ff82bf19afc90ae2066e12fc2d14653d9d35ba6890e6b8a4c3744bc4ad0ee7c5be1f36f3c9d949fd8e6ce879b2c4af50ee4db77e2876fbfe5e3710c356a2d64743498dbe1cd8cd717fa9ea66a951698f0a48a7a7a3538539c2029a636b0db5f19facbfa18c21bdd8824443558e35d6e35b562bfa1dff19bf8bc6ecc79a27380bab53c3615129c019e96de3fe397f28d182d4b7e2e51d8a6f1211fd41d9c55a29d2f06fd76ffe99bf6102047723efec010aa5af70bbfb1548a8bda5209d16e369ee0b6acdd896a3dbf6e0291d936b3fda9d63af97a28dc850e972b4122736a8f4a565a682f1a17ef145a594479524c9edad5cbe4d266f40916a320ff7029837e81bddc32ffefe89b0093ca5963cfc44119f6b12629bc9646d65e3b150de212c70de1b90c472651205bf86c7d6a8e4b2d1c76d58882f67452d8073498737df077d82014e88c407dfc3eb8fb01103a8bd5a74ca043def8f6289e068517a03bd6f2966d4166e477b3cf9c6d5541a9122c3ec8b828ec2d0fe44a596b8802527efb7afbb202733de15a18893375e126d5b9eeef44c49a1570d8bf28d11e9ef4000b6a5ccf598dc40e181367687525d091441f4b34219b30c42a96bbf445292e79b416052b84f7128ba1d2907125e14b79347b1ecbf489229da73416948026dc192cab0e0ae5ef87df0e186e7903e1fb1362e09b4ea8d6a0af7d8568604cd8fb9caf4db922bf8a4cb77d93eb3c7d4cff15eb81761f030328eb604ec9c7b9ba7988d3f5280bb96b8757;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hbb0997064f3795c04471dd9d4b0053f65cb520628ecfd1e9de72fff0015220570b330685bf0abb3a8c5d155b2e3b3f957c3a57114d7f75f2ba49f254ed7ea3102526cec9ac7062d9372483f0e8f75b9589e5eb345dfd33d6698062f676eb104833e520c03e51d8edffb7fadbe2b7304be0b86a9203db725ff14dd159b797b43625b87435d509867b1e9aa46ca03317b572fd693656ac77b23e1da434a55bd5a678ac3fa66ccc7954b9f52f5c5b3d67a34c789751ba6ae4949a7d544bad2c8a7be8dde68b08fb9944f66f232ac0a3f6ec37406b1d9be911428db4ab7e8e66a810a27ec1e8217ef02ca02a3978ed644fc135f1100c7cc386131b492a9074d71ab6f401dea433f62100e64baedf345e9df37456431b6a510543146d0b420fa5c0ff338b881010eb80cea0e2c09872908431f80a6099e8f732c496dd7da3891acf6c82d96126ce756a29d9c5ec9e2321fdca155509af0bcbdec1f0e773296c570c8370900ff5dce7b4b4c41d2f01210a959a8b5479da02c7037e8fe4adac36f46393c0a4157b8fe07dcf4c02d20374e24f4f4afce4978785aa5b9b0c27bb1b621d99d5406acef985af8f8512e7d1aa809a85467c9152b8f0e6971f9464c9467daa3cbd0fbf1c152931cbcd3f332bf67e36a1435fcc3f2276b109d8bf58fa14f84c6ce35789d0ffc0973c49180ff59c987f7f656f27d9e35d66ea0f8e1dd7431f4a8f0946b426b184cfc7dbe472050859d7069ec8f80a9417b8c3eea8f184967bca3d07fbecbb6e65734dc0ef7de05a07baa5f86d4aeea303bf62233d89766602d0d7b319e092ead85e3d49fcf673ac493cea69377f0cf560f5c158e39556666558d9845bfbd35dd7c19f71ba3ef7808d343713edac520027b9659a44ed9a76a288e71214beb5a849975bdb2b627b19ba2159061280691884ce00537596cf222bd53775514e849adcd9012606b46fdd32e27692f7e37d21e4925abfb9202c81df5002f3d8cc64957390fe7db2efca3e490dfd31c586699c1e7d1d130f0038a3ae5bcf224d1325f07014f524e62b07ccbbf8a8b97c679ec1eddbefdcb1fcb3f2f50d29b835968f79c284e942acdcfee89714a03617c0cd6004d9c8d12c2d6b38bdc9b58905b6e6c244d393e71fd0aafbcc91315414ddb089a0abe60d089e7199dc82fee473aa1873b227884ef2f6af0c980d5e50a8ebdcca9167940ae35ba9dde59553dad850cda4661881a1202daa6499dd4a0ce3da449f9e7f0cc9a83597f19760487b9b8feb3a4a0b61926dd3a6105e750d26b97bf8f5bc59e51df8c708d2ba0a027a73fb90e8fe99bfe768b69879e6d0a0f9f9899d93b9acd4df99a6c825177d216455cb3c851cf30829cf1ba0451bd6b7bdaff70d5c597703abbfffadcacd950816ae9dd7262a6cf63e48855a6ef75136e6c88e44a1a490a88142ffc752359280d5c1b48286035bddcaabe89f42b0d7f89565a779055e8df573dc32ee2f036e91dfb87b5679b83723d8af13cf43c50604e709b0b78f0be8449625bcc07a4095cb0f06ae31dd00d36ab4dd76b4fb6f6062ae2f85c12d9d738b39d4190db01b0d0e6bffe4336701a5f181c07b89b1b66d7a559a8ab96500408437e2f356cc703c5bc2c83599ba01c36a7b9b8be2b14834c9d644c2c0296d1c8246a5cc6d1d321d1e3b09112deaa72a052595e7047d054e3ad04a0450840564457c1ec967a32ee6e3ea7257a1fe8d89376ce501f9605abf9d6f8cbfec94dd8045fa2c7c31523e14360032eae48aa01ed8851118550e7c6589daba035c136f9ec296c66fa7a9add678f595b6684ba607905c5dcc6134bea874;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'ha19f2ffe30293516c30dab846cfd5d51cbb582f51049cab646664aac0ef8e16d58a90784de77636ff3841dd4008a37b9e34ea44cd5f765af8ed78f61a4b667f94ed08c53c762235ece15246e926d55108f8372b96bf0ad57e43cba0727509a2ac765748c99e117f8daa416cc12cda7788b4e440dd8e91edac6f2da5bf0a148d4b9522bce7e40f468acbd3c28eefd1322cc010752174ebaa9cc39d464d596b6d8339b3c3c8a28b9ef624adfc0a1f508b593946d18fb900f440ce5cf948ef10ec3ca47b4340f8c18e204e840252e7aa5c369b234f2a71802d40b3da2126a5c141ad2707b2168b8531e8aa53b208854e0c3f57a877c13589b9cd18f851997144d265dec431c4f5879664490f8e97e8b3f3f11e6c73e49cb086c5239db442cef548f7a33d3deb98f9da442354abc8f89f9b45638a241542e95482fbcf4ad4fb37ceb597b7a6ed37fb1b2a906941b6680a193337cb51243b79ce8ee513cb277e70c7ffa4b955f7384a880426522e11529fb7f15c9b3406eea3f122b1ee0bede18e3d7df73561013674f8a65d5f04ece8a46b049ca9f616d7856e619852b4422eab5e34594b0092f5b37aca22ef87c17e5824001bbbe847edb0388d234d986b8c1f395de8cab8040a25e6085bdd7c48428665ab30f74fe309e4110a74991b9808b0cbcd983004b24877f67066b4715eff8ddac05447bcc6f7e86620ee4d33cf11e06d0feb0d7fd95d2162ab886689b12d3f9522f03839ce6fd5f71764370c917cb315706971b2f681560722a6003df2a219db749298055a52bae3a6b071c57d242de09a95687a257f83a382cbe760580cab0ac7c3b7533e21b0fe7499994ff2433043f01972b4a74e3cbb802f1a968292bc1067f5e45e0dbd0bbc371a1c624c2374bb33fb14bac56dd06cf325b3d5ba1e21caa610f6ddcf17385f371b8eb03b2b169af2aae45d54e3d3fb76a1e8bd0ca2829fc271cfd135179fdfb926483174dc176614b69d30d762744e8801f45bcdbe088f8c4a024fd28767a52992ecb5b810c1303026db3b3ce887357975ba845b2d32d5c0679c5db8d71b3cd0015aef34394a795ea64a49ea9e2c9b7187e4d27142e30f3cf89211691e07ce64644c0dc3a7b804718e97c9418f8107c1040c22ab7497c89efd3a23c0630bc4d64c487236f2b1c08e3f4964d3ed629d7dbf6ed26a06e6ad09248ddb7bf7f89683e18ce271e27583263e6afe104ad48d30cd0714bc0b0a6ca38a6b6ec1764a576398e740b731739114bd90c8dc5ec0416569688366177d0b48e781bb6c17f76f013e6b135ea0af9aa2ef37f45a54ffcf11434ccddda7e4f183b059c7fb0acab90031f6c2ce2a37ca3ee44675f4c4cf2b3187f9fba214e6f7cb796dca1a9238e9336fb4030423f615de54854303bcd293d168835e9453ce42159ddd4d3a7a7481ecb14a485118293fe393b84db738cdaa1cdad475ab2bef7093b0ee1d9ba8fe72bc23cc1f3189244b5f37b36854bed6592f648f1894ee91d57b8c40f4e21c86872ac664550b72ca23181ceadb949567a5972e04cec6ccaa649671250e9f081e3372a9129440f631c91992ffe5cbc6a2484877b65d2b71df840a0aa370efb5625fb15f9014d0853a2586b2cf895fed351771273579d210f9493cea6f4111c01f6db0205d5f403045562fcda8deba3ccb4bc88a475fa7cde19bac971460e4cae6c0846c97fd95e9263e5b0ca7fa0ac1ea395319f14b08213179c5926d6e5a60bc905dd91fe25ac0da9e0dc38ba89a3ff878a38586fc615ce861405be349e9c3c3c60449bcd65e006895c5c34821c475ecc23f4ac18f7b02ad058;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h9f6921c1bb5e2a9839d74281f9955b9cf1c8e66bd16f94646fea6a9dbcb1ada00011e724b9debaa2a822f4e711340cc1e447486a6ac67029da19d26a5dce465b4e8785e13574fbbb591b1bb677f71cc58cc51f3aa5496054adc7f699566a806888fe70d85990b8c2181db6034cfbfc15ac39ee75aed929e8797f1398cc14c884934e9d80f54fc1e7d832ae1f6b64ee2a62956d7ac8835cb2df1c7b5b6599bcb76abc9fc01690f76e35e30f24e4f3c8a552e369c0b11f79ec777ab5763bac8120d765bfcd96678fa3c0b780b1077d98ad58d68b9816c52276b850714963bfb2df056cacabe66023e9ce9012b2dc251cc297574709fe03996ebd18a6e81dc70af9bbe48df184fc5ee5ca703f3d3592c4df6e421078d38a98c5246fa50a59301c7be88936af7ca7e12f4eb9a548a476a3d4f9bc1d5aa9d8e36f95e573d55ce81e97718f12f0e504a5d8c3d23be798771d1fc49591a932168d2151ddd7d2cb6f8ecde6361bdfeb7cd2a27e11a53bd1aad27229d4a9c944ab743ed5081caf53168696f44887b4cd69b4c431789429b0623ec5e782ba3325a1a5158dea8eb95fcb8ae245c0ef6d210c0f2570bfa1328303dde8663fbf104dd2207903e461cb4fa027f1ca82f0b08172e19ecdd2bee43e89b29165a3d74ffba28be1e6c9b3d631059153b4b6bf754f4130666d4388d964cb4590d488f7a2eabe292adafd5e25672e150bd7f914bcd81a84ec1a9ab45088d556b8b62ebc04ec3e2f2a7cbf0918fe226dabf3e010f7d71ece0155d530d459aa66e89c337fd92a0764f1bac1e5e5e6e1e17ec1bd7cd0d6dbcf268eb30228c6b644ff1bcf9d4db2098409065472bdb4d2ce5889e2855eb0c3c54bb00179133f77fc4d1a0813369fbe45f91166ba3e194ce376ecc4ee762d1fbe89360e624e89d7ed3e6cae87a2cf5a93fd328e9622d496b17db9e5624a8484bfce039429d44fcf280dd6f726554b369d52937977016a221aaa4c17a7a0d1b77a3af3321c048cf4962090f8d98dd276f52b2f9d96691a9d1b4f6f1c27bc7f98f00305ce76902ab4c226513d1f960ae1e3843133c65ccd6d46bfbb8a70b13a8b2501d35ccfe7b44b0dcd03bfec286dcae1fcf329dd85738549b5c8caa3fb354e0f74775f0816a0ff038499d8087445c47f562edc6111ef46a757da5c19ee220ad02591cdd697ffdad677f477718b296dc77c08a9b8fa83a2d9cb5dbb659ae3d3fcaab1c7adaf5dd49822c8fbbc92f156226060b05c6effdd2807d9fa98dd40338757a5ddb8e17ba377365f45740aa9d3e45e2259a7c2c905157be56a72fa26ea7926f1e991ad27365cf7ccd3480774e097d684a69897167b7cfff581375000361a0059ac0011af46bb08c41d1f7740b3b6104312464ef1489d34c6948b891608b465f5a2f80150a6ab4300154423defcc73428982281e4bdf093a72c97f6bdc74d4861e23ff570febe77ce6c5abcb58d05900adec25ad24ad7b426c3cfb1e4b52abc57f9fba099a33feeadf3ef95ad1f3b712ad0ed1eb3a37953ee7dbd0178a39bccbb7ea8b131424018c2519b2af842baf38bc26c683a166be8c219eb7ae9e1314972fdb06092b5f06436ca3bf00f7a70ffa3786558e6e687d033939500c7412970bf83acc145adb15e1798d109943e2430c1348052406d2f01f0c4727634ad015e8752871497ee8cef69ce0b63030988123c4b9a801a60486d4ae99eec68f8fbb5b6c616d375da97a5b49f749031d70160017051c03948130f7ef987d7cabaa5e06e38f209d7f80889275765950d76401af01dc9ec2bc9655f786f8be037e8b119360c8fb3866213b1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'he6fa3ee32bfa809ed00c1b8d08aa0a1dcb0d107cd7d970aa574bb214f2bd82bc1374364486b330289c7a19d6283c0d74d70d3bbb2dbe885ee294e7a8e57ce385551e8969bf2c60912f73e51ee511361ad9a4ae9f8deb3858a4dc6044a9c2a0cf6c3ae73df3da09df9ea1a8ef551d572737f3f58d936e8a055499faa2443b441773897bb15b48affbe31c82e13a1b0cfefc1711e85db766231fb36efc3c803163d3bd8a98059784b839d2c693b140f0855663bafe7d60c3db3fcd882a25c99fae176b6b573c674718bbfb747a9b585ebfb44d1e1cb8d2b2a33c04bc98d1042734dcb1abc97cf16fdb202643dc7e8c310859685134e5b8ae17763ce7f416e7b2795290697080435aab925c802613b82a4648531006098ccbb2d35b0a86cf30a51dd7908224312a15a8813af72b0760287d186e6150a94fce24616b835f00dcccf9aee7c05309cc27e739cceab943975b1dddb68008e16d2972c964d70c4891d5da9f6b9092c3f6a709c21779746d3854a0742bb11701e5f6aa0d07ddf24018f355badf2ccdbb44f7556cef479fb7c8a8e3b6afe87d483e9717f12735b842012bb79e0ad2926c1a5d8451439654cfba4633548abfe8fd50b061342a96f2637e3437d95aaa07b9f7f3684d35c6c8e28b6a5e70df245299986bc89f6a31f8b34e0be9271ddcd36aa5bbf96731b025534b4068ed3184dcc0a83f0160c8a856e62ea48b2ad49d09cd6bbf7f98581f7507a5a9d08f539f220f9de3a415e2b43a87eae9729234c08741a8563de43a2f1b7916602d78659feb5c4662179e28e1ac32ada45b34b300e43ec42da96c9e5a68679a696f731ba374062e00d11582be1043de110b25f5fd8192cb9ed0ef6c097c2ebf1c037c106f7b26bbcd75a7ad998194c0834b191b2d63748ce8cf399700eec5a503c52bab475732b6927ae1ff6fff872bf7c4db57eff09bf254ba0eb5132e1d1e359febf6715cecc56bbe68bb78ba9426d888fefd94d5e66c17cf738e563d3cd6cd8026d89bca92b678471c84e088319a634b499e57163c56de7b5e88119632da92ce97fd4fd7894fb9394f4e08a239f14c1f5c9eaedb9145178c8677c304f1d3c6ca0e65ef3374b118e40e51f6dce1ee42f1369bef60818c64e3335614f4f4f5f1351b6a43f2605a95927a8fa01253ac0db802f40f99a652972eefaf75b33fea64dd049559b95754079e6b3840f16bebde594ece9c816720c24ae548f0056f4a4330cce893f25e2c24642326d89ddb8e4f7bc251487c9c0d6a8d7b1111e365cb7d4f98a2bdc2a9f89c31d038cc51b7fca10947de6e91ab585ebb47064a9e7cdd689f31904c491c550d8f3cd73ecd66905a12b19201f2f945c061adc8eb8ff7ce41979f18deaef84a76f0ca6b6da707f23b3f6434fcb94eb019abf57cf151b0189d2dad732f21875e3a2dff11c3569a4ba97d6c16cc23b5d03d2202603dd12e289fcb8fb42f17bc63ff70868d16bd581357716c319cb6863a9363b21a97b929cfb0525a310031619a9bcdb74702e4c4c09295c55c94db7175343a5faba0a942344161c5f9ac7917be8fc7d58bbc16948f898ec8e7e5fea17be586494ddbe65f6286dd0c4c395ffdd99e3f4d32bac700b9151d34cd8a1a962f8abf82795ce6a94c2da53b6f92e12f39997e5688839ac153d8e6d5b6d8a9e787454aed536ebbc85d9852631a2e9f7bdb304c7f8f1aea3310c6a1bc7836a71c7e57b17efd4395b3ba7235afb57025874b2380d9622588fdbdf8bf3766ee1909719bc8bd04fe989bf2e4dcf5b769497b636b951b366d212275b447ff5e5bbd1adf2d0d277ddb8722e3f4e4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3aac5e941d3ddd7aecc5b682b5f3a25f6d6b30fe0d143d7e835f69a330025794a9ebaabf8229554e20fc72e21ae27629e0be6769744a57593f73142df2e8c8227f10217427ed1e4f40090caa0a6b9e49db95f7c1a462bd947d40ce45600243914c879c5fca9c443e479cf555d2e42260a55fde0bab5c1f56b79fd3ad2df835336ea89b2c58071e5872132717a2579bd612c4c5541122457b4cbff855dffca0b9af22736031c14ec44c1550e221c966fa9d697deda955f827a29da937aa2ccc1801ce67e2c9148da324a8ccfcddcc3948181d9b55c9640aa3e793f9a798487cca5f4bf6238399d25cf84e12ac8872a8cadcb6104c0bd14862272d27668a76d737929bcc8f807c11beb58fb4c9541208bc5c67fb604c179743d7e915af77c880ad2b0a45d474d8dae8fbdb2b2045f5332bd4329efface67f6bc2be104d23f06c473d70a8121b84366d649eeee679b91ba9aeb0b7f493a7a8478ac86069a855c88e0dd7596f07d5193d4567a23c4abd868fc0552637c9cc664506bd4426fbfb5a440e5b28bb108e84c1f042048e7ce3c10a84d408b139e5c2bd9760b805ef885e2ddf20b9bdfa9418793899d2ff3be11eef37da19c25342a3a78265a7094cd23a124d72b3f0102766f92b2f0e7a5949974ff0806c2e7403a387ec9013e01d7887d7c507c70051e30db87a160333f0ecc76297baa566a38d6c25695cfbc707685234e88ef6c22b2a6f0671117cb591c2484e23b25aecf24bb9e9681b650c31893447960618053f1332d9c46320379223a95389a7ec52e32e8aadffde32cd021f36ce119f71e888eae87e9a99e6fa7f86b83b92a79b700beafefd4e371cfa5b9c3e48762c9f35d3f2271c3b6b37c5a9c440e4ae0be0e7879a93bbaefec680aa773267acd86372b06c4afa86c3d3e93ac2506a1a9e5bbc58e002ec26564df1b796a028c1d99626dc34bbf987d089d6a0520177ecce7aec84dd161fbf122ecfb0f3862bae7720df09f94082709f58f7de910db45cba7646dfa0af3befa624e418da88644cc5a3595e206e5cca290cb97684746a9fbae6a7736f020191429f337e9407a07675be35ff72ff4464e10248a8d9e9f13e82ddcc23385860e897c644007952034a3019d938eaa3f643088948667aa8ee3a1a73a3e42d6ea0300814dc344a3f1ea545ecdd8920bee216df78f767c03540a60b8a5966ba5d4726be2866fc25889517807f2fd0bab76368a43d21d6220636e0c275445f02a33601f12ce2c8aedf65a50f3ff840ecd42115fcc9090617471792bb1e7c3cbec81865931f75bb4128bbd69a8a1d693bbbdec14359efddc8eef36086ebc766bc9f1f8d0272dcc9c5906b91ab00b0b9893ced488145acda0f777481ca1cfecbcce3fc62fe7fd8918a60a2722a3c2aa6275c3dba9b8d71941e22cb58f17bfec109bb9e9c044736ed00912cbc296cccf015eb94521bb65416cea7d2517bbe64053bc114dd564c5359b3eb02a13293520c6a425401e3d94ba0de880ef3a87098db7af99d3232f0da4136ec9ed5b9f5b444c597c758a98142b0f98ebe4bab203c748e906ab63f716d9a60c91e6b4f944ad00d4d707a88514be9b46c3ac6d655cd134833e87f6d872db5b7eb918eabe8e635a4bef8994988878a9123aa4aac06cb6895ac6ebdbbd02de02143df0f2dfa3ed2566fea6f1a08aac6e8102df9a5bb52e622d23010f3906cf414c7ff9e2f2ad2b78fdc3c8587bd9de0ded4f23982236059964017f07d3ba3fe2ed72917942ca816738d9b1727482c2ca8b385e9a5635ced8c23e6c6d2ee7e5a82b11f3571d23b57536f09b381189a9c1ce9cb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8f8b74039c2c7ad0b884878bbb669e841ddccd93f85ea9d18ddcb775978ea2deedfa63c59d300c1f1848e15b7aa160dedcd0e133ee986c46e7e066c3175f94b7ea252d4595b61092607c99a5bd9bcca10e5ea924239536d5541054aa78922f5d0ba3a689543b576017adfed9dcb2a7bfb0903b65d4128c69c69e3b17cc8ef4a8b0782d0fe4f81b60c1dbeece7b8915f36e3d4129bdb2a9b33ec19a0d62f9781a4739e16374e298a35e2fd520ae365d04771795c84ec8d2f9b2ac9acf52040438edac5a0cfaf7addac48acd712f27c7d3dab8926ab9fcac49683443b0520c31915c103040e1428974dc0264c0b640c7f6fe2ea861357ccd7bbc9a0eeba06ea30bac0d47e42a78d2cd08071eb8f40aac2c6ea269d9a8710c9af3bacb63cfaa504f31f160ccb0dfec17980e43b52f01e4a400f8ee4220e8b7983b1167fc83e19b94c3dad514205b8011caa0f682692a35ab2efc4c07c0f420999078a512a090206b71fb3b1726888b520152adbd8f91f73423136c15438d5729fb9a7c7eabd7db18d1dc291e3af2a768ff6da5172021e690f259ca6f322ff2acd7ffd311caeb248fc9d7f36f6b9b17059d45989ba48889f148304fe609f4b4c0b6d7e97e1e40285bd7d03877fc6c2ce81c611d583d8d14f934e3ea15de23dd20d8ae5484cbd1010f62806e5c177758e9400c9b98d28fe7012a0527d42d05ebdb2a3db804a2c88e1192bf512aedda7a364a2aa0e25fdfc3062e20ca301001690467df2ab024080cfeb61e36c9c322b272fae1ad46ae67482fdcbc92419dccf620a562ca56154da652e554c8c8f7978542b3eaf0dc3b8f27704642182f8ac6d74a32c0d77bddca5b0ca2ff2f15b6e2ff22d7b554272a5ec6d09ad06f970b41aa2b7677286b8819bdda84946b9abcaae551523eaa4f4de4dfb33e30ec2624a2b7e04d544f4f290943c70d25b6ff8b2c898265389e39724daf2e53ff1ddedc545ce59afc3bd34230027117701e6c97bc21961c0f01821380f868c7eb710345eb95f6603f2219daa868b9c4bbd839dc91a96f130f0c662bd659441afd163a9cf5b6bba5ca0b43941a11d961dfb1067c562dab35ce4d4e60a2109aa355f03b43881caca9cb7d6cd4f9cd48093785ce37bab4107ee0a13d90dc8a86e3f0a1a593b7cff99b2f2351d36c779af6e3ae54d5a2551155c30881835d5f48850edb99f3f21a6519b595e8a7160c2402b3f628528c4f7222bb2da0a230aeb64b6d766045a5d59b943bb6c56f47e43adfd72d8838e3c8ef7b5d5140178702b62daad6f3deb5e513a0f181bdb396ed608112f67f2b5d6c392e9421b770aeb7ee3bcc4282979c41674db65aa282db186fdd453c6089391893370aac28359a3051e7368cece6a179c8a5e912f629626ac737112deb995424c1c384a9b6152f279711361045b9892035e0b8f6e6272a0a0674ef82a57f75b85b5a9200c8fa378449f12c5f52bb1e2a148adbbb5c038703db0f449c38ef77b029457d928404aacec0638b740c48a7a68f1e884261fae7f005021acfb7d955140a2e5079fdb223f085b5e90544028ffa31e883a0388bc243eb6ef0954b42e582634f7601631193dac6087f6f4d6acd502daf33a17fb8f63d0ca28c8ac3294bbace90e20e7a862c138c748d54f22172df9c1c0067a7cb1e38024ddb51acb8d32c4b837dc43ce90cbc03f875d75139b54095abad608b1dffac628909a95165bede2a439b529619b106b4270f7ab8be74ecba164bee98d967e70444c424aa09d87b8866d2b6c3c0a1c52c6548991d70adac46ed950b1f949c62190754d04ae436d9be2e0b852388954a96;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h9a40c3bb1fd3f98130859d006da8a8305d453da7e66aa4c8389bdb838c41f9bded88bf2c358a4d8dc4eaa3160a65a059ad2c7cf1b914230442b79eb13d80adabcb2915754f897350a0809722cc197a667b613118d182420e4b2cb92700b955fcc917c7a7b8ba13c5dfb1a8a532cdffecf53f29cb37e4822d54fa29623fdd02e586229ea8f90051f6c14661a852dea0a941d505e54c8db171fe83fb9fb2720d126ea11fbdc8ae96ae9c3c80eb1bbeb2c5c5e70322d45b92ed875b43ab5715857dd26b56f44ab18f29528e128f8f9961e4d14bbed6ab91bc668b146c884022a8f146211b0feb3a26d10e89c04dbb8fb918d33db3b84dbfbeab2b9cd13cf8e0417b87548f5898bba45512a86823abdae4913506b3058787b1b56d1112d4c268bf14ffc8b550b12333b4fe259743250c64c8ed197714e5ce2cb41b63b49a4f036bafcd869f7d83dee2fc429284df5a075e1dc8dea5b2002024e9b1982379d2e6441fded50c775476e88526042dd3e8b764aba7a7d85718b15501ccf1565652521634a17730278cf71f8f08f85e446e9fb23ffa5802ce876752b56f48ebb9d166cf36cec64d919b67ce85fe9a495487eee22f124370f2d7e5e89da6d33bf4f71cb59bde89f9631d07df05ecc20bb528b88d0123bec19aa9169912c2063ab686872f2cb3481b11df4d480e9b200d015126eb53cad59a152fb68abcd1fc79fc4dc28d13cf807a52f39d7eb20cd6a05025758b1d03b1991134420a56398ef8b4845469d6595aaa304d7c6591a93ab1a1dc2fbbd2d0791db2c05f390ae8e0660e5d9d1baadf196d2b17f19845e87e38b354b801cfd56eaaf24dba6777b7f66be5b2e21f0080c1d141fae363164cd6e006308029f10a1c147caf474e33e18a3f37635f4a93a4b9122522eb5d73bd2d7411fc8a0637f11f8b3e7e2498123e23dedb944c30a05c4b64f078328580af9102350e92f1dd3c025643b7814947778018662aaf9edcd90d0d6c82d731c0de82e46f38f0d72cfe9862070d71fd2e4294eb86a5296c2ae9f138c2697cffcd1a976b7bbf7992f72cb4f22cd5c2aeb1c0bad77bd0422c6dbd74b0749fa0de80d03dcc634a5b69ccd60d2eebca39d21ef35740c822a7ecb950ec5704a25b1b070cef8ab0462d9da469c32136ffcf80d10e115939639fb87bade679c0e08428f86537fbe30b10aa2525e473d51cfbc301444535010c12b35d4783915cc15f0c65bd14d4a865dc5776839d5d99ff925e47ea75796abfdba53865f478282294059558eeca8e3d5095f4e5b53518e09db36d32e2482768f2775f3b9ecbce67b058d4f2dc5caa181291c6a23efa3019a8d7018fd4c40bb0d7abd5b8fcfd930b2ef8919c49c6b04b340650a993b2fa3dd52e06831b2a557309b8db50b443b29da008e8bc4d735f48968258920f0466adfad4ba0a0338b15ea04682552e7b006d3ec69826cd1d195be294020a8d76b15b230b965ced6598fbf481d9381c2ebf0baed2c8d3c963d689ac2cbe89d35d7cfb39fde910dd059ee95ba5adf7b23f516865d2fab82f679488efb43da2e3299fa084621cdcad424266e9e3fbca4a5d1b770bb5d8a8752c9927bbfff8a1185a9a8984937042278fd2eae43b03ea3d93494626dc40362dbd7bebfd057a2b5ccfe7d2a42e82d86afd39b9dc559d103a17622884e3693ed1c98eab582f715df450917a038edf194547cda08a434cada01c84691c414b8077ee72183ab154d83cee868b4cf4f560624f9aa92f74897c234212e680ac96e72e62f55f52f43456d29ddaf9b6ff62b6caf676ff3cd3ed8969b4204787194b4270a16a1f59a59;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h98be0b0b6e6d73df54355c4c7bb5353030f75e3a1c146ab3eff7ca40ef386af1b78f5a38abd60145b99f44d16adbba5eee90d66e2cb25c1068a0ac8bf6238dda708097504d94e9af4d2533c8a079c5760d97bc0d5640f6d9578a0290c5b2b4056ef2848a17580c107553ede1df933c86b74ec0080b99b7fa198d1594b889b0614a31eb51a892c69f71eb736f9c729fdc14a4c862bef64c51492311dade0d94b1122d4e4a119a6ce7ff59a1754b9c3ee152a3d1eb4a6b9765f0b7b3b1c450a65a8104902df7252d14cbebbb83d8865bc7187e995253f9c361b0ab27feead7a2540bc8c7cfcbb90bf9dcd4bc7eac8fbd7c78d418e04a64d6cb14e57ae23ba0a106b93ea17faba3aa0d5ee7421c2212ddf1e68f699d8d32e378ff5304d77acedee917d95fdc213a8686d19f9f73a7a4c0d967e190a06cebd551b2793f4f7237a469502e20845daea575f3c4ed44796794595bdaf6a9c43fa85710dbb4c4d6ec356da22f6b1bce9cf6cd941ae1f7e9a73c82f6e7ad65cfefa7d4a39dc366450ff5d8fabf199f2ad663d3c2dc6e579f5fc8e6baed0554fb5de69d3e685222d65308c3da0a389bac3f1363b2dea49d8979c10f987db7f7d1b39bab24b60da0f269a31f21852020b93a6301349064e8699bdda56f0d15e58d42055d27ca364dbdb6ca1003d79cc83e1ce6829a5b10a1a348885b18daa11c954668c6a4b5cedeb9c6f42c56ad6f7ab77216d6444650e1e98f64d15749645f71dcaa01345c55215cd967a4b13949e20cae682170f062ae1011bc9cac72f13cf897fd88bdce926ff2079076c53c4037d65f86a259b9a48bb23ebd5991007cf83cccc4a958a81b8fdc2cc88ef6fce4076a7f32973d9833f56ca9c2611f174676d4cf87dbaf47c61c3cf9a3b196c672b1f3d7df76944df0d855468899fbd8338afee48b33b2d5ad2944ba782dde3e0daaa667a0936efab315d07a5445eda0fda6c39db2ba8f837ed96aac8e5d39fb895f148bff56fee71fc92096757e5209d9fe8a76231df82a88d5394acf02a1ea94fa9cfcc3aa82d57ec62f299a0d72c5f9d6da754fa0caac5a318cde7c8f0615add131c204f5243299d5866e9d7fb9bfa073367a082f19f8472f52727871da0e0272199fc3a0ff1b94aed7dec198c4cf19c32e86ce40276478f95226925dc86f44e31a240f918ba638f14ec77d8753d19d4dfc74e2ccc1e03cd0452b4ea0efeb8eb0139f4dd381f546a5d36f7ab3eae9be19b7a2bfc80348bc5641e3ef397a3b2087c0e644584a244cff7737867b5e3be6b393fb250d3dc8f0bd30ae14d556a729204b3d9fc3f4be497f0439a1e6c332fb2755f32aa0b7b0286cfb4625e6716ca39b19bf35a67602617893269ad9aa6709eaa949e5abae22c600b4f2363a99238a3c73387793dd0f8b7507fe45bf36b13375ebdfa5d8eb98f764fe46d7308fdc29ab13c0ea94d48d5ebeee1018ba39afadb449f91d3e663dee6d5ef64438e23b5d736be9317eb28083ef2f5f03354caa02d222b69818133b4b352bafae6df451c1135917a75b6a3cb5bfabc9c0ad702e8d409f511f433e064501536c21f9282cf327ab1229ca5a59eb9afa5d01ddf6084b7e173c76ac1ddf27182a7003f441298f576c51f12f3d35bb062ce61f128b9a5bab1c650cf9966219c42ae7f0ea44b1e0eedd7ebf7dfd60a5d0d7068b149e794185606f694a8ade8314bd0256f4fa0f8a599727ea080ba7c6598c7acf2524d52c597bb95e1536e6a5ed2196a3d3182cdeccc3609b55c79af0cb44525fa3f8dd46c338f7797f63b59572f5d1487b8475191f5105c37a451b6e66431fb57c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hf706a59447ea41694e27cf514f0599e7767b8b54f90e30386ba1ee965e8ed33e7b92854e324113bcce3c747360a9ca59b3a7d358a2f532e7247bb0a098e091f9c83a101da4d8a2d9edccb43f5899e39928b97d4ac8570b29df1b5f2b9522cd380c3d9f456cd200ea18b6d6275cb5570bec2d7e11f076582ba3e19e5f07be9a80b9ecf1b12cb74bdd848c842ad802b5a1a2676c0aa7f48b4a12208d9ac0cb5000727fe3eeeb9d8efce2c65a9e314b77d04d0e5c91e5dfa5c2ecbfa99456d178fa9396be68dee57cb0431370bdb1fbe448c980458d6157c6e616f45135deb2059e0e6bcc65ab12cec95579798d547f00c076efdb62bf09ff536476d3ab967ec13f81ea8544508d16ca6183c46cd355a09ca3cfe3487384230c8f5cc4648e478c76fca20cc830fe0acfc7142d26fee28020649e9749a5df98848bdc02b69bca01914b2bbdfa6d4572040126b16bbee21c33b68630dc74a5340a48889ae5726e6deba1fc4f013e1469b9fc027288aa1a8cb2d6b14e6e6d803fcdead478ffd713336f2f9ace0dd1ed63c6f85286810bbb17e82583704344d2e9f550d39b1e0c8d8e1a05c1e4018b7a3c6c7928cd77a3e6db7bf5ef4d0cb615234180b96781e0f3715169b9b2fa43d9d6979f20328f3c9946b828da8c9c55c5cd7488faed8cf3c0eb1d07bfe11124a4d05428f70a25844a0323b7115b61cedb33b41e73f9bc32f1b9452d1c24aa847afef745e28ad9004b56c16fcd0250ba0536b87c7af5e391eff943e359f611cbcd19c979c69134145c058f8daac878e9dfb6bf6389e1d76b97cbf37bbd05ab5d9c80cea8731b576db300315f8b6637591a2e30b6c351454adfcc4385dc5f2eabebef50ce087dfb3035d0117ae3c0290cd8b1bde62959404ae001508e717db13905901ec05232456bdf57d1ec558f4aa5425fde07bd2db5d5e8cdc90cd658ce7b97818b982a357dab94221dd04889819a52120db992538b7e4e6b4d55eef4d186b3cb10e9238a4f53c0d05e2b89679bdba56dd131b46fd3764a1aa8c127765eb6f48168bd131d30497f6b0e6b0e2170683a1a43ef1fd3ffd21ca08660f9fdb30501f1c4a2d3655486522dc321d0508692ac87af295dd46dda345e6cc3229e5c0ff672613f3d6d37ae55be98454c55a105d7811b32a22cf3680a6a49de5401c30eff121a3433b966f1d6d61cc65436215f073b62e097058dbe0e371b6a6edb290bdad759469373c750d35a6123c16b1d58424f3f0220a0471fadacad641636e3d22bc017bd16670375333d14c271ff6c0c5f48029cbe61e1a04b73808c287cab3aedc1610318a6b2415a90edc405a1b954c84c3192014a4e3a7bb005cae910bb5aa107fc915b8711e4c9c7be5306b5b5bb1af5b999adedbc10bb250c99f6c406c363c4b4b15b9632ebb5847ef391b9276ce27ee377b13acdf9ac5d673518ea18f5b2fe2936413f71473b129a0226d3cf982e4350e4b83e5610afdf6dfe8014464e779addc222da5ad7957fe5d226bd85c7f5bae09c86c8876c57a5eddb7521c955c2f575aaadca80a89768b03479ffe19dce8eb9b80d8500012aeaabce396cfa55e843056723680cc3e9071743424c38dfd8a0e18d17afc67c2b9f16740db071a6c648479ee6d10022bafc25795f901db7389f6a53ec2d7aa6e1223dd09667f0ef75a2de85b23fb471af93980e7f29da69e9e7e61f54f9a1f37e2005248f40fe050a2de13d672590c1c6facc6941f41842c25144b7768d0b0418811827717bcff4cf14e9dee2f767c127c75ae40eb00f37d9d760ce86bb93f1500f67743e8823a6ca39524f8ece9584b81522;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h26beeb125e72716ecec84cb7f6af297829de0d4588771df410bd5829cab89492204721735c3165921e0c3c7a7bd21287bc574eaa22c48ea3a8369dcf52c4eda46f2573ea4e54540d105648eb099ad1054f83a99eab4e626fa0495f7b25c51df1bbcbb26ea4ae7e24af54e635ade4df6815d2524a6dbfa635d0351c259463c20911068a088b8112a9ba5add8ebcfd4970d75407b6654492777062bb562a3fe203fc603c41c84dbb5129cecc5e401bef25df3da3ca2c9a5d7535d3c1dae1a2c73c3b12fbef67b1be3cf8c913f359e79e72b00c8974539424169e582e950ae71a9306fc22ca826ba8e7e1a79b1e8adb39fde628123c1f0c3fd84fe168e8b59c6344fa7369502a7956f5bb0b99ebf9a96f498e32c074d76d696a92daa0e95c9dd811704d2d73b49f701eac2cbfb92ef31bde0c18f36a95b9f10bf90b043a392e54ea7b7394e0a5912de30d28829568f1dd73553213930f514a68c215aa4c088c5c4699a8faeb7d469a8b992d79c5a5ccb69a6654d46e78e2a09595284791688e8cfa7a88da0dbdaf03b47c0226b1ca54c7934020bbb4f1f2f399270072db74d083e3afa1d52a1301c8bc921a5a5e82bf2404ae0e30f094c107901bbe3c5e4ef54c08175df18c5451462cea392d766ef480d3f2fa89c718088d854682fd717fb9dbbcaa15a1bfd469bda3626e725cbe01ebc6ab0697f8d966b446f7b33667cc639b1953355ecfd23b38745985f789852c42f72b8fff95d48ffa17c6f7f0c6c5da233535a5d711423173b8aa485b61bb453eaa0090356c8f201dac1313f837ac85ec4e778fbd1e69db2527c77771e73226719726367c36e40347edadbbd9ceae453b7eeaa80d2969b48766e1b07ab4bcedb75730023dd68bf86bd946ce54b35303e89ef762649c4807d73af1e2058fdbaf3a9d669165e4ccd469fcb3d91f01a00f72fed18e7b462b0fbeaa6ff936ec62747ad1158ead5a403f6fa53ccb697eef718a731a6bf2df3c2ab2b2f3b1781719a2baa82b9b2fc085d7dd3eb8b0af341ad2c38ee07f51ac105ed2c1b1c39c892870d2e946ae386ba6fbe0e66d1f8b28ae6b54899ffe1f70ec6c987eb205bd2b34616ef7da830a30340444928c725ed2c1dc4f18c3b79ee0b9c26195575d5214e3378daf9c4dc15d778eb710d0620e029fb147dfa4320e634f2b1408673750b8a029456232dcbbb3cd223c6643070f48cfc660877458d6331ff8c0decee945d15f1ed8d971b519774fd76de84822d696a93c3d0a1d7d62ae1201e591129e047c3cd1d6e5e6f4113fa1f3265206c35be4e04b5d1a84a9f16791d25c952b406734bb568293294510d1ee9ee77ae616680c60391c5ae1adfbf633c226fb37cac1c36516d180a9bc27f7fb6da2eabfa6e108d6b91200a9b217893cf77bc27c183bf65a646c77ebf376f531ef3795f7af432124f7fb213baf6751605725da8bd14d267363c9cafc706f820614628b41ce991110969ad737641e24449f5e1d7d3df1a61dac62ac2055d2c612330e08afe2182afabde74f5320d29bc1d5526f385ca3bef11ac889a0b0d8c54b37d0b15d719d4c6e441ecc8d3f33ef60c4194ae09e0220ec1587fe37c051b6309950b0314b6bfe4420956a34e932a23cd5cd0c06ac59ed53a10bd246837dcb7f6935eac41a004cf3d23e45af83b0c0c3c8766737b385f2842a5a1c3f53f0230bf25920ae507ac06faf76a97465a4c933a379e3763dac811b45f7ab8473d57170c949ddca30fa1d1bb1f978a2d68125e4388861c154ad5349796d3fc2425e6736ae7c52256a4862ed042f88d8bfbe594413b16c8f1c10812caca29e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8f9c4991258618058e77ba2fcd5de040e8e743175bf8e813857bbf183679054611b625bca5403d0c23241971f8c4b53a15aee094b83a03ef201edc3d10cc78bc79e1227372f5b860cdee386600ac560f37fbf739b3645443263b5434d82b98d78b8399bbd1fe457a95fd1f1b3a23c218e2cfc6e5306486f6f2541ebf1cd3b99560ef5424c9e8aa1633dc29b57674dd5ceb76979735cc2c3bfbc3e25a0fa7f19058578a91aed1bf1a0cc71ff7d728767c363663aad064548cf4765ecf98b3e8caef991a3d388704da771cd8448d7b03542456ca5999097cbb4c865111a0f2d70470de061c6e026908a5c3918b929d13e17971a616b9bacaa8e9b213536d9d3942007f46dbb97dfe1542985b70f8c22458870e931b998a36fc7e8c769742f4dbec298a9d5e9386f7fd1fad5832af6cf0d0769f962f095a9055f2cf005ada5bcb3649c2d1d819dc53b9ee135fde777c071b7c01551c61548b3e5d5d5d8f169c29e9e0974c7df4049b83e6d10eafacb79ee45cfc27b3afd5703f1f72b67d491f1a2965891726abacb96807566d5b2e04d9cad903763d73d8cbdd00a6e99ecd44874619090b345c4e914f997a644d2c95376a303e235592a138ca3659e0655610e068bc3e649c53546d2a8911fb968660dd769341563017399069102be06e67749c0089a04e172260f8f443aa07e35abb7b944d00ed779c4a8a0934c6910cc2b459a621c64c798ae84abef47e198a6d4da5e2808e25abcfd3842cb967057b1e760940b35b3dfa4f12115f18050de7658e616b04021c5d1f4556d821165d0f792f23cd6385cc4428862b6541740289183cb96951b428522587d02f6cb58302c425b3e8556249938864cd23c61f41071f5914549d08b3814da80db1466650cfce88cfa8d1fdef3399360050d33ac19ec48e9beb61a3765c836e92538428e6be96d19d455738b2bc147e5bf3b473b1771fd5532770ea8b1c8912da43565e1d151cc93efd2ad6e43f75f0e4e7b804a30edeeeed19ed1d30cd51f3c84fa6801138a3b68a5937ae1bee426f1b5215e0a80d40eac6ff88d087551b79ac5f73603e305eb546ef18687e06d489f41f4d22a77e403a4decd6b54f62140351348cd4b0f57690c8485d12a71a32752034826bd1b7c136e4641dcca1f5064829b310af548ff70bd59e7be5109d00ddd694652b7745599016de734c480172f803ea8a5c8a4febfe352887992918ad17c24278b42a1e2593e712147063d0ee5df4680d6f58c0687f5db095cc3e7a5dbb5cf24682a2dba83554bda6d39592e209030b8e947d156d45ca9c2062c59d61c0fb972eff0c6b42c1a866b009492ae4b4ebe3054eac26493f42f15ceda010e57c08e43f36877c2b2839c24bdca493bd380ee83b4f3c4b7c4d5c011fc6654fba147fcd3d8a698be94cc92b83389d18002a788c891797bf2d590cc0def1673f292a31baea367fc917b6720f2f4d74005806544d3f6fea4f46557a494668bb652d6cd741467d8537d06b31332aacfa131820c427c57e92698c115114dda1415bf16fe896fefe13ebf035cc486d2669cd56a46d5bfc9014c2845f4f7d03aa3296b58dc6c022b8119b7bafee124924671b4de79ff5cdb6ce071811f77faf53289f33332c6355c54494e05ff701a9942f6f12b626ab9bc46a28022399d4262001c1255c686b0c959b1ddbea62dc711d0ac690969cdb8bb360a806789a9bc3c8fbc4a9cdff01dba2a9fe2fbf2bde448e4ea9cb8e43200e9ea35c8eb6efbede9e06652310487a4be81cd17d0787112867310970667152ed3844d1289aa39ef7385c4b2ce840ff6f2ebab857f78846;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hd7afa47ff3e1c31ce9dc39d1505935693f02b87e26e3c63431e2fa9f53e45187f8a81f3c5b5de34c7687449ccfdbc40d00cb97cbb70b558ad561335d496bf82987f579620574402d52e871bb8b2563a33a3e940c98f619a10f5cb637cfbe4d0be1865a34911ff6006d161064231264685308f818c7967de5192fcaa5a059e7027c4fe0ff1d3a5bb2155162a43e4ac0d4f32ba7211b453ccfc3c264757067d9ff351ad94b1b80392b9e539b6046e042c87b2c390859492a01f0e9477ad529a63f15d42d97bcf71292499820faf6812e2701a2a820685f1ccce568a36fc23ceeadbc1295fc9ba8c1702b4f75411722a97928ae40c661d8c1460f9f11e708e99d3d390bca0c44da0314b9260179277482b1954247d001564273a602d6b7109f991eadbc4ac46e0139aebdb8bf896cfdb3f6e0ae3b26da9755670174ee934a37ae88131195ef91e8d1fd9311f76476928e3db06a63a5d1bec5070365c8c1c4c9f86beb6ffc7711b286db8c7887158feb2c6853a56326d667b6389a8a16e94a88cf1db25413526116cb776cb0549a73ffb69c97d41aa29516ede6ec18d31eeebcd032784f48996398a51edad417cb0e424e9b9db892befe71d7b09d0c1c17d8eecfa1b963854e3249e5f6f4b5ed80fc4a7052c97071cf5809b11a39be34ceb0d2fa869ad44f7ce69b7bbdf656589080c9d0458bf6c4fa876bb321c01f4c013b3f02b2fe49e64e7b70945fe29aaaeb75a7b8b17af6f3b70673e1f3679a3506c59e5a25274f75ee9f1295f308babc3392f512329806407e747b2eeb10184bbf73926cb1ca78e603c1710f0c75a268f829a63d9bb70d126ff4e467872b0a35a68dc3b3b40a119699f71f07c443e0c84db54bf110e2015aafe73e52c932cb05c90c550eb25cfa77461676f298dfd46902c1d879a5efd08ca00847926257f1c50d2aa60c93f7d0dae4b42d4d8b8d6cb8b190244c6c7a216a7457e923ad3cb1e6e215425cb55aac661dc01f5668a8d954051fbf9a30dcf1b4cd8ccc41e6288aefa3a8022a808fff103655fb9f08e6bb6d2d69d1a635761cf7cd7cc09be64bea7528b2a6e7e4529e77715092d45a26a170cd10a43cc74239c695686b3d3bb338e949c08b87ff42ab71bf1d8769328516741f46dbcf9733aae56f312ff74ea2a72a0a02e97bdb9d3747458630228e9bdf4749b082a7c92d39f49384f4c01a9be2b4e3df0985514ca92b5903906b3742cbe33f11e0b60682be9c4fc1977d6cefa5011a93ad14444a97a5a38111ab9559e8cc5dd8799c5d01d888d673eedaa0d250a8bcbc6096765a68d85cbf7c2bf5ee3e6a1243b0b8f6e0b370ea4f4ddf577c4fca9443556f3ffa5c1e2d6602eacce8beda9cdb40f6a8a6516ba53bedbbc4628f2ace75a61ba66b5e90079675a4b548910b85d03d63f67bb0e500977fd7ab881cb3592c4ab67a18ec3f2bd8ec769ebdf9157dc3a0a932826ca2c43cc40de4c135bba34619400a467c9a14744db99ad865dcc0a63266785f7b4e888b46a1a25edd2f4b3ac43b15b4b6a4f9a3a671bb1b0779176b9fff810f04fc330b95271e97b69f0744dce0bdb0a2aec17ff74780b5ac19e22b63ec9786550ad328aca2a95805ec36d2792b45b1e16220172ab2a3ccb8aa0ceb7a6b7d536e156552c62bb4775bacb1077b80893759255a116c627e114787bba42ca8e3a7d64eb23e22419cea5d56739f9c681ec6417053669eb2a58a327b66ad34de136637c112a9deca4b27b86aeb72549f27059130b1eb6238e3aa1b2f7a8bec72fd09b4f9858938eb5e107d99effdf4655e9a44f55b3e612ae7a5044cdb17fbc2bf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hc5cb703c3ba8cca698ac2d0440d16162c9f7f4c73126a6eced204c36761ceb4350e73c94a74c4d189cf564d753cfb6e159f40fdfadeeaedf45b4d9ffaa1edaa47f82106324b3fd4e4fd52d0cfd5cdb0fc7f41a86fd5dd5381f6e9f9e87e970b8c96762a00ee0d83f18854e81c76dac1e56b0640e7a29c73827e66961d6a9d00ae2ff26f6f24fd2a95746b1ba3365d1e54bb8071c8e24259ad433af66c535a80ab0cbfd96afc173c78849d6f575b2b1de582a5ead0fe566f32ec7878bfff14969cb5e289f35f07e4710fc0b3163bdab86947476cfa6e9906f2e3830819b3fceba6bcd958018ff40e1b7b21dcc984e97ca4b6b9be99e81eafd5c6fc347f11bcf9aef4c2c9766fb7b03adcf9236b8f6d40fa9fb7a4b1b0ba5c45f65fa2c5816f0bfe17e499ed0ff0f790be1feebf90a1c0cdb2f047d7fe85879f6d32d5f6fc320b630a673fe59aa48f01bbe012dbaea729cf7b80d278d2fdffdcf8063c121923288dd93ecdc13152ffbf4a216a7c917f9254e5e39e07b9a1f364b81b4f07085c977a3e19382cba35727183f93897c55dae559c378e4daf20da52f3d4166e3e292676157572febdfc7e54b34cb4e0f4c45096d8a9a2b06121309b7150d9be689a2c33017da193fba2702c12cad9704164e12fb874253837894523da15d54ee8f7dad799da9415314c3e82334eb67ef5c9537dc42a753b70202feedba50ba1205e9ffcf1eceaa5351a562726b785b6089b5a03c18cfe0b85f3cdc9df2c23695682fd0bef06862c60bfee1227690b7d407b295c0960e20b62457850bc94ffb4a10392603a85a1222c411bdaf2d2bba4b3b16fe5ddbbc52c4406d6c2836dec5f903fb13386b40cf08bc5103569f5a07f68df0756a5f3abaf8f7b4d64f3de6ed052665ea22efb62d6877967c319e99382664008fca995bcb07b56547f901c1219c2582afd192ce5b2e89fadaa379074832dd869c23326528b29d3357d77ac10d3c7cfa9ba4874dfb8b451f633c808359f37212ad5b09efd893b9e266055b0a80bee7de52c47bd0bb49d5c3cb0e96b9b7cc7123dde34402bf61d2947d90d8d16f19800f67beb55b237ce1e8d5abe734a34229af5fe32bd425c205232abaf816789fb9d6b8e51f95f0beaba7501e64a69cb399061c5611512f93a87fcafba79d9eb663457b520a0faf3322f247e56a77a8c8b302a9608cc48da685bb77b1469f1b601a28d9bebd06be30b87823983857567e96cff52fc27232fd50967a61bb31c8e2eecb597d8c73c4d988a416006273bf67b0e1d7ab39053fea8e73eff2c0baa59665b918eb413e80c8e7602f912e12c73d14739dc1ab7b8e94a65a05f3023685ceb6af847190b499b35929ee8a7bff60afa50eddda8b3e0a6e05208c72690d039d4b6b983d7a35a9a80cab236d84a55c8f1ef03aefbd738844db3e2640bcf8e8fee3506d74dc99293eb858dc0496acc6255e513b869ca0f8244094d481f900b88ad080e9ccfb1aff47c479d26d4c03a29877a4979e638a5effc738bfa7eee1e1a651c88523442edf19d61325687e95c8201798b7ffb3702c8cad4a0d5a82babd9899e97a3c2a80dc987cdd23fd0287e0abcf97253b8fa539292048091030f7df4f5ff2f87be0889a8f3c3989b030aada015b2001a9b10673a2349c4fec82ddc35f73974e3e71aa73a8a47712fc1003b4924191caf7db19be70e4c7d24a21c3f4aba0a71874701effd4bfae54094c3d0d0446ef409680a6f629b34ea4209ffb3035bcc9e13d9db1071926f38a72da26e22e70d0f81ed5ae415cb579e1988ddf6fa074edeca448e5ee549b507f892f06c3c6dec127;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h64d8e54c33f2e6303cf1b074ec74683606a2438791d0057610504bc1cfb1bcedbe0a6dbd21c144ac2bc1355f8ed5767d4ab01022dee0ed6f790a16c13f9acab1bf1a0757fa6a14f16e8adc18c76f4097258d073153ef8851ce14a312b9a5af3c479e3651c2931bc09265d2693bd465bb015fe62374902fdbb48fb39f51f90ee631f33e3b0ec6cec54fed4bbc13c332a8bd9f860aa065e72eb2c7dd30645fc06fa050ec64dd91debcdceabd3c31df0f6fd5b23d797e61636eb672dfc7e72cc00a295497c7370d078fa8eae84a43b564e214506908712c68cae32e7d05a971411de7b1e25cba7b1f754f55518dce55b4c2ad5ad9adb35fa9d16c2dbb664abfc332548534161775ddc7180de628289227afe6e6361a62975bf3ee820e338faa2a9621ba52c74fee1b8b8e2b1dbca625464382d9d9113169da4613503d30a6f3ba45bcb1e83b62e3fb31f6a96519fb3e171aa4aaa5ddc842ca6de954190cd74c914abfa3fa6276a9bd43121065fac2037dfc606252471eeca11a5a12acf45629828524ce839ab6f47c1722c1b6c67ad18016629862e0cc15043ee24448a41abfd4f180942889c09280e7df64ef96833b510203ae58249cb3f49ec2adcc707aff74ced073567717139ad7d920556b964898bc721ce7baf14a02b0bf79e2484b82135878db1c7db5eaf86f45a8dd3ac031413a9bfb8a15517d457e7d822bb52938756a0675112169f685765a9c9e927e1d5021b9fed15b7b1c53f825356dd925c2a5f067be3400141a88d1dde06e9e418366b625faea6f344ea2bbce48f400b65895dfcde6acc88c7bfe0043e75daa74b4892297f0b4a4946f24727edf3ac442bfa26513a8461e7e21a65bdc268361eb4999a598969fa9221d69997cea8acd730a9472669f6b8e60bd2ca8794a4f21ea41494373a598043ced3721c0c38205ab2c87dc11e59a69674538e3493f87b10ab4a8c7c5e64d033474cd0fe87f35976aa26d42021ad12bd6d27bcd36f96f0bafa004fac353bf0ee61d5abfe988187869715de788a5d757d18061d3e57e701b71c7ed65a467804341176ce8889a97d88939c71ceda411afbd31c5e53dad1e73021e9af31e690773c2da2df6880f201ac39c1101b5044ea93f03294d6902165922f18935cedb74e387a6525b6a25f8b60882757263d6422b5e318bc5375d6cd2db9f352312e334782def614af39ea319c17a65054cdc24d07143d2591ef0ede8362cf4a918f66b9ce9a7368ee432383371c724c69655247f564f8b50f5a1d8c4076525632993ed8ddba4907b87b71706271b6283907c64df9f07932202119a89b3d8c48be01220840487aedb059d1224f70cb16a9c711619aa61778001f99ff6f9516655aa72e0063b6d84aa78d9028cfc44a22887e73b2d922ae0697f9af67ef6e17cff0d5b70bbf3a0deeae87a4aa3ffbc7f67698b521ffbce961193cb0f05387427d02303f2adf5e81de5f570b5d3f8e6739a23c430c81bf6add63628e32e4e55d140aacf6f43a6ac1dbc0cefd2d4a10c6940436696439a46a16512aab2e006d407c0f01a5ae6a8f287ee31dcd5f56f3d0b98ea04e5dc74c480ce3e23a288ba4cb1c3990cfd7af35ca730d875036cf44434bbc1e68e9aa4440c6613a4458c81b0606758fbd67340a27fb9134ccf1d825b183cf05cf3c6efe92a064acdc50b4d4493976fda9b6388e6bda29b3729a85491e627182b82511df316bd7299e1fc2adee2060aec21351fb7f42fad6ad9ed89497b5477bf7f80944b1bab8ab45af89723a65ed4ac97c65ce6f53a1c4ed1cc37382d798597239c6ebf7d9b76aa5dcaa297baf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hf4a5ef970bc203907515a2b13d34a0e4b1d420e2b525758dd9abb6487d8cbe14a428fde55a2fccd563ff39ea214ac587a29e11bda27c58545b5418878b2cb790d990158cb4e282aa5b3a82363897d510cd3f7407a0740ccb98a29637fa470eb60d7cd5cf94f8603783275f86f55e6fd22cf11569d4c8b4f9075e7dbc74a98fa7e6fd5d252ee09b500d9f511f409805b2c3591634bf7a4888391ada178cd343ca57b06e86b1ce6643e16e01512e619534d0b085c59a861ec94ab73dd8a5aa691f834e01ecbb9f2d670e48fbe7699b670c5934c86d2323fbfdfe87806de8361d807fd98546fe5706f9dc0f03f58bfffc073eb2eab92abfa6a54c14a65b227bf8c4ba751dcd51373475658e6048d4381d20625f856791a8ea879a4f95a9d4188a20ad2ce4f48d384234f70e0788e6242deaa249bf7c642270d62c52acd255f2ce108bf1451046f574fc57c26b4086b76acde46fa1d7836a02a9e13e700515be6a9f6e028f5a4e6f58389f5555df36ef962148916f94c3da5bddef32702ee08aabbce2e1daa9e7f85bc105175eaa5c06e7d925744273ef83f4a6e4f38553e54f7bf8adb43ba9913f57b8f38315da9c7d538bc3b300b9bb283e8af3f68a663c4f66b4fb91567418817f23f5e94a7268cd92ed68e3766c6f229259f7098e6dfd097acd2fb52736568763b4a0a1c7587213ff7b29be91121c2b3d02eea6205c88acc47db1861d2fb960443ded95b9b09815d287af6b17640ca8517321e632dbd7195faa0cc31296d5d9f495c79858d92e4f17a8786d5f9688a935c642ae715572d827f48dd7d62d5a54548467831e97c5e55ace83daece6ae7c69521d1a3ad48a42827faab2ecf63beb7f560d0829f6e523aff9cfaf5b3b90ed5eebf242099d3da0b5c2735dda24f9e5e5901ce8dde5000b70cc20bb7c899897e861b9120a00de798058374560b9768ec93d7742a4f07e6792fa9892411b02b528d877f51a4da24da2d9124ed2813b0a544be9f340c7192d4e5801ae73a2fa748f0d3360067a50f15c77eeda1ee08603f42c075aa67bfad606a499bc72f9e5ed255071afe9de970f175d0e2db7ab4a9e63a0c8076c85782ad5f6b9cfbe30421b14dc6f9b2517e9172664d7349106970bc88572e914d656df496e659e0e77b9606fbb220e1ef1e168f8c60270a663682a8be02f2b28c2b04e68920f4119cb03a101aee10dae83a99fb09dc6732308ff76ff975d75277c77bdc8a3737656a68323e3c6222f73bd8f7c5d938014d46cc70bbea20908fc4b8600380aa32ecfe45653502403c7c1e4e2e2b5d40e8788fd9b4c10da3571a6ec40249105c0b4d0bf7c818a6027283c81eb05228e0bbd93a5ce8f122b1159457110e90619985a7c91dcf1061abb7f13b3b3fc70419a35fb9ed7c7063915d2eea2c122a35b497a43cc2723c0432ebc2ba567bf43ce8a99fdee20fe0ec8e1fbb03afa83b2723061eb4f34c6aaaa6834e2fa3ab3cf1a121099e13e9b51d55bad93bad9d3c2759ae59ef5a8ab1e893c7d0393a59510623e95920444430676a089a470284edfa27994062c422756f43c82c7e6852107e90464806959feb8f3e3448e0ccb71efb2be9f4d3a190bf44614e2b58bb83a567a68e03df5df3f8c075f1bbfe402f3a04d108f06920b91eba367bcb6a41f0e0b852aec39888153961a1bb382df90bac92f5c74a6ddcbe7d9c9711d3cf8d32ae4ea682726c2c577c43620b02426d05f7723db3004bd4adb332ac2d608b6b357af3fa2c2d45fc85258f5a36a7b5333b2a07f5d742159ba8a5bb3b6f2f6e560ea4ec2a981e12160717afb0e2599e430ff5b97;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h26e6263882df958c65589ee98a8fd62981b7ec02145b8ca802fe3fb8b198e6e896e756809088ee62a5ad309f74542813b7820525ba0a8a4ec92c4df8bb7724877b9b9b994a864805d94df69083fd2f832353f19c0533d96d548798c042f2271f3cb6ee40239c01d55ac7dd52c21cb35aeb6c4e451e8b8921b8f744597b5282576610ba3ffb751c7569d26a003a57c4a127d4e8f2244a857e5852a3270366d4bd0831b49fe29eb0b748a4f25066a0ac27f560cc920fdb069e41d0db0cd79217d294c74e5ddda07839f045893fde497fadb53dcfc896c6608d0d1f17361a30acb4e16b1e0db6b83af6f622dc1ea9f04cbf88fabdb9cf2a889565a2479525054589651a7919c28c640b70a329b000352a17891d6c872b0201a96f79f9ab5911d79c30031673ed0a5370ff3115e501083a454a0a972e26fdedd69c1dc4e6adb8ba2cd81ba09391b232a1251438852c9587664eaceece2ba7748c447a2d60a71561ff9ede4674f22158f2daed60c47b7349e984a6d51ae659c8ce9f5fbde318521b50f5b4594d67f152cec3405ba9bb5b83e891978e1ae075df9b97dde0f3ecd25fe5e7878d96ed33e806f1ac202d3c2c7ef36d3705e6ce196583815a7d049cc6614d1ccacb01f0b7650a1033d25e5cf11a5f1958d3a9e101d51ddfbe8527ed9e07ffcc70f38f627454003f20d29b983001d2a70234af9fdeeb9fead8fbaa283371d145c30dd74607dc4e529ddd9c5190c3890a82c4fddbe12e10d99180887d27d3a5e397c5371a5dfa83f4fe53e590892fa616a8d0574c7eba60ac751040118474dc19c7fb5521285954c1b33358dbd080c8235912c91e3fcc40435be6f4a04d5d286224f6d9fb027fdb5cd81fe5e433af7476bbe1c6c419e3665bc793e37e93f601155e295a9eae6e7c5c9299ad6d244acbd3155abf18fb28de311a67204de16af6e54838d2a022f4fdd93907325c035ced43ec965fba1c6ffaf320d59c019e4ca92af55e22e053f040ba9cbee4466e8a762b36d3e10c7b05b1981e484faa47fd7d1c2396c2d41efacf78be03ef6470b8ec9eeefa0460ad6c7fb6a254c3e6074cd0466175c422874e529077b433d85a6408a6023233c21e9322acef8074479c226980058b923b3ec1d732de6dc0c825c1f141f718c978c418c360bcbcef11c77d4c3af4ed61a6522529e347ee653ccb4b18da80dbfa30b7e785b893ca13527cb5e367ece3cd039c90b97bd7619056c83f96b4726f3efaa3767f69d48fc9b43edd58b1018984083373641f63089a062b8ee303ed7cd07e6c45c96fd6e06e5c8904fc3f2fc396992f41623c07b10a63bdc1416eec777ec304f0af366dd829409826de06cf46107bd66ee4af7fc9208a5b1485b70d58948cda51f42429a77867423465d68bb0ccc6edca72e15d0db473e305e7a26b98e3279766c1c09ca26c2e9af2c1521e38fea3f8884765d7867db6a113711340eee90efe8bf92712b0472fa3c709a82053aef568bbc3837879fe73e85785d572aee5ddd93c2bc3c739c33e50185e4145b60c6f34506f8f95f277c3887c652293ef7310bf00d20ffb04891849a651a096a37e9896cf1febc8ffe91ad0e58f8842e6f4197f2fcfc2e2c0b6129aeb5551791a3d8d44c72f04d9e60fa0e5fb043a32d1052327b0ae6120822e53647301e27f6ff302cdd1d94049d17ec65dfa99accea9fb0df6e167fa7a79c69ae2979d9a6156c22495d9b8af8f08f889b0f56ad9628e73edae582d2cf0b36e840c19d06ac21667669c23ec7c7695a4faf45cb2f04e574632b3633729d245a064b971016b54bfd8c79f630d3b7c742a0fe4cca6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hed2978e41c55e6cb83f8fd67f8fbd6da71672919117ab5800de807cd44a69ecaadb80bbb07bf02c485899aa11a4fe71db462323c42f2a52fb97ff72a82d13c31f35d7e79000ec44966c1007eb98491dbe68357debe0c5b2d0a7f189cd7f46416bd23b7a6c1daa30081b8952852d4911516526c94eae893d8efbcbfcf66e8beb81e2cfa5495192a70d6b0985416c52e64ec9408a51fa06d9f1ccc75da4a5d07d3b0b7846b55195a2112df408bc0b92ce5a2df8f63afd4d5c4efb772a31d4e3cde7729d669c4f1938fa7742504f85b0081a699bbe337ef59ac4b8126ddc254e7f48e82e738e3ae68832ab4f11ca6636b474a62ad7e03082671f8fb6f47f83b934102e9421a638a119ba30e639ecc29f216316489dec29da93906328064d7f5b1c7b6ef5179a593307b5877c3b510d567ba0c00183d462eacc301e19bb2916b92cfd0b32e6a63a05b5c47413ba72a7fbfca45ac8134107e45cf87c085e825f16ef2e09bd819e2868890f6a879cfad32233baf58e48e378bf052d1a907a1cb1e82cd7efe521b7d67f8d3619585453dd331210222ca7af3fff0833fb34764744bb882dcf07b91fc3e5179ebd9e0c89356658b8072dfc8048cd991de451d6edb32c7e1d081d4187a532afb1a25d8710d97488b3bf29ef6b3b837579c6911a6fd61f1929e81ace97da3b3d9cc4924d78e8e06f7bafb46c169b5e12358cc013eb7a5abd823269ae1c84162ee70d89fed2b7793d577f88516e377c39c5f4054a080609e3073a2a5d735bcf381ec008b8871584e8318f148284bf7fe997aa015d06f68d7a9b880706ef2bc67859e152e0bc9596eb67185d85513cea3d859a912e7578b46ffe6f4841745c4dabd959cf4fcfce338694846b1285c10092ab9c60b44475c47938a9047f278b00b361cc47b26faf066f66a0b4f7f88f7c5d2937e4f23124b570ff19a662daf2a815265f2a013336ef8a188f3243057a71e3ac1fef01a1cab9ca94e7235f44b556963488b3a73eb6970b51b557884c6e9b5f0b1345118fea33f4a6d5b80546b4cabf9474ecb206de54795c65f17f7b0a16ee30c03c5d19ef22ba63dcccbb7509cec2968117af75f74bf4c7a0c9d9e136e2eb61d70cda413d3fe8ac7849901a6d2bda638b72c1975730c94529b5a07e00db76bec65189dc7fae58044b3efb27d1bd4b84ec23bd5f12e20c0c5f85647fc99f04e0f0604e7e6c59916eee08cf5fbce18f1748501bd05f8afff710177fdc1e178d72effdffa00a4b09b5f113e277b5c8ffd22d1bce1deab18fb180043d95f0fbb3eca6b7aba5b598173a4baa9223f137297d2f15651283c0ade751e346f8b55388a1b49877ff77c6a52a8054272c3f1fa2234cd3c530ce808883135d8c0c4f6bd50b0bcb5d1b75ac40b501bfd7fc3e4193c044c1444f4a285fc97d071a4873e9df341f2e90d7244c4a54da49ce33bc6d720a8ca6427e821d04d5b0a7231d6fd0893f313ea2092818b27d9ff57a4341267ae232f6f9ac094cec3af9331af212380d120d5e7e2544f706499ed7dbdff12a74b5b897b096363b45b8f6aa4ee9e5d0ff1004e4ca7886eec95901149c22d79582183ad229fed9384996eae25659217dcccba933a01c1f436b1dc2ecc42c1fe86d8a181f87c4b41ce9e06d853ff3ad8ca83d8b0ee94715ff07f86ffd1ff7d73e4a40af655ba8d94a6e5769789880aa157c4d7120a928f75bc0c00bfd0e9477448414d2b2d919514cca13818eeb5be75df9e4a1c0ceed4df3f0764fa6bce71707ea8262a0fc9a55d3778a4f263190cc36232bba1f5ad598e951349d4aec450fb84a3bb49796813db4afb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hf3f9e509670c8c35f716e3fdc2d939fb9ac8fd124838beac04bdb724e528e9d4d3a96c0727db74f786030914979518ae823f0372d09926082264534270d5076db8511ce65142cddffedc267b4573724564293e1af288d3dc559d51430b1a232f8273e4a7531d14f5959bbcfc651104b31060cfa904cc44f2f46c6b7cbf3acd1ebc705cc7b081278ab594421f5714fa7333c98a24193f6b90612db00b19a08680dbb7e174e205c145388afce132d8b3edff6ed60e2f196f50a3277f93fc05517fcd4d693c3ae1af3efc2412bfc03871dc32bb346b7354e08caf8c3f5a79fa0c0601640096ee42d6e86175d9190d6d51e413d3b5ffec98d15f9427576adbfed4796a9cfa02c7e594baf2dcecf43252584d4713a3bc084cd571f005532c4339decd15a7f9aeaa1aa99b238c0f9fc57bfa90707908eb62b6a7daae30ca157c67bed19dfc6c2c62f25c9de86a7606aae03cb38d65795b77404f9c1821cfb3aa62ef7af128f8a57260d837c415debeea2ce25b2d1aa1f531073aa25379d3c8cdac02ab872598f2888a38bdc60c640155aadaaabf2d2ac216a3365579830b94ddc18e4c56e93e35c0c361a6a214b0ef556306bd173da5927d46b698564f37d1051f74c9ef3258506cbccb6828de80b0ee15f41ce4620f5e097228b9afafe311dc313536e275945dea05427a629535cb0fc0ec29dfd020914c0880a74887fffa2c5f4f918029f76dd695dc9b8fccd7439eaa082f3b48c8659465a536c31c1c6e16860dd17ae9af989579847f0dc9cd6fb563ebd2b2350eaf353a175a4e22552f3e2c67c09113034a2fc9525c2515e175206fb1593b98e0d5206a9d525b754148be47fe6948caa37dff24f6fd8fb38c9111ea4dd7029b7b7727212c5dc5a0e57bd358d18b1398dd6cfb3eb1ed2a112efedc1a203c92d3f142254129c2e6c95474c4340465c24183016d8e18f294acc4806710b77ed2cfb960cc8f429057958a2048e4a4efa25a3ed56ce638cc0e3b81d68be7365265ff60ec2b9d86768e973f45b112212cc3dbfa2c397811756f8734e9f09ff6cb9b9e6360424da03a811ff5ddb7bc9b40880a9a5b79202d226cb72704cdfaab766585c5c6ac0ea3d2cec8ee97740c24e6c48abe969d36f407f6fab21f5030095d9f72a4548693c9aef3dce2d899d213b6c06f1c7b7b73a7f6ed239c2fd6b38bf7a03f9cb6ca88b5b0f164af977cb328f38b509da3946fd64823857909afcbd2a84088ea25793aaca0d552330352576568eeb28a55573ece73eed0fad81c1c085230a9d4f9ef8cb0506d29f4e17e522af7ed1de537cdd422566a43acb1b0595b25ec9e8cf7f7759f1840d233831ec5f3f9cedc742da43aef1e0529ff81aa2864c949197ca4e70c6716f639337b11cfdc4e502c5682f3a58f7cbe861c209c978e52319174edfdad02b144adebabd1383b74bba9031dc301f6dbc98a50aab02d4400f4b17c934d6c85763201dd0d1fe7431df9c8f76f69cf26f7ec0ab0d0d24081d3f854e25dc19bc24d1ed2ef6adef6553e8dc3498f2dbe7b023504e4f7f3c78db55e41b1bbb51fbadf5bf8b3f8cfcee76fadf4631b7f9b5fb96be6f1ff0dc010da39dc97648fb7eaaa0d759453577dfd5d26e3c2651c497f03c3724b084a251afd6dfba733cc97fa2c6eafc7c58e3bed8d532610b2448bcb3645d01d66f48a7b9a99e58e8b075d6ec9f22d2424a6850e1b03cea3e38f6235353b2b0831b9865d2d0f68a38b933f90c526c26bbd72150904d3a1f010f7db578841045bafb092b90bc6a466eb5013394018fc1f1ab3a9a8a717769a838383e7a79d29e5d26418d6c1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3da02747191e6abb8d8be78ac106f65cb22bc3c7e48dcf51e2c517a72c235273a578d2d3789b71b2edcec56c6a6d58f3c0bb9f354ad3fcef53b6a8b587bb4983d2be70244942e7fa6fca628a76ae1cab97d6f4bd79da4311d30e6fb0deb9007cd597961c75d142f0edde5cf72282045d1677636cdf2a6746e424ee17e25d07e12a11350ad57301ad0718e27193e69349a49de3eec72c20e7a70393fe3fcf128ad028ac39fbbf5994bcf86eeff1b62fc4e7b62be27a415d14d936a9431a9d59a98228b356d67bf29188792305dd11b542b3d8c72e5faaa5c147f54c4174d639b5d2f6218a371f2541533af6ddd31c2853357f7abae1f8d837c91da07f6414041d566739916934aa24e52948287fe4015c946a4c4462f3c3d311088efab56d16c9196ff85ad757977ea2b3c8f4f624a7829973d647b6b3bee8e691e4d0509cacc8293303b250d4f7a64605d4df102f0e4582b7459e4c9b4a733ec8e71cc9b61f706f4cb8564db51192375381b614adce01c76686bd0aa9e431437b57ca35f9c35d8028b097e1a310253931a9426e7d7d40ffa597def9d1f4ac032d232ecbd4e596dd581d71c594267ecd76a7381474cecaf9f702506a22a4fc1c22d20c2024786bba86de5f28260e72b908dd2ad966d64b96f89176d9134141b2ff8645981b590ad7fa4e73dadeb610739660a40cf4a4eae764a10bf406f7fd65fabb399e97d06fdb5acbaaeb332fcf228b8927da5b2ac5cccc790744494e0ac1db737f103ebfcbd1f8d64a4998becf2758624f47a22c04dab6d92a12db866d0f4a01c38387d2b033d6e382f41a92a456d1d8e9a4920cdc5bbee0063de436378c69f95600828e11836d662efe1b394fd16f49bce81827a0235e2c9098048fe0bbe944714257d2a8a1546871b66590da42778ffb933e64ddb0d0de6c056d2a1243c4f57cee55f82089a917678b3be2b2d7782aaffafedabee2c7f785e9ecd26dd5ca9854c3d93abec7bb39b3cccc98a968d0dab364a7630822ef053a81cc146ccb2bf946ad757756de92b142949b5af808650b93aae99fc2d8ddc33198fa1f70c0b602a011575f85fbff9e77edb09e0ff546f9fbd21061df80d6011d93b22362dcd84eef1b61749981d7492315a8209906b87e70de91f7e1c9a077b4286faa9b8a1dc3558cf558324a06d94a0794b05cc2444e1d0b5d31cbd788a9e920192fa5e3356d10848566a414f2c8f4cb657f6331c429cd506f29f876165b2b212763f39bf5b9f4531024743901c1cf0b91f8ef5be0613bff5f34e288332384e05797c5a7f0ad66cca13600bd2f9616a9a978e0641fc8f219202cdf86567d103b5dea98a3a081cc837f13b7c1baf42f4728779a30922cf2710942fb64ff808d2589479878fd2c58e2db6c71a27e8030c20cf6ecab8a72af6412f4a65a01f548e8497fe16629a44c66339d4fc988d4bb45c4e6c0a6acc6449357658aa5ca330f4c5668244e9ec468a465e8595b9ab6808f9377bfcc75e2da7b2d066f57f30baab99cb61aebe28ca8f9cc017b928bcf8910034ec2848da9a5b384404badac4776fc5476ba1dc44baa5d127005e3b92288b48d76ed4df81e66d13f869106603bedb2bc5e9d46c7b5411b4d9c63f0fb62034ad09ad7b5a5c69a45900b0aa1178945487ece40f2ab8d83c36bd466ba669c57c08544bd7e4d05ab7819a2853a18530073718372e55ee2e2ec5a7a4ef0d6d42a507e484b26fde93beb28ac11173ee0401de30253666bd73a55205ac76f8f265d56948cddbfafbab34f2ef93228f15c7bc165ecf86cfaa906d5ec207efaa780d33979a22f15d40e6ad1e1429d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h197f891b1696309ae0294ce56c9f4a2371a20f7e497bd3dfb7b0cf2e2c32e7d531de8884b05307b937f22933ce4456a6fe90e66aab2e017a8af58d993bca6822e91826a6697fc431bb878079dbf654af926b9c8e3b4add87f14791ec58f0d7505c28f69425c4b6dfb29c0fc6f139172ee7090eb3d5ff7b266a646ca31d1527309b1e68c95409120761e1f51c6d6148ed5a1e35a22d541e906999d48bea5bed6df562a6e329b81bb0f0b85d247bdf3e7a1d8de480d504b7319852088697a77e98d815bb8f7cb391577182406836b21f190395f186af40769cb51deed99a205aa7a4b7f75e9f180a6249245ff56b3c12db05e54803884f04c41fd2c95b65080b2b04b329a52ba1dac3a923160fbac46ec905bd8e0001fe789645ba1cdb54c9d0e113ac1c3b9fa78df9eb2cb955d57a191ee78a4bfed5d3f49d10e752b326f518b30c659b91a9dcf2be79f0f26d9b6974195892ebb7b64a5a8c5496c701539f1aa9e055a3d6f303371244861f7ad9cf62fc13f5569bb1d9b46149f626aa55103577906560eabe928d1e3bf5a0d3f0523b4efda6e839f08abf1e3d398b26afb99c801c28cd278a69d5f89e646de9409f85911d3a86787b8aa9c252ce4725c7685312353ac1cd2613104a5d5f2bffecc7427015f97af9676c62db2e58507d6a4476b88d6fa98558ad1aab306a76a2a806d77b33298f22fcd88872ba5369902aeb6b32c0332ed3e077ad64e5abd21b6df6c8e8d70284e0ece1388ca559faae02ebad1c7458a5d2feabedcf88e687b4f04c8e47a06bab79db539ee68f52948d0e21911a4ca4875f34a7b0040b25b84b0f744e42839d2d096c2b64e0366f169a75b1daa29534332471fc1711b13d79f0ea9f0c9fdd263a996422f562495352f3076483e97022dad15931244eeac0edfdd64094b07704fe003161cf3f752c7bebcb77f9db904d18e2bddb40bb7d1d51e1d2b27cb89cdc6ec7fe134eb5cef59c9cf753a0af8309b06123cbbd62f6b0f398b6efe0aea51d870f381a0f3d930936342f2b3b0de8cf9ae9c6e57ec6c0d6bef46c7f288dddb3c0fd9d71ac6edbef6d8b1ec38e716876ab24af9f5b511ca2910936ce77e7263a3028ec8699a65b469afa8fcfe861cdac3ecefe46f2fa51b9979d97a2976cdf855404684e57b027579ab9abb1d764aa44383c74807579fda68501e9be0c0e2331e187ece4e1adb592637e6be162d49af3bdea9d3fbce63a3bb7c9e84492ae6993b88868e29caf672e1f22f093f21d8feb7c41597a2e7c5f53f4d7a6b71dde044443aa5c8d592e01c42676ec0c1c8a30fc6560aa50b01f9d254133fffcd9663367869bfe61951494849aebbe30356227e3de984cd4230a6f7a00d8c5c74cd8285df54995454ed5a128512e77f8d2228086d09a621e0dae6d99be7eddfafc47e2599565178a79d925ba1fd9682126072425486d66d5fc8836abab39782cb7bc9f24f2c789361f54c7c65ec2cbf4c3126ac380f36e28b91ae6f05d0ae87ab7013b52806f23e6e485d070361404e4f08f8277c251c0855e33086bb486b1a423d92dfad47c923542a5025a6a96b4c9c7daa207260d02640d70be3829d0b01c2e7b997725f6c84dbd948047d642d36f2ed0a19632a9fdb5c61a82c312b4052c68544c50c6e9f5c52683d7a6154870398955dd29ee428dc96f535b542e881eaddfb9ae485acca9a692b951ecd19cab5eda8ce4b31c88be0eb98a3180c9cb92df18a3c396febb0a23dcd981cf15ebddee7f2b39acf9f5af2fd2a5440628b4d381ef4793a9ea24291d9bd96f7ed9549dc0c02bb5155563b2271e4c7bf25fe0b3682917;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2c3105fe15cf55e8ff10aba81e541494a201e4572567d7cfb19b87c286b3897eba60bfe95d1d3bfe35b968c97cbb9c0b8bd5aadd7cfd6b76358cc17ddc694850783fc823a9525e9d122cf1c8489d68b810fbb3e262f13eb40756fd81e22b8c240a04e6894f3f6bc3183be1bcaf1f23995b67da1e873d6340e61c12f150d9336b3c2b34bae603d84797c9048e665c973eb23a897f7e56017640c01b5cfc4b2aafcf138167d1f3a3fc6bc53816f86d44f4f1eb2e31e03c97d61333eebf9613c04de4499caad68718a6227f3652ce6186d3b9f1683a5cef2e02d31352bd2617669693f6ffeef8cf00a2aae30f15a8f33544ba9fb1cb316408a5a270a3f042ea2517f2e30d1c9e490f090dfa1c5e84a3fa9f6d74267a7e961601fe89c2fb05e925bbdb2961c0114b19313f3ad6a7ea7af3c568ef7073c0431fa57644c42aac1ce7ac5cf776c56c89b637a65e67f63a22d85f097e56bb27540823cff34cf644637a5b1c5deb08d7106e73010ffb404847c8c157fd7d8566a36edcdebeb79a3890eaec06626ffcaadd348ffbb195aa168e4f56e8d4ccc9abaec8ffbbbac3b3cd9688e7cedd9f92d869d5010fc81b1361ca6d2092fd1f8a500ce3cbfb904167c437bc67b5cd978cfe3bd84687fc29ab303d23a7c1b82952f9c6163f37215b1c8335456dab6523ff0a47663763ed0e191607b15608261fc5562badef279db10d5b598f7a5cf191828247623a1811e87f9654697276e989abe6f071b97ddbedeecf12281f1ea594c082e239727ded220636d19598c13d1c21909fdc380896700a0bc557b676bc74c78ba5aee0552dc59fec2dc34ace720a60f94b770d2238da0586b5eb47f6c326dc02950590d9d53488c838471272d1efa44ba3e97412f65776e5d307b5131f04361cc1695fc5346198a3e0c720115f262a01cbbae5dda99d4dbe88f844a92ee062f99441ce6c8fa07b14a432fbfccdb7e680816cc5bc834391c88d8c6941e1de53836409ed58f5852e16920a60f6dcb05d73d22ee5062bfcb94fd86d3357ef239ea03dece371753a661da64e31b68bc2dc5712e50a3276c7232e970fc39bd36415cfb9560f9c92b37b2e7aa1c11261776459f9012d85a8989c1da10b3acb89dd59f04a8eed38f86e6aeaaabc732885408248a45788d4545804d8d9da37bdc9c7cf6935177b7468f515cd2508710e3a8cc7833875b299b12a9e19f5a1e3fdb18350e8a52c6eccca0c44b924853645c487d61e4e54cced8eb20efe1d16fa27e6b5059de00f4b1186e19eaa1bd853327061c771f630779e115ced0d3921e3362c9ff0c7e4b4c6a7933f3b01f8bb1a4af5a50eb112ee05a404714ca5865f859a9c62c6bd802878c69a3e92de0c657c5b56134691bb07ca10d106ad8b0321d0cb7513b87b188248689126a82aff5e70433dee2ce778c21fb4236dc1ddc65c96dc08ac02e82433beea66a052912b62eb9d0d3b4a9f858a1564f70e1a5274174874caeeea07e7ab52278d8962031e27c1789bfb5268b8a46176284c1fc1dd09b025b04e60ff284b21f590d1fffce8e6a24869203dd6246425f2d3e4a607db828a74a396d6ef446a801cbf1f84d93440fee283e28578f145b47bca28c3850382eb3ff112db596c14d44b28024e85ecee0aab12d84475b37236805cf43e44ae85fd46eb6cfc3eb282ff99000d8df1d77fcda3427044667244799e4e026755f5d6b00db0294368119bfaec86fe32024d4ddcae96847b749927c120cfcaa4375e67397a18321ce53dddf8aa2fb78b3e2eeb48880b1a5f5d68e43a5832f8cb382c5e885fbd249c489c86ee08ed6691ee5d50d5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h6c195299fa08d619fe5d324a13b44a45c299ffeb557aec381204667216bd6034924e3b0641512f6b13a32ed61b558d788a406f2824af3fb99c37b643769c3e42741952ed8a60c0305259e8da8104b4db73d1db7e737575151d97e68b2662838c6d80679dbbdeddba1e47f711ead52cb77c6bbe4418de700dbbb6cb6d87253eb737d582757759942ed33ec3cf619613ad7618ae26b49a70e0c9f795a5bb46cd6869e48ffa6fe90bef1b9b7a5f082a4a3b0c9c135a32c892c40125fe18ea1fea01bafb6ffda0d99726f4ac489cb9debf0ee0966313d3e167af6ae17a1fc4a38a3b90d05f4f6fc340c1eb3fdc2d2a8eda415c73fb5e48b80cee613fa3ea4eee08bfdca1f48a4f4d0cf2f309eb32b44ba9f595a0d18092e08675d3dfa8a71d28549b065e2e36813bc05a1057ad7a5d319072490c831e179228ac1f92daff030da57bd03ee0d91e24e0348a2718c9d08474af25433fa2de61f6b7d73c89fb10ef38b6d8804fe3594dc6c95b5014dd9e71a13987c385c494cf278de18fe07b25b460c2ae9c5e6d031220f140967db7c62f597840f28011a108ca45db36fc3a8937c0d5de7df1c6d828151d61c4954ee2a22d1c7c4d069031f20858e48edde383f5bbf4bfeb48a2a39337bca4a4bcebb33ac5265453113e250040321672cc8ed8cd75c17652dd42f9aa5026d64f380b20e61bc5e031772a2986dca8a2156626805a5d31f9fc1997c76dccb2c8968ba2383ca39e0e1a5482a1709fcdd937e1ae162e167393ad3c1726c950447b87ad26722338c0c23fef0f27ef1009df9d3c0593bb7534cc97a4d63b459e2d20f666982378007fd813ae89b46d5c452093b91606fc543b63c1a162a1307094b923259fbea65edea46cba4a69808ce0076e6774324518fd70357bbb694aba0320da53889be9b64a52990ebd96ce38cb3ce0ab7c925394418ece0673b3fc27d2b6f24236787c54c788d24c8b31ba38f4dc223e4f78f6ceff66bb07603d26fb6bb5f10baa54945e0d27eb1bac46c9207ab4b5eed573716fc21187c097c8ac25b2745c6959a09d04bc27df6b759606e5b7386aabb9fc3969da286f125d71b936bfc32afaad66d585b517e74819286bce3cec8d399c257166f944a8fde66e49ca89b11de7564fad3061b4b18b05353ac74f17ba68583b37eb68fedef9206b59f60e36b93ef20e880087f3563bb758d46ebd5c7bf36bbb8bb92408f7ddf0c65ca58f898ebfe5c0c0604a435046a4a6792b5095d61093facdf3850817ea6c5b9734d59547f7ef6a2dc2fb324f29d480ccf1ed59362f57ee0b9b353d0e93ca9e8f7987217705f0697ed6ca55a32879733f149e0cedd96c35657123547cfa33b9458dd24f57cfab3f3b1bec12a784a014c3501233176ca6248c7d432a1b4bcf2d8adabcde24e7b9f59edb4f6aa20cc4cb71d68118c18690e3623b902fb3de61f860321adb3965bb5f6fed92525e09c73d264f2ccc22b330409a7f1054159e2d4398e865ae4dd54dbc4a3640d0b0baab92da5f67e79c47a6b7d0cb3ef09d511dd1953ad4388507ad49f34fd535f529f3c972ab148010717b25b0b1449120cba6c9e04a2629a483cb4d3e2e11ea3a836b9e3fb95e8a4501bdaaf1f1751b7bb7ac1b258cbf34e7bba61fbd4aa6c905061fc56784dd283c8ff580967ceb95ecf7b39e06ff9e36b6f74d61f86ae7387b088a610a60d5c46110633fab654a875ef7d29666fc984d30e3cc2d8da0131e70b1271b7c2b48d831a57b93fc6ddfdfd4bd041c326f7b3b43ca60e7d513d44077ae109853c020ba15e96dfdec8ed30385adbc8a6613f44a19c55e7dd14e8a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h6db1cd219ab6e699824adb2a6726f5235abb359a082a22296a93c49f1972c420303d21ee5bb2e788c2081690d0e5bc67f2b27388caf02270e1f98a65f5ee153c780846f1b2054597f1cd5de65bf58d5ca4cc810ad59fe8eefb7df543ce720206bb548a9fd597065d7e8b7250f892faa6cae54ad990fe07233175b4058b48fb9078540172920becb1854acfa4464a3bc369500a2930f3d742bf29ffe235fb3391e75b77a6be10b1440c4f393d010fb855bcec778cd430cef89c8bca63ee564e3dbd6a74c71f3225f7eeb4e95dc9c83ccedb015dbfaa558eddc407b6dd3cff505938f261ebe5604c36c71da617cc590b5c8e42ecc105c117de09b7f9fe7b7689c04b99226a11704f18c70c7f1442e8dec8a8f2ea6010be358d971d835f25089148360f68fb918e043eab3d0c25db6cf3ab88c7afa0f2824baf13e8a3b3563ffd0544a96018ea8d0f228067a1a9c73add35cef7146f2cf1f91b74056e233dcd0a54c2efa9c7f6d5694bbfb10542c0d75926c4ad2f611631419ee7d2c3c4ff7cdf0ed0c194f1688a701952520a62e2c43b2f73b53208328b56fe65dd131ee29764e7db828e89dec17236fb8d9aaa9b86d52208d09bc03a6f4f0fdf8404f2bbb90b0ee6e0d58dfbbfe20f4d7d4c9c33b6e8c3a03161123d61068375ebd6d19fd5e6801c53004074172f024a5ff947ff74e2a21e2f741708f14554470c5dee7ab92eea33d49d7faa573605efcc8932329baf45d66657d4ed5824ae9ab62e6d7b64668cff6e46ae13634d299a8af85db448fdb87d91357017db5cedadb0c4c54c8c19822c0df0f58335bb682ed6456f872053cbee66d5fd8758035ebe50bb09284926a38247a544443f4ee965f8129a00e6b5d7427b8aa0f2e827a58d22f0b925f0f9f4add340daab8fecab3d59409052b86f3262156659053db31fdaeb074409a2fa5bc4777482bb3db880ecf5cfffb5e0749114b74a06463d9e926b3847f3288393dff567e464d341f8ed5c261e2addce0478d4e735eacad43b4c3a4247ecb5aa84841e6a236099fbb69fe9c3cc934f665f7badec72cc75dea6f81aaa743b8afd8c7feaa53a3a861bb4fae5068bb1c62f5cea6fb1d422ad511f42454b3b5f176936f72ad2aa38645f94de85c6fdc4802d19805871c2b9fba486140eb76ccc9959c94ec1f3e9f439060711493c5b359ffd9ad5462c8a7653d442c05b89b72df62d0b8f00a55595caa6ac4d6ed840d31464072cd5abd24219cdbf29d964ccd9179b17d134bdbce533d950aac2fd50b772608fa54fe13b891aca5b40a6c329980dd7cc3c1e5dbae46c958f5c8a7c396aa23a886695cd88e638e3aafe7534c618ce481d8423147499461dfaa4aa300b30b525bbe2a1622957b0d266ae25f6b98f2d59edd28179cd0359807e127bd04e984fc3fd1f1012e24352b84ae677f46286ac612abc625768bfcd4fe2cbef88c44240bf10cab355583495cd2b6ce14626f8226f57b3425e30fa5f5aba65a733db371d25c35d0f3e2bc9c629e481afa971ea4162b78256d131688925a2ce05b6da2b6f850631182e4f1a7eefebd5d4f249849f9a24d67613f3dce0d0fb0e0d97aba0391dc1174eb6fbb1de6c46a52bfac36c5d9a7914c3b73eb43b93ba63d4e7ac9cf85019298f133436a613758479a90189e69352389ca24b7038580c39c02511e64988a1ff89f1cbd845a4952706547a39cb5f4805a216d1ac03a80dc6f809b1622ddf5fd0a81f45b36daa499310b034d7b83e92d5a8bed6d75af2b622b5be6bb79260829addc67f394ffabf8f151f9d8647ef9f3c674e1a5178cb91500b0a40095939db5d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hfbfe32fd480f1a82853570339d69ebcd29e808772bab20273205bcac63558e7434a81102392557064fc5b78a3dc119d3179a846bb4a38dd6ca53a9ccece8fd6d0428b63078843934f606e5611702d03c98a14d63166f940d86c293c37a095ae0b1308a88ac6bb3650ba36955e475d681b8d9ce1d59ed5d4e787a719a5d9ab803cda88dee23e37829d3133733bb21c2e93363f8b1a1839e72a08b5f0558bd3cd7a6ff8bc51e450b518c00cc59fdb5ca9ce9068426130571072a4884bbaa7ecae7c75c602e87d9b3714807d2b21ebee728fceb94958f8cb41761c6d60239238e8191152aa764ec82d8ad255f54d8b842e0b62c6e2ec79e23c1400e0ee94c2b696c8c8accd1ab3d686044067ad021b4f3368c111d3c593d371462bb0ce6150fe2588017aeb0d40592eabc5b6fc9db10727a8748dca66ec78c571fc437856d5e4547dbcd7aae81107ec49855161f6ea60f2c5c5b1fefcc77f7309da4e6d67a8180c1fc63208e8767da6d3b1d0a3f1e6daafbe14bef4c500535365014211511e2062635fae3d83e276a43b40a260f49dedec9ed92a1f3209d637dba2c7500bcbabc868be09a2ca8e851e6cc2a5705643652147ad702ebba9d20cc2fcf67d9af2180e86fdc4c831278149cbb862294d65cf77e714ae2c930b2005a4edbdf269aaa9e9fce40bb9a608ed8c4cdd620234eba12728831fa02e16154e380cc19c4f4667b522987159e0a174a6b065d12493b177b951983872428dc6a46880964adc18b1891bd1f938aae03fb379c77dafd43bab75020863cb57fc707162c5393c74ed1a2b1c2c09f5ef2bee9f2539b512107179f1d2e33711fd7ceece22500dc5f93517b0136903c2feb0ec5e42aca5a23f5cf22dddd28022cf0709366e4d73c96dabab3e2c43c0082a1c2574841285eabd4c71d56177e67751c72e84506504bd70f24627a7082353152ebfd3911202c37e140f1a7e803ab1c49953691652a4570b207466db4444787bd2f588bc96a730eac3c65e3be26d1c8c80a0a16658fa84b8f95526c263d0aea68092103b9fe86cff3a422bb24c6bf64cca85dd4d55a69f40f748a406a87207002dadcd908f6c2b3c109f1eb66619dd394097047f8a0442edff06c7dd7673a3cbd9da43deb56337501d69cd3a22070eb8e3e3418b3304d0536eb9c6d2842c9066b13d44f83ae36d0600998eb8136e2c1dd06d1c784e157f841c4cb8fc44e9a7677a5f73b0e1c56ed35a2853ed2c2af1a43a60ccc9e9d6cb66dac1bc7a1e9672827972aa075aad06e086307ee51799d982165741c7c7759a53bf6ece144692783db6eee542f5cb628d64fc5d8a3969bf95bb117bd3f0bad1cb214be4c6b1c48de49c3377fffd5e5c61e7940a8d3a0c47e1c2ef16025420495eeabb907da4fa13fdfae20f0ebdbb79c018158f2fe70697f285771c23313ec776037953c9ed9a816cc231279da42456ffbf26de0c444821d6880b0a0e982cdb8ae0bfe59ccc392ab5796b36da8e0bb1b88b6b93175c5ec7c5abb095d76580d9770c4861468414f15a3b023555db95a03369e279331ffcb7f46c2ad4ea9e35d133ca4711a57274844a3d8710dd84b12eb5f7098f92d78589101f34840625ecf63a8cfa14fa86ba78e8c22c9c3e79676fdbe0c704f2399aa5dd810db62d9877602880b635a00d1b5f8d6442d1bdb06f0414d009d0fade20a7373d00effb71201f47f920a04280e1dd48788ee8130999a4924505224a31915e12cf1cd05812056e6b12d92cc6a7ab412afca66e82c9953e6bbf293bd95f5b289721b36b0dc0ff66c44e8b286416bd68f3e16412cb0b98e1778c2558e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h54a7d1f2d74261b5fa334bc2968bdbe715aa0503f1d8acd859d91bce48348e447d2302d159c65b371eb2b9cf0e81a9b624167aac0b557173555aef9cc36c25044ad4b294e4f78bc9825954eeab15ef275334f4157aef52d4f22a584d3847424148f64345559ae42e80456ff4b1d5746feade9b3c008aacb97e477c66c7316689283a8e240eeb64564b33a2f4a346e80ec813c61ec6135ed8be51f045e143016f7643bc6776ab8f82e5b4fe34db63985d15c2689f1ea3d3f8f506b4d59fb20788c1160ce7fb63f648dc20a4482879ba9a4a2d4d1edd6918946d9e5cdced22281b6ddf43b35af0017bdcffd864ae305f89238cb95a9b426a7480faf131d146274a28ee78daf231c73f2ef7efaa7f470c6bda28ed12f3ff1d7e5eaad414b4d56dc187789ed9754d6e673fccb98c48b974b93e02818e2b84b3b7ce07017749bb6b9c5b22bf3cf8d4970e7710122d5d4811be55b81a588245b6e543dbbecf342c32869a17de7cf8e65f5df0d26a44b6bff8d820c2a822a51185f1eda436b48305fb5bd4f3853dfd9c8965b6cc07fd37835cf0d6bd3d5ec33ec71634128981762580492875b2128eb4075b55ffa1fdd39074f913ee8931a4c7427db858179a078b48e7e94f2743b76b74c17aaba88dd47e1943ef2dde76a77b2bb4edc0e698fda646175570c7a34523e48aeb452e58b13ebc3b37ecbeaa62c977ae094034f09df5d80308427c525255f3f906d19130203f317c27096b2abd46d0620a79dad7a1e8f31d036fd276c622eda8aae9c1bfe668fc4e46f527dff24249a9e5a73d36e3aeb47a8cf24ba713f8cfa2df270bc1d3f8a05fc13928ecd6e359e805a9c57a9d0ded58c35e8f32866ff2400efbfe6e68711f8c06ec565cb1abab171a082faf00544ee1d4da6ecb3ccf45e229750f91d29e78dc85095c359f6d867358dbd04b0478f791a2f0c89c7a52be6c54d37f5bbbfe69c408681aa10bbe8ff7d65c7a68ea1e0c3cf9acd060d03b915c75313d7b6907700b3674079dcc717a66b0b31b427af02fc1395e55c5aa9bdef98068f3a09ae7d6bade40da4e90323f94ad17c562ebc4febea22e9dcb536e80a6fdaa6d7ff46b542e33d55555531059dae4aa4ef788a52fbf98a15aab0412627408629d81c5437c50f6b443b420d2bd8cae53e096aadc422850bb4835caa759666d517fae3d626bb230a759ec9b1f73e3fa9519b78104dea70905811c53d7b6ee5aa9043135d210c40cd792de243bbcccc41f46da4adef3481456deb6d7ac06211a8e05efae962b3dda79648662ff13107beaa5c2adef2c2cf23fc8b244c10dbddf9fd19eb181d074f8924e279ad9c5be2ddf6deb0ba8820a80a9d266566dbabb42af3dab4881c7440ca390e97341e53eb55c035fd7c9a99a0d49d655b886b9a3af936f93373dc9e8434d98dcc019a1356f1a70060a38e1d7ef00dede26487ba7b31f230fda05ba2c2b213235181332b5d943db42203b7562b716e4f06d97b28f939066cb7417c25b5956186cfa2ebd657e9641f91382db3daea4ebd869c18af05269b9aeb0e9ed32b2916dec623e89d7d7c1b122ea7cc9a92ed917e4cf022e80c47a0e0364b8aa4c9f3e57842da5d37f505f72ebb4102b5359482f43b7c7d6fb93250894fce69da7814348ea596a7a77cfed1ea5f4f8b3e7cc59c33a11cfd5842e9645be75405b3694ad5a058f7f2820ecb666b53a6dcb2c7cc569f623024000aff55c541e8b6d3208f712800f694ac7f74ae58bd66e9f70a2a25bd94288aa6ecfa50cc90787d800e0e7660838c6df11b79f3b63dab59d12b8f15634c391827553ea37b23094abf1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hf539e641d8a180d96eef6db928be1af4b1928da210c51a7efc24fcf029607c5d8e6cefe2d08daf93f010adae5f437efe9ddf8806db12acffc1f1e47fd3f4b2e9d0e15774ee7ec348a5334b14c9217379bff0b1ea6afd00969b4bb8512eed68dce43c6f951f8f4a177b4178ee33de80f8ae7d0a9f905f4bbead45f5fdaf5ed5fb0441e6ce25646478ab881c200c2ce415dd20dfe277296c00d035bc118af0a1a38b15aa11bb4764b3fa98efd2f67fd28c974d85d7d527e59e218e09b690eedaef86963f795d3cd150d0fe268a64b32d8c0602434d5759fd29861e3bc9f07273e1a446771cdce2691b7a501d1a42a9a2b3c1fc0b9bbf5f6d4dd501c467e0c5b68a301c4101079577e05bbfafaae5d6865d5ff8eaad0f139b557acf46e198b4600586b895f104858983e7ecffc916c349529d993e702b7af7c72dc9e97f7fc958aed824575b6c8d9dde52a3e251f34ebbdb7f75e92d086bb705eaf2657ebe31da895393852f695073d89038537ca75e4fd6dbc066d257f734879f9a74a61f3d9abb5b49850e0b6da1cd0cdf885f652d8cbafe370a73a3b0ec20d736efff6266ce889d32f00fae7a84652cc8c401c2a520c29f4636ded0c38a13939432dccc34252c50c8383454686016d9d3e2030c5f743ca05a585a51518ecda3213bc924be4058a47050eaa9b338b2fa20b1241ee14c95980fbf067338391a8b096dbc6b40d80811da51bd69da0a74c56941378246f7f1b99ca4e4ece22d660295253deb2eee6deb67b845d2ae37c9d6c3d7802c1968fc65193f567380ab955ccfaf77ce7a954331105d9d15dc45f12b2685dd69d591294d8f61b891eeb1b27ef71eaf7100daf7a3c5024d79c8e5ebd91eef63dbe60449f17622b9b0bfe2f2ead58071f9f499c27c777dc017b9731225dffc40c76030db22f20148babbb5af52f60ea14e580e3174580aef4fde220efc2ee7ba26eb78a74fa357793a83b2e9efa0856c4709f3c71113806c529657e2b18e60299cbc85335b3b6fd0022892ec10a2d464c491eb60992276e8fc5ade0d8bcac84b324ef75ad86fdc376d0f0a13da3bd9e172bf179d047825849a958e2d182c7ba7b077f0ccc14615631067dcc484bd88f49aa24cd39cb2ade7aa122319c7cb48a42f6fa46c5e7bacee060030ddf20614adb4cf293d7643e702d963ebecf5a0b96d189f7d298ce51edb3bc010ca9c613f895cef57f5b41a4812302b1d717780f45f2a2c089666559fcece367df6fcd9e39ca73c3feaf8c3972734617ee06bdb3d8891ba93fe4516ab9ac3406b02fba82b62a04d16112e9c7305488926c4a347a42998347229f3a2b016734126a6bfe5193d5d1d563de0a6b183e68c7491c3c821dc5a7c71f60997cc825449396d2629431da3133abf5745b7be5daa5468caa7b3e59a6306d47ca5bbbcd8217448ce2ca78ac206b9ee046a823b9cc14842a482045b81a533014e2aaf01c0fdad0fe6888c25f99dadbef0a63123c78f5054ffa908d623f63a371ab2415af8dffabe4dcef5d43f549795827c4975c79ddf9a5c0c5c079b347a8accfaef8c26c95bbf14f2bdf6b4379aa077923d7114741230943cd13058c4e5a6f1abbb52e9e60e9ff5e5e92ac5b54bf18736d47097281443561ced0c42ec6f847e1a92b9fe6543808f12ad8f4a2e654446fc4de07a68ea3fc2965a7a45a0a66d30cc28a348241739ce2bb9f55090a349594a6d95e99dc49846f83d1f28bdee5370e92b0903555cd5f39c1e47608c4338fad62828acdf2549df913a2301a6f18a84e62b81830e894eec7fc6c4d3db92e59bdf2e62c606bb543baa4496150418c7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h91325b80d2d7304fe688b9970668ca480fddf7a535bcea68988c2b9106cf73808a21671c2e85f13f31582249c0a68d8c07e1b2c4ba6ae5e35962255fde0956e1683ab6f57a6fa54df57f926bc099cc77d23ee6412c07ab6d49f9791697b01c943e32396586e140510253010559f31225b5ab0d8e91658b1dd5316521036d8c31e9d540f120be4c2d5557961f14960da694f8f69000df0a82712a8835400ef8a2020eb8a62b8052e2faf0423dde374feadba8a03f03d04b3d53d978abda4e81644983f085f48c16a35494bb2ed6893d8af1e9558ef0fa28fe46c5bc70fa348eca7b748997b88abf5218ee556343e5a96a0b9336a5b3c7801926159d860aa8915068592540dc19d3cafc91a45a011ec271975b752c6cf91921f8e2a87e10c16681bff8d78cfb144be51e4af243000af77feccb52a0176fca23d80aeda4797dac8b84089aefae13b1bb9f83e522eb7273de85f5abcd8d5bf4fb6aba93355630c412581e1154e5d21224e9cad137c79ee4cf1855a385a995302cadb845b3d7d746147845d115e2affa41107466191878dfe89d3303bff1632db076e672a8147a6938d8a53edacf5ebe1054ed4f332308126ce3fd4d3e1802c1766d5430b6dc615b36100b5b92023d213eb4e395783ca6670e116049ef6ea16c711f3106c144d38ae096023130b3d8656f99c10a3d41571cb08c1121305ebc3d7311acee57bf8573631d53ed26f32ff5888157ff2657820d26be4242e3b52c01a42a0217b6301f4e95b8c67126791e76e3ddb418a87a69d3c61bc0f03a79b28f17816e42d89e16a14205b9b36f7aff3d54782323f19a2cde8c98f44ab91595ce8baa9776d4cc30d2f639de2db40bd46e1c50dfcb69150333eef4be43460b00da23ebc3e65ae2c165c2ba320d14cba8cba666ba896971644e7282f6ee025ed0394b53b09b8b783d52012dab0f6594b09f4f3f8f9a76d1fbb76dcd847bf61f4c27aa40051e441953115bd35c7c0236d46900c9a1b6390c32add12d2eee1d84abeb48fdd2949bf5c6d29bb9db6418a9c7adb369163cc67e21e05e16a2d1540b85f884d5ddf2f879eff9effded1b255dce027c5a693c43501fa4bff2f6782910e844ef9b428ba479514ddf1c5c394468fab946af7bc73c1aded5b5ed9c1544a07797f9104b794516ce7c86a7809b0c815321fdd3a5d321f9e05550825be4ef1c97b943d099dd2ff2db2f7e3b05d8947241411f142a4d5cab213af5048780ea5f0b95dafd5a718e1a18873c3d9fe4d0ed70528003b61cd40bc676715f876a63180758e41f8558bb5725e0c0f7a29f9fb1ce95d4d924703e50379e2c78edd9692bb7711fa4ba4bc6a53c293eac928e7db46c1d74c44b884295b68686e51eb152ab180c14a10208bdfdce6d59eaa946d2aee34f0ae476394e321faab54b5f524f151e9a90d30cbcdd0ff7e421d15df5db5f825b2091e25cb8407b013476b064120bee9bf3a211af3288a8505cf718c26ff458547ec2c0a6a06d79c2a6cd10a187beb8c06cadc166f83e48f0ec82d5ce50f9d24bb854d1e848117096a478ebfa3b22a36ed09864f4b59089962cba9851b0b64632dee8958fab4ae97a6445bc930040fa35707288235e09bcbdb74ce44179187ea4132a72c5b3083a207489b3d2e7ce948c941a8b35fec022dd436d802cc5d5a4e52ffad1584e9cbe22f6d67e15157a25747b5efedaac28aff03fc4222fa30c74bfa2b3cdae01fdf36d2eda4865431b0dbebfc04da21e54d94d1e910293aa7e45be0f6a6a7abf135d864989a44d235cee37e3175c62b53e01e51b64f1ae97e6f140f565d2b5b5d4d5e770;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h710a643bd739ebdeb6b3b239fc1b75639dfc287278248257bf07df742a644f4ebebc595efbefbc8136a486c9da4b1f0100354b950f116c20892f1ba117f78006c256dc6f886a9b95c63af5ac17db0c90ca9730709f0648f28b4c9f44389691fc937c67858c33329e5875bccee0e34c170ba0ac64bb44b6376e6f4d76da2335c7aa10c170562e3b32634626a93110b636ab02b1e8299147bb7fa5d8a449e1cc6dcb4d40c200e12a83f478cda49ee38b0b264fae4de014479a8bc60ef7eacb9cd912a4a0c31aa42021ae3008286b6c579c9a5eaa7dbff4b767e64b0bf766d918439f6ed9a021b7bb22357228cb63188f582369882f38d3b9869e9b3680f381360711e2f65c9314a847a06da98d7687f1e03c911a5ef78819a385554999e5885f58c77607437296cab9350dde918a95705b6f4e11b1f3464106a591ff0525c52e8b2f64937c7b6ed3f67f781ea6349ad6c130bccaac3d89e9287e94808102c759a984fe59a073c8529c3bca4e48b99400973a48f671d9794f79ae575a489b4ac8006dbfb2c0286c177f216d8b5bd89ffca876adb146362b291217da11ede169a0cbd8dc19e08f505f0f680546428070b2892657835e3c5eee9dca3d5102123b0da5880efed043e0dcc676b27a5fce28811e77440f82f03bafb10132f4b85917592a6fdb1ec120812e06a0ca0a9659b6cbf9279a6a8eefd99961432faba3efed6f20867cbb427aac989a62df6d0dae1b317399a43a8c433fe848c994be8c23bd52221baaba49f0c77dc85551994b5ba73ec218957854713506a7adaab775f251188cdfbcce2bc7764a660d12c6704e3c830c861010d8067cf6bc57130c036b27571571e59148b7876e683a73c1913d067e9d8b557f85158ecbed4d347fabaeeff0b4c9b8d6cc7b88934b7142aa5ac03eaa6b992899004f5a575f8ba996756427c05421ace23d5c71ac035ab3985a558860aa40641bff43915b04469cdb81926aaefd5597c74305c5ba494cd555fe2d6c3251a7efecb786bd2fcd2333b3eb38342d3be9c33202e622af3ddc50b8fcc17e83ebe1f91285bc0a449798d87790a0b2dfbb221c515d92bd37d44319f44b2495572cd083e82626a3a398945498289f30b80f3d6f91404bc247e6adf391d7ca0264594295c2a6ca1ad169cf021c4107fdb43b2a67047ed500414cfb66a10daa99fdb0c0551c3256ecabfedf2474d188f066ad646f4ddbbfb66815aad5fe40caa6ea7ee74d0164383ffb09bc2a65e2a6c4b2041cfcbb799ef8edd7fc046c0dbb9959e00b413153851bee53cd53343f814a6f0fcc3749007a8560dd9359d1e5e9012fa68c37e7e1b73696ce4847b083fc52f0d873a497300eef08f5d89f2a1dc607d0e39b86916b8d47c7cb00774031609f4d0ecb73abf2149917459154de169d6ef37e2c6418b9b44793c4071e6c654048dde1243388df3b4e6a5cb33b27ee3640587f773114ad3c9b947e82633bf95f7781b83fc931d2de6e19963e79900b1a7aea44888c45aea7d9993b5669d70f457035746799ed9b7dd095a7fc58f3867156b9544140bc0d0e877350912bc7748aedf29e7ccc452c1ef040792af15073aba8917b411c819777a4e5e400cdcb698b9b2f3524a0ff1f94744e699b098b1cdc92ca2800c80f1a0fb0c37f121c8b0dfaa3c84d2a4f61b9f3f3e16864fd03b1aed74c8803770d95967a6360f48eb95cfeb478010f2e92e7bdbf28f5b021a21eeb92e1788c5914ef11c012f7c8bc914cf32fc7d1713c74d072ad8e7a5df23e1a8c141e230a5519a31336c2b01c7b8d07f568d1ee76eb8cfe7af0e1f88ac92aade647a3b3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hbc083c1a4192ea7910d356b7add4863e6b04dbad3307cf665c7b386f10bd7d64f4ccb6bcabf805b2bcda6c77853d237104156b5affef0b565d18beaf21f5f3802ae53c435170a65a4b54c03903069be80ce7605a1dcf0a0c61bc676b4591fa857dee6e53aa9aa52327227e21aad78d0f3274807698bf8ce121ee49afeb91a9f682f0d39026fffa0cecca89ec15ebb304ddfa618450fafe769aa2629c76bf15a5fc0b098063dd54830a3a97e71e42c51dabbd202703e06a18d4e00ea27176fcf3e8fe93ed488aa8bf1631643e730668f5846dc39ccc14d1a4ceb4ef7938c55bd05bb196b1fffe02ba24f013601fb857d32935656b1b3500c4fadd281794f589dc92bd261f977d35f070f7c80c12be825566211159e4c499fd6d859f489dc6727eb0ede517471fbf6cae840369f438d4b9492d2ae40ef06377278e58b90c22156696683b4459db894d12f21a759bd107b96aac97a569ba496460a0ad54fab135d7d47c7a1d6136c2bd39b5156b21938b33ffd12fcba765bba8e3384faf591dd0f511fba0c2741f044cdab6f04633fef0fd4a842d3f1b4527b8772f891336de6f08bfc6d3dd9f0d7b8ed8ad94d47c0a30ce77598b21278841212a8bcb3eaea534de1097438588af8bccdd14e2e497eadfbd31776712dbf1da696e849c82159861cc710cf3f3f82184d567ae05d39d0dda69e3077c0255435cca1b94eae628633d4d6cce7f91637580092357758f43d61e1eb2ec5100d35bb022b4db4b12b924fb79848a619ba8f2f8b843ebd243939305316d1f086147fd7d56001710a5cca72da3e5c988e273391b3436637fad65a5c80a5d801ba24c953679dd5416d1ef0e1ae074fdd3fc51e284c497d2785a6c7e8d81d9db49e2bc6c376aea2992b9f6c0222632b4872f5b0e443e103e09b8d29dfd7b68beed474ef5b895c3390cec2eaca81371df1d65781a7fbae38668a5972b58b2ee9e2eef65f8fafa7b4c8eb07941a57601f831e172a52e1f0a7db14f1219ae92059ea6d29b98f4d3a5af399240e985c2b2bce17514ee0ac3ccb3e2caf555c2dbb502686a2b94d43c5f224c75e9ca4151229117bafb743174ddc6328d59862c8c8372fbf6403bf8edcdda3c67da35c25d911ea202d6d8dce5c13deb487a26ea4c65fd5d9ff9de50f6d51ff3d6dcb485c3c07fb4db5a48bbff22ea1e93243b6a28f6979b65abd4beaf25632551fc88657bee45ebd5d7079dcb3334e686b22f6dca6f65a411620d81256c854a3a6a344fe478eb55d13c5d8bbe1a6c0d2b329668704adfc01abde6199be26c3692f6ff9218f1f5f8168e11f75bcad43c49b4121472e44e42b8d8df627c98928a09aab18a4cb2477458e9c7fce1250de48a29f67886d45772fd597e9f8cbf88b0233dd9fed38055487b78c774c7d7c07ee30b7fb5577af6d78917a809737e0c0509b4fcabdb6de7fdde3297ee94cadcd5abb16a85ed67b0faa8d11bfd479a44c153d70cf348a8752522dc5ad80b18e8f313b1076bfdc781ac9730ebe5bee09cce7631952533a26aec3f02bed621fbce27851922f0fecdae2d178e61f418df64f879319875484a16962b6398583b0647087b8a57ef897d2e892062a9b4355e512e0ae823590dfa898efbe400b156c0502ec24e6cc1502cb2d29428f01f656da04368000f7ee52a9c11168e4a39f32fe8a2ebc2a8b0573f0a31a383019e4369ae4968a3e2b825060b1251ef7581088e5030c235782729551d8fc4e3822b60ad79294c6b0f64a1587fed520d283604cd47bee8299ad671c45b53d4c06316bbdb309c63afe02581e20f5a1b70a8d88433a9d4cd63d795b7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h27ae01a09c72bcd34102d0f8abdb3a22921439fe3ec10ac60d4745eb8bdd6f81528e3383ef72fcca036df00674c25637eac97e2571a83d49d5ade4112aad392b6c504259b8e61d29b8a8fdc4614984ef6f6e5d9db834949831209b1581ea69c98ea285a9b1d121eb65afe333f37703917e8db0fb87da12bc57a085c9dd18bdf2ab8c02220a081104b82bba501ab8bbb282702ba7869f70dbd700c700822d9d49f63664509139a8049e71691b5e3d7b263fa70a189714c07dc5ed380b6558c87e73578fada33828f92343ea14ee3d604811b1cb8efffff7db41c56615586135ee4c355fe70a671bc952737626dd8c49d3057e0765454b32d881e6ba7289d6cbb3f223bf7bda14e659742e077c749fea9fde5db1ba1a8338e693086ba768c9ccdbecf85156f28e0a73e9b9b67cc7c4ad6c7422e405c64ddbe0505e07a0d1c0a2c89a262701194c27c83bf3551746def8a4f79332f1a37f194e7350f18421c1371bb191a6a817684b6bf4b7455182a2329acdfff93316546fbec5e3374a316d87ac29da62af1f5493c8744b069dcaa1d40dc4b33e57bed6ada8ed45e11f3f09dacd5e0eaed85276a746c2bd799a4b10ca1710b236f3dda58675401bb787b0c45fe1404e9de9935336a04d1ef2e788b1ba89e460ecbddb99cf4339ffc7440a6f8744e98d28c9717b3af9f2d4962781435c187c78c8d61f61fdab520ef31823f0b1251c79e84d5e0d98cec0b3892a801765dd7168dd0260e61b281362a4917da6519243affb94287847693ef45e7fabc3f602fe04e97c1a6e7bc99d5a2b8f9d92b41c6f15b00c95a974bc984449e1c542d545657d35bf057367297cdc04c34652494f4d95975ff81f057ec05d2621c5a9367d949382a07585e8125e1aa500034c3b765c8d73ba4025889865da0067d4f39b238355aca5305cc16b6483fffc88d7886f90e0484fd634aa95d71e2338b7224b7634b8767594593b5308a010149487a18c64896de05fa87f2e25f77564ce7fd7ee456a3b344b814ac0356d44fc02c680578d61268f35f4ab5941cb53a2a60add693aa35633ba26688918c165ab6a07f9c051e6ce2e58fcacfc4df9919f3dbf2aee2e51eab74147641bf01e39b17eb5924222ec21f21811545119f7113ac19830efd7c8e4abbb8ba572bd593aee044c1c3ee1c77551db4c46316d880af79c4eaeb9d40d6973d63382bcfddeec91bfd139477bdb7fd889d778e044793db259a45d02aa4d080c28a78b9f3fd1b679bdd087344a2dd9578a838709527d1fc979872346470f978cd9c1335a70ed4c09a393b92a53bc716e598b98ee9ed5d0a69493804387644a1b383f0f8fbb275ef587fbe1339c96d0fed1a036cdf3c7d13740d951efcd9776779b3d9138bfff8b7b54b5f52018742b98eb0846435149635cec90ac507b9cd77c2b3c381321ab6a173bded794683a7a8fef16be02da68e719ea7598610e1b6684d2508ffc0ca74c48946c63e320c4ad6327a2c5dce104ec368be42baf595dd95a6766edf5605e8539cc842f8cbbafaa2e881f925de7495b42bff2bea1f59074235f0c06eeeb9179522b68155b165a14eb333d1ca7333b88e5e7f570fcf38b520e06707b40db9f79ad8b8b25256d3a9e17870e80ce11384bbd56cdd35ddbfa6fc6e1f03b0fb2ee9bff59e5b590e3c7bb06f8d3d0955fa362e3713c18582c58b602aaa6c01315f0d22a14adb485ba4c44c8429b1f87d3e8c8987acf21d35790f2724a232d3294bae87e0471dfc7b1e60e3bbf79093b21863769f2a986677792a4d484da26dab13058b64c557d14b98f1c7690f710f922482158a8253432;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'he9de75935bab3222771712f3186f92b7576cc82fe1f047e3ed383ca7ebfc1451a77ce90fade787a486a7fe71cd38cd00d65ce3f0f0f9e1dede5ae068e4297d2844ac713c76c4885e91de8ea7a2e0c065a1323f883af1488ddf08319c9a8a9f8e24738f1ef5fe20e7b2af599ccbb4f7557345e979acc001fc08610881549c94af7741f56b7193ce6818c266c75b594cc5a007ec9b2a75af9664b0db3b4244489cf3316fa7d4c699574606be7adb265b7cc59d0a3754869e667c9e3253614cea7dd5c022345dfe2ca82007360be7dc8dde5b22a22677454a29ec5eb015bf9297c32f258f7eba0afb72348fd77500e22ce7b2f7f549da591080549c02a481634bd7abf92fbfea844229beda386027c849a1d09fd9eb5de22318052b65e7e7ffad91b097d0b42258e27b01238801e62d2e19216a1a66545962b8b4f7a32eac91a920b91aae17e9e0ab7e2432244e86b017d0af5edf2cf8852816602cd5fe62449141cb89768066348f3b049d499d67a37e62109bbdee1c8217e9ff8a33326a9ede31b0fc2d8a52053d5d7dd34e4060f8a22e8a87ffc2a4753771ebbeaa92fc141d1ee3066ffa849bdb50ea9578587c30f3a7189b8b7e57b62c266e2f01c03f74a945e28fcfb39babcd430e599950343c23957dafe925b7a2f799b365d8e70e36db29d11a1f236094da4f8a424ec76a1180a09724bc851424c477557ee7ba5bd1fd172db878338614062c9b480ddf3ffe6caea5f079361ed0d98d10a94c706ca17782c1d8d8323b53d73f0b3f5f65d6d9570217b485491731fdac4ff0a2fc09037a21c84a25d525a1adef3636a5fd44d12f2cb1e7e7c774cc52b30a161d688a1283ce0e24d0193b5e01aad3a394044034b56bbc159c5375c6a820b935adb9f177e1515ab0e6af69f92a9e9018a0c1196bcf4b8027874424ea2697177b12d37ea691feea5ad3eef581e5299d74d50f9b5a53df54c9856144dc110d6864c3e67bdad04bee967a1546e695466f315a1052426176fbd074b8936240c90368d69d187994b74dc1a4956d92f3e86266ec6075aaa6f837868d7535c0bcb59516d078366ee28142c54142e2ec715db88674bb89a489a3e3e40de0fff2ba19ded6fb42b2354cf9e69cf1d2142306bd1a3e839d6ba9ed5cc8e8f05a3106854740542ad87800787e9d56af128660eec5c9e6ccb8544fb77c667496320ecedc46fdf03adf9fc595a97cd59139645a44b518f80c73015782a30f6fd6b7e88cc3bb0af9cd65973d8b800954c2d8cd1a0cf2fc362ecf950b27c5dbbbc8ded764fc0709ba2e54517d9600870d0de9170f78479e669fa01b48b5463a827fa005315609ffcfdc9c75f5e6dcc203e875199f666d18526df2336bba05afbd959711f3019847999aa2be4651e077b6505156e78b797a1e6f1c03057e4d82697fe878a4e994d3b1c5b157bffc60b35a9f0f9739923d76c8ee476af3f87523d45524f37ba7129b9e27640bdc352fc749acbec185637c19c22cbf592ae839866c39c010f7874ff99adb7cdef5842c590458380c35ed67e7b52c29ef42a1d7d2cce4c3d70463d292aa368a21ad7f8a68bb71b3a66e6c3f1f6de919a79f313cef755b348d1491497999e3d03d1d6bb9cda8cbd10970db18ca9ae53d102bf4f5b993cac58b9e9b500bf3ee48e8fed41fc7a1a30bd998399601804ab62d8e3c673ea83dffee20461c1bbd51888834c8a3917993925105b3380b0b1fb7465e7cd43684ebdcac7fea266bc0b27996e309ebcc50b8fe82c4fe1c8ca0702c02d4b5920ba22cd2ce2aab1a2276f22e8f0b122d6a423aa253d65ab091810aa000e15a67;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h45a7bd3fb84e1ff18c3cb445383dbf6d86fdf2233a3e96b43fca2993a853a4a8e8fec336a0068ae2e9dfcc64f3925ea3bca9b8636d7f3eae82b600c45b54132f3c2c691f5b2d902ccc061bc0bdeadbb196c024cd6de4cb57c0230f5b1502a469dd4512cc7b19cb7b480ebe5dd33227e449f06847f579c82e097292eef7a08d13a5dbff30213cd561486cab8fec97a0d1ae84cb672c7799d939492e52e3c2760d24b99c095a72e3767aa11b7abae34c6feddbadec18386b2e1f97d04aecb5b69f9a45ef57c62f3ecab7b845efdb22058c582859a5a8b209e0737164fe5079c376b0b6ddaf3fee0308dfe2a9a9db08e0be89602436e25655704a12bb55d4e1d5a966c09ccc53cbe77e81760217b40b50e704a6938cfd29176571bb982bf55a544b331d569f2090922f2f440d24e10c09aa71608a1b0bfad9c9222c8cac84e3544da0352b7a4f9cf3df8e48cdf1cd8ca6b2ed387ce14c7703926c7ee99dfcc5e3e256f28ae73c13a2542c7a12b95560a52a3e09038ee50b16ada8df628c7c22cf405170e795027ba095f8f6a5be94eca470b27e2b83137b2c7cee365bfea98a493ff25debbb9026dc493db7adf613776f024b9f2ca3fa5b3a2dfe8d469d2446cdeab2c266b3914ff471467d0a716ec2fe8fa8c40ae2e5b83cd7bb17292cbd114b3a8a7d1bb992d7086f646135084fe3470a642d690d6a125e2807e958780efd8fbc3a857373829a6467f29f821ef32ee4d1834ac4f41a734025cc51c98a6765874575e8e02f9ae940f36839633b8c2e4d708c54c98cd49de8d0c9c90ee77b1cd55c6b37bdbc1fad7c2e73aac6ea61405a36a7b1bfc40ffc80eccee9796224a95bda5dd47cacdf310970f0c67badf2a276f60810602fed290ac99886c3d6b484165f09d4204e9512a9ee0866caf35d97f4024b068a92708b6084aa8730e434280dcca3a438193882f2cd1bc1117edfd477d37e4b1c289d406b9ffb8e15fad452456734c4107f2d0139f42aa0ac1f72db47d859bb17c0951a681e83798a2fdde097b9c7009f03893dd3b62465db2845addfe41dc377805355ceace4e565f7a89fe20409e96a7e76b79c92027bf5c5cd4e1ae2d5ec4a54b24d1df67a9a7eaaf2966be5b38dd6b09ae06d133b3dad97f1bbf9c644c12937fa7262248f07aa3be62896108c2893e253a8daf1e12f63669a5bbd3d2483789fcf1f15321d52dea0e3715b0d6ca3cf61f1f66fc3a6fbc90b975672ed1075210fc258b07ce3d0561e2e9d669f78a1b9c33ed733566e74ed67a0ac25f5a39acf31809f4057c31b82faa7d7ff4c9ea656bb819a5783d60c6d48166b4b850ae00404efe0aa9cf7450de2769824b14bdac8b3b4aecc6ea21581ecb89114cf388aa8406d41876dc98a77dcd6b3caad51eee9cb67eb327535732f618582d8e0df95e40840d1905ebe8a473046561979e8cbba62e39f9d3865cd42b76d2d6df8da7b50f529430a2307b1dc9cb9cbbc59812d8c41fec0a158e7b5d82eba2d403874f3cf2c5e693b5ae22f527936167cfb7652f2aa69e0df3fe7ce0efa0d8c7f29eabddf1b60243df01fc0983265402eac086040ff87ef208e4a50e8b07cf87c4b5e870b96b37e6a53e465e6b87e6f199cc26b52554dc632ab11e35caff26a1dbdf9e295d30a98e010507aea3c8ca08aba7885514a8a028bf450a8732b589e0a4d0569f46b6b4f41ca06674ecef0e528c11e9cf05fbfca0e94e91a24ddf85842a243cea0d2edecc82da07344761c557baaae07252a459cd91c6a71cd76a917893ece756ed7e855a3cbabaf3491980a2e49fc0d3654525c52b0c0699e3c1f9e83b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h7967023572737e8081e180ce6e64ae4e19084b25e49b9e770dc36a907d27955db9d999ca1c4b8aebe567a2d71ec4e84c9ab19481f0156c32fca0975b9d1905157a342ca346b6f6ae6e2fc1fca32cdf6fa7d51b9268f047999a754d1b3f6017e5398bd601b6d46d543cee8b2b39b680fa4b0865527c12944349bd94bd75d12c4a158eae026607a1fc9b6931bf2deebaca93824ff71db893d883984384cec1bcf4102f895c81f9fc18730f0303aa39d73ded9e278b49779e869909582852116095098b2012ee02e44ab83a2eed07554f36b16ec7dd6fad70c6ce0116d3cffd38dad682f58b701ed5e227350e7423a6b9d5f700a6ecf503970c05b9e709314c133731c9d92f09e9d059270d1ce3ef4db27c7f32fbaaef7c22f6f6dc1650435e34293147275a81e41dcd00bec6d82e2e11cfb12eb4bad6ba2d56797851f53103bd85fbedd2d341a1fb40f26dd291548e511f6219c444b3eafea6ef742a6431f11b5a999c3eb34e8a7138c8704101d05885cb35d2ffec88675da94e21f6e62536cc53957c68c486d23885dbd48ef313734b4645a0fda8488cd3a08797d9427d66400d3907b16fa1ed8e7eaefcd20ce5ead7f3b29d4bd4841394ffc4d7d0b494f93fe6e60c9756eda7ea345e9c1990b58ab51e33b16b9903b04496a5df2b62c9a2620cb4fef555af074458f1f88a0d922ed3c64953c70b920788b1b5552fc4070714bdb402a185763f4eb1e90a85ed2a92e4ea7fdd1c4bc5893caf69be409cac6022c2ad1941e97728ae0684ca63e1212aa82329e3c9459cb1f226666766fdc58c6913bbf4e05182c0737c5575985e7ddcf28051587b5edf96e7249c9748b7d13dcb7608de2d33112a543e1736cdaf193247a07a11493ba88b21f6c785a74922817d6f1e9bc07bc82f5a26b2c4174aced9f69ec308154a2ec56dc0d7d4f644a890b05c245953589f982578be8839a122cf1caa7b94785ef6da2b53f70f59d15c7d5db5cb075e8d0a8c01bf718a2bdfdf3255e40d95aba8889dd4c15e95cd8192d08b7088fa73b99be29ead8f8c09dbb9c5298433ca70f347b0f339784fa2da05b12d1591e374a28033e8349e79fb6756ed3f7d04d4bdc1326e1614188906285a7d3af16cb03f1aba242c7cd1307f6893a4c6c4e6e5311df63272c1929697a15c5f0c01d2936fdd391cfb506fa1a459c6394733902abf14bfb65443b78291e07236e3dd3e320696ca5f76983ac0be65954370edf429fe190e807831b711e5cb9f66b017bdd2c97b164913d8d68339f9534e5f8747fce480a5a37dfe6dbf5b6993845abc60d7fa0315c721a796b6e5326f912cec85c925ae8c01898f6e0efaa4d0d4e3b27985b973cb255b062ff30f6586370dd5d52c9bda5464d9cd3a531ebe6fc4cbecc6b6ca03f717fc00c082daaca35a8544e59471af75a25673b7f11a0192ad49d1d665c93dda54acb0d51513b8fb58bfcf4b22da6760f474da2fc9dd965649fc4b5581aec85b255fb36f062f131532644f706a662c9efbbe8f6e8adbde507e78024a0ebd576c45c4b891df2c96dc518dbca964e9c840b7fe95b61558ce6568d11220f600aea513cd52b66d74f6f097c71657067c117f16f5c80403ca4b10572cfa5e911e303c75455982ee87ece645f6ca88a2285e7a8b154bc71f8e8e2bfcf8a743ff87ec0abe237b851681f0ccdc55fa694a9ee84f17ef07482089fcf09d64f541eda128ad42b23b52ff82011cfbb1f6920753a111d485375b74b30c5641cd538749e99cd56a266845efcc46ef5fccee61570354dd54e216e168d86a7958a244fa0ec7ebd1e8281b34129e2c0d2c7d1b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h412013937aa8f6862923ace14a3c0f4cebbaa1d03947adcee51713cf014e9d04d667fe6d0826b90c2e547af8aab2d60ed37257ec223569e296890d2c957115a12d003e5b8b688dd3777cad809518693b47210bbaf6fddc8fb16911cf818ea124e8281b0b9d72980d5f47d82c5f134453ff6729a83c5ab97b26852f96d8993bfbf1d39c7eb2d8e3a01edd004299441f79629f8fe4489debf93b253747ca60a28040fa1541c655313cc4c48a36c309a61959961ea67ad745539a8a0cf0ef5d5640fcabfff6d3db547ee986c128933a0d9c78149d08b11f4639e39933c44cb0e48c4365ba5e756ab364acf2c965f7d3c8e85782dac8e306af3734c036bc92fb6c3a9c34a9f2e3a3249f60ea21e99de570860f3b75b18eb9040e968f8a98a09cd6c80f9a44ee487952b4070c24aea8d82a2349c1fa32bd82f4b3a5439b7742332b5a93174a2a1b04dfbea1847afbbb94657256c530ffba230bb0be74a3e4d1bd6f0b0ee25530cb9e04ec4c0de4aedb0784efd9cc80b80bcee98af8e57e0ab827e53a01c78184edff8fb7a220f0eb9286ed52a3bf8894e928941889e9e74202e427b4b99b035e67eee2b8dc29e282c1a5905bd63b8369dbcdf3a5790ce33bb81f915d11b84d1265fde34dbc84cb10afd6f7d02947f0a67ae6c6c0aa54fff072481faca0a3e881f747e03c89778e4b1cc923c1c3f3f047b5f7457c1be11505971f9b23fde12f49c04b12cc0328637c985920ec46fc855aef8dcbd38647e135fb1a13eab7e8500f4fd9f31e6d20eb7d1b76050c427843d8d6bd58d5f68b7f9b65646f2ac2dab20a8a49aecc215bbf7532925b018a6d531f025c71e88095a45fed9d9e05de43aac7f3df7b727ec40bf5d4e5cbac5469e9202866e245c68da415521770d4cde46d510cb9febd898f2f9f0af85658bf73d774a9b5ef42fdb5da24f53c587914d0346fa0a42260e381ad739307d6511f8171abacbd3bfc0d75d85ab406cb5c226e1ce34d1f19008d6ec691b533e61e009bd19211fd95c5e75369b93ff9c48165aff51066a51ce582cd69c14e527544e95353f8a77a35d801862817831c7a19aa1bbd881658aad354ad9e6f410aea9650158fd6d71ed4fb72fb120358573c69f950383ef7b28212adf1f4dd2346d6481e81f6b2322f144bb7ee3723783b50b5c4959f873191dad97584855ceba50f48451decaf520722e21e48405f84fbcb6f9614662b536600509802af0685385dc2f710f55737c0ffd43b2d74796b83bf65116a8119f398e75a9b34b46b2c05d1edb0bfb18c6da6a99724a3a501e8f0bd08a7de2ba450a55405ba6378c0ebffeb07c9ca8d2df228ef2552156c819c26f66aef4427659ecf2e89a47f89f70e40ad73ffa9ae236cd453e8eb8b1a88e75631b38f8f241e74c065ea031f961371f911e9533e740b1a56966d6ede86d6f0355f0500587f2e05af24f82c0102c759293cff470764d9569f2bdb156e6204bdd70e93fa0655cda60fc806d07bd0f7f06bc2f072e0ad63d35ea2634a3258a4a462ec055e0bf8d26d7508afd024b5dd6bf1e6c8f6133e4b6edf2a8aa9e10f36cdf6252a747d8ee8e71893f6431cae50474ee63ae2b69127fdd1ae2638b1bf74ae53955edc4f4702026c9e0c392ecb7f16641680bd090dc805b05d56718d0649c4630a699e4e2ef89f106d5c4d2325b4ffbc9cd5b3648ed53fd17a444183a02e2efbbd82c08f69cb65e2ef8c2b09867d52fe6c38ce6a8028d6a801168109189da71e27b8d1bcfd86e1207a219ece246bc3bc3c01eab2d87e5e3398b906a89b600eb7c2a0b2646c5e20697478cc80a72b151ebaea;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3c69ae2dbf3d63159d41f4f4864b06e00591882afdadecbb82eaddf904a3fdcf4303ee29ea117757d91a237c9cb2e11fb497b19aa40f65c4eb5dece00bca421787cb98bed572aff1c8ee6785d08cca894cd3f3040bd9dee13ecb531ddf410216f692bc1e6b3ee4b4207e804cd89576ae54a14ad50f59540348fa1fed5e90f75c2878377392779695c8a5ff614adca67c8e84bbea35e1c6370582be8bd42e695a498cf10f11b9ae38309c9abca2a961dc34ff456ce1ac60a524cd5c5057582245adf39a2e61213c47b335aab23aef7cb89a9bf75b570066ba0e4e11aa21575ec878e26fbbaa08bd07b9ead5b21d2663a3a86fcddea4f22d29aecdaf4a1ff94a686fa46a154a8861bcd02ba638d1a4137deca0c93ae09512fd2e7d3e8c122a9239ddc43e8602da2859655a24d1220fb8eb891394158b09120f2757b85585600dd50331894b61592830cab100c5a8a6905c9042d8e654e7b48cc072380dfd7d1c0491a8d1ffc573403a619b59c58f3f4b9d29463a3a97e41228df9eb9bb0f9bf60c1289aafdfbb747309d73d4d5ab94e113bfea699c7380486154b4022efb3b0ede0180a6d10517a75ce7bf6976820605cdefd96b5584f5bb648008aa6469c56b51f2caab60405a404f958e115597dc7c78cef5970ffbe6cbcc94a6e43b073621744bcc1706da219edc9ebfd516e4802de8a42ff084f27bfc1a5ea9f2f22840edd61cd045863b47ecfdab0d81ed1b7065dcf4febbb4ab7c47d7a3bb59c5f138fc6e3f41e529d6d090e9834d56ff5fb83fd1ce8312410ef69d11fc75c2e937faa6d4f8209c6cc262937472dd54d93694aebaf2e55f988e1eefd3df2fee6989503cfefcf6b644bb0822ca69afb7afd939d67fe084fa6671c86fc2829c377d26d3feddb5ac92984db98257fa278bf98c92279f83fd39a200d259f123ff2ad79de5d8f95e41836d60157138f4a573757db339c8813c2b2ab6c3330a8a495f3dbc07cd05547abffeedeff145bed6b8fef5dfbab2f5781d11e7bf4ec7bd7c2ae14023d2b164fe21854c5cf9e54903d0b3f94c022d2154ba5aded4917e37f763d135d8de2346f8c52be8c6b960805a89ddba5f453326048ce77ee33f57816b929fddd79947d9957c8eb6f93b8a289417bf2eb48536ffd728dd6fe1ebc601629f9c2477eea48b0676ef9f8de27e8ae04c7a1b6fd6cc305e8d0a83faba41dafa2f7f743b0e08166cac96fc542ec8053632091e61cbf3823e941968f10713ee47e73737877424d47b4a53158ac589de43868173d2cef42a875b66624d4e78e78fc84966b959470de2d3ff49073bf6e4d783a87a5ffea81f9d77b7d6fb15ddd44c1137dce3f761bc5f592f540e2ac99acdaa6be018f4a629dfaf2d05e4c467de2a63fa97d5b82006bc893784179940482f817ca93d147920ad358f91c0c86da73165a26b9b40dd43f40c385131db2095512ed63d86b50b0157ce426b91f27cde556a707a0239f9efaf924c3b01219c652746f38b38e5d5adc835cd0a75de615c6699ff63de27ef38345b13f176e78cdccacf3ce109eec95181518346323b6aa175444139552b76d9577a06b644ad9d570277335957a31241f3244837d03caaf69c7f20bb9bcccc935e7ea62ace364cc582fc26698a5ed041c095ab0f1e99777498a735d552a4165e9001c327c7e6334be27162611d35091fab143529bf2e27ace1a35ca49f115add45870cc880e560f9d4dd3b8e54b2c87a53d22e03b987b7b4add9b0aca2ad58c5f692964db140e487d523395aebde1f37605ae9a8829c2aa4375e02ba71f40e645b9161d1e103fb04f54e2d5b6e7296;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h782567944f5188eb08a21a97229c670495132977b5ce4146a579e835654db6de4cccbcd1e38f953ff5356bb8100695d51b78e00bf4cce94743d4c04c7a03b4481e4d89079fbf5ddedc5d039aa3f30f1eda1a401c0488615bcbe591388db137df2d29d6ab5f52b9a83cb9d12324794a023e3a8739171c78bf99d3a42160c3a9468f7bc648af158266a267a865e7adf9f946f78b9c0e99406f88f0e326ac9fd233b2dbafa6993315ca9c1eb9a0c01ddfd7f50659d24ed732db988157efef5bc875be5852c75ddc861280fb68f2087044d176864003ecf7f041f815f30ec4db4f7069fae16656b86ac6464c2b6033eef66bf9d8443abd741df5ae0aea2c19c255be19c0bda11a25e38773eed16729c4e2d403d5a423cbdf0f622e03824262bf9462adc24a9f83461cd2c8fdaf0ccc57d7009f4c978e0df96480299d6ed016849aeb47a6e8f0e6c4c37a6ef682f13607aee22f21ffadf7342800e184cd0c5ae47fc5e93e54e88c83f360950296ba90da729aa994e03d17c566aa7c8c154c13841cab1c1b4048b35c27d795eb37b34b603d86e8156174df43ae1d81e88c7e9837117ccb6a23f94afb1e8a93e5327b5af62090aff72fb8768b031575bd3492c5bb6bc75bc01e5bb751c204ab99b25141a38181df668ceb9c9b6b1ae9b10acb19e04483e61db99da67790821e670f7af8cf88bb121166b350ef00418fa39165e2e556d843978bd647cf8ade91136bef5aabab7721271d293f57e493a33a6c1c4c3d1af37b8ec36aa7098266c8fa8f361ded01da0e1c6485db58f4b19d28fd02e3d08081ec87eb77ef531fb5190d2e47f6e0f1a3b5051c88a4bb88a6a80ca00eddba7dc022a85b9abd15782f61fe8f8e82ec13669832792b8c48ceea2b3752f5b61aafe8403f60eecb5bb612c43dca2ce04b28b622cf52f5c38697e630207efb176f82698cea295d807ceeb9683a1400e02a7cbbbc11c12c0852012df4ebe9f9b716c4ca063cf5700d46f161d49f3691c9186c023a700b3ef65a4988a6272f75b6a57e8193f64dc2d1f16535d1b092d826935fd6320e2260344f9ebfb6530e0c2a403c5c07bad1ac7ffebdb81342d594c0832590c03bf6e3aa106f7b41725e3bd5973f48198e8dc9e175514733b1397a363368e0cbe3d682f6791ab7b02118cb1aa2cc62a8aa041193e5c4af39ced497216b92fe4eddf42778ecbf8d3f78ac044b7bef74d2d0fa25f9a5c222052d1c51aac508e29c37261fde6a62b98725b02c5ca09bcccb9bea20579a783e217cc2d32638255ea203a1d1bc92ebb434cbe0b55848c713e21ef5cc5be63afcfb3daae22ec8513edc90a716a64560f08271d3ed8f7a3b86ea31b1c07d78139b816c961e15963b9763518ff7a5e15a2dfc5a43718c5f5a83766161615ca0985bb1be3694894d1c3a7464b0037b6d4b707b8508d0e5ca199a5c05b16d3e3006b14f6e77fb4782b53004641d7fa6a047768e8eae02285facf439b20c53106393d3572d440e6f1784ebcc04b540eb14f415c156748130178a1b231c4446cc0a59b3f9128917948d31a32e47417e1152a8b2ece3d87cf31e9fc4fec34e7277693cda64fcd001a06eb17536301976e8b8063a6870e54001c35837a7a010b3dbaaa3d03be2331e9ac9140c3ccc177a3d655b80b66cba415c40ee9ba959fec954c3435f28014725d6d555607552f5b7072c6ff34510f576ed091b5bce9859bcfb51cf03742877cff661b97788d5c0a61e39585b5ffe601fcf739d2622e158190d479cfb79008de11df78ae8c24f495cf543dea13d10d61e97925c47c45e1a65b29c05beff43742c9de04eaf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hbad23845fb1544556cf11953d1e03ccb523f4c13bb0fa61c4e092f2a2a907f9c51aff8a42963e741a0a28a694b2b4a9da1d3280741268c34d99069296d28edde2462b271f18bc63e96a9722330f1b926e962804145491b6fb93479d3771da8634462f746b7071eaeb0f77f9846510897606b6e2ae89ca3755d49ae6dd3f521ce695294f0c54798eecd0e9fe82ec0c2f5309864ab5046369bf62ba5f4ec71aa8eba7d177df623e705456bea6d63c6b9ceaee340137e89cc5c6ffb9c1b56db1165dd085750c4a8553f34845832a5dd72b24a114e361c200366697fc9ee20541c063765b34272ac6c4c7427a41258c7f03403438e2fb6a016fc38437ebc61784172ab8376c51681b74f3d2e935d6747d1590de0c062eb3dce1748c0638d097928c8e176170c74c5f9660ecb29c745b10fd9e662b99551aaad5194af88ff8fb35bdcab356fe40c06653ac0f8bdc694f90d82b4d4102c90035377ffa1adbc3146ce96a8848ff596be635c5c1cfe06f84fbe6f56a0fd2f87fcf7b1531f59f11b693347ea60a8def8e158046da82506b9b2fe89770a4d6b13241e281dd1533cbdbc4700299cc28b4767617c6f54a8e177b21158b6f9b4d252228c04adf1f31d3cc4bd69196bcc70d5c98984652cb58b9b1aee75dfd7a64b79a0acd8074be5ea3f7fb2f1798aca02220a2f628cbaabb0eeb847e6211e2fbcc47f2347b7f5e9e44e537c7a9bde6653f1b0e3d55fb955f06fab57e290485558c0032e25ce5f2d8e48a63d54aec0af1b2d4adf7814cbbb766c86b004af37f2830045391d21ad8c94af3c5b0c85d6d7c05d2ac0dd0801660a2adb8778e3ef80e86ded3cae0cb9385b83fb4c3727efd35cd4552206b0c91383732a22f18dceada31fe4310540d5c6b113794657ddb8cddfce66e62bdf58651bf804d113cff043abc2741246befe2364d384403d3ab9dbb813f83915eccf94f2610c3ba74ecb2b691ea7117d341e21154319ebe446e294307cb51abffdfdf1637ea111c7d2450bfe0a7d21d500c670b10078a55c8f1dfee77746286b1013438355f7a09de4581c4fa39df78383d46befa571a0db98e06295d10d79ddc503b517b199a3310b16a75b859d30adbb8515f1877f3b227301bd1b935e5d2b53b449e79a3d567d31df14c28ae6e63d6e4ff2f7759992dec3fb5c97248420d015ff7c812990d9bb5357a7c8732cf263ed3f8c0100bc15240f7aa072b06e995bc9b5212b0e63e8ed9bb5ccd3cbee9283b628fcf1c243e577fbc2d103eb4263e8cb7336dfea4318bbe38eb1706cebc7837c4f565c885c75fd65513b079bea9a4a2cb0b3f6c5e47a4ae5a6af42f279b14a9e069451197569de5cb023e3de19cd5cab370fc4288abe804adfbd1f36cf09619265dddfe66c4e43ac9cdbf95b3f344f26e27a8376bd18a6c6f08a2b7596fedb6deb2ebecf2330ee40b55da99ae235df9caa98c047a5515ebe931e6ed0ab0e07126b37e730c0c75321e19cc87d226f958b4f002237b1967dff4a540a68f0046f126092a4bdb2d59fa619b437d8fa5aaa0aa5ccfe36d7b492bacd1e4fe030eb86a2cc108f351f1bcb125fcebf60c9fa4412118c45f36a35b460f89cb38c3cca6667b768a3101cc3a02f0ecde99ae1b29dec2e523e03f7ad7ccb12716faf49db07f019a44f8517cf55c96e5559c8c0c0657806021e8e4310bfdbfc3b8ff9297067830ca1d777bdac10f5e3c46c3339467550122a65f4f1c0ab8566c127634e3b884aba039e17058a25774b6b1c06471fc4c9b9dc8ffa06aa01dee5ad546b1caba1d5a1bcbce7c3627075131d8d9dee175f99def401a1286186;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h548d7d5406131f3714170b65ec833f7ac266243181746ddfa19d238e7284af76489961412b2168fcacbf52ae6dec337ae4f6676aa25d30b2fd23cd2394266f6b049a5a64a449406ef749c31b08c16fbe5aa4fed3e0744bf76cf0bb077552744cfd6cc243561ad39d5ebf7d2f338511589cc0113d4fda7f6a56d59556bff4ee400bfbd3c7000444e7a46fe2b8c5d7941e5467d874608161d2302fe2afaf3e23218ca8f9d251ac75469dfdeddc8628a8d00ac93523aa80cca840651e4a6fed31c156c3148e4d1cc0ceb1ac2b62637139e136e523ef49dccdc01cb1dd4a75f745222ad91eac692e4cf483bcacb867c890bba43806b775b526c3123d7c3fa60773d5f0a4f7f92484e43e4c76f7e86bc3369b7eb32c8296150121449cf1c054c99362de41cd4aaf0f0863bd11ea1799ab111e15e4d7f697569489acb84855b4696884b63f3eae5d673fa52e164328bca1044d18fabc8b2e72c841f1ad7dff50eb80f0e9bbb2d13c72aaacb7db34f84be291d17799c9a03cf19e3a3e58b6e307bb4925566bff6df9e4e58a036fbd695da09c81774741595b468abea71cdfd41c1737917bb60f4f00fef10cd8d54a59c5c5f884fc21757290095bb1dc4f8b7d5a4c879da17eb793bbd5dc6be7666e4e427a295ac7b1188d5327e60e2f02ecca7bdb71ef60c44974f7edc50596028b441ff46095bf9e56744ea414a83923cd332802d9d6cb10bbab04c453c15362613fae35421d1f28d18713effd8521212ec7523c96c238c8e9b19efefcbaa359549efa8ce5d20cdbd2ec32bc91655e33c7733631c3c9eec6876d2fee875ceadcdbe3bfebca3651be7d96be1871243053f22f26cd44289e323795278d31df8575a34e8002b18d0443e234e08a5221f9649272c6d8129758fb551d4295e48a7149aa769af30f0c84743cfc59189deac8d53bd1ec2a1e7758a5ab719f07ec9dc459bc5c78276c1453f53ddd778fc2b021d5e033897c3cf3e1fe1803aad95f48b48b7d122bccdaacc167695424daa1f7b9ba266f60d28d95eda9541054ae39eeba981509f00169e6c4d0c7dc057a6dcb8330979b7b4cf46d4eacb0a92763c7c8444545ccf6f853ac44460a8b71299b1b2235ce7c29904e6e4891d7749f8a13e09621eebad320c54e2e7984ae48e0da0ed7f3faafabc4e2740def8c53c56f75f03fc1616092fd101a1927ca6cae94b4363299920085f34b3bd9d7ea0eec7a75121ef00922cd8fab6cd9c5b12449e93911b3a1a7213270cbc6292ec60e5a71ae8e88dc7dccad5168ecf8e3d0dc43e74421c414bb09a2c539938ee7eb04b2d39ed757f1daff21025c576c0ec23c106ec56c2c974649e127228613c4a22693675c55310529001bcb67c9f44deb6695380fb11a266a34cf6b6a4a1ea06ccb8bd112ebdeb39aef42e14c52e8a5a9d41290e703ee354dbc78334fc544019d05d5298a58eca4aedc80e3c688dd62f437af72ca6079b453aa8093ae3cc266760674212cf0265b325db8a59e209add6e5c3b2d410c0762e2f4352dd32e40f8a7798ff12dedd553f5d9fe9342ff198c6965fbf0d1be607fc51b3ab78b45c7de36f414685d26c71f2703d219fa17022a7834b14968986de123a61556ddc9ebc1bd3f39ff00743e8af2119a2e53ddb1d65496d4e075aade7cd8b89ab6ff128fcacc28255cdf96f6eb810f321d3230e310e795754d7a02f2fd7034007e06f1c5321a13a6129b046dea12bcb9ec0e7e0aeb47667e3bd5e93201a068f080c4ede897779fc31b5f02095dea6cab3ac62da0f7530d25571fd20f3becf7ec8c2583fad948b235da1fecdd132307b0bc453f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hfcfa3af92e0bad00068cc897f66f7d8e25abd78bb91d717d81e66fe9471cf191268f29b1bc4dffe847db095f57b024eaacb0e45c6a6b2d5eb5e2a347f279f9ac7495a4c013048184ce95ffd2226a631aa919c2ee1deb476435c8ee96a04473bf357c71f20c9d44694267f1b543e08878aab80ca532aefa6b003d2b990c059a1918b6530d768bbac3f2a90b6b29ccb96c152c7ffecc1fe869927060ab6450efb4491aa1c37fd005b5f9bde0fcbfe351fd9500ade99d2a9261fdb6c7a6b27cef0aca69a2d5ba5b81a92979e9c77dedc21d6f209e3c8276d451d8737157eec7fe89b4680b7d237c2715d228a040ebd2da9cd830feaa642c91d64338de25ebd9b18315541cd8320c71865c088d2815dc731483a80a5184494c51c004da0302828c15af8909073c874deb510b74cf41a6cbcad17d9b142ba582b6497837675b286434ccab812248f3358f7d1e0442caa5783619592e39d6481f8de533686ebde603aeabc5928bc2314c1657b0b1af34fe9bb8559997af2a6827f29ef80d8d149f1f6726840cde495ba11067d91403faa196ba6d18d2cdc2ee49d20d0640ba27fc253b25b632d9884c322eaa413ca6b22451200cefb02e5d11d0f09e2215c8bfbe984fbd78ce07e7dbafbefb7fc077398995bd77eadc8a1ce57e7782b9c0a338e0dd1819e809af9095736fa562de8783d46b04954d2484f9c5f0b78c88641d73ef50733df24fe6c0939ef48466fdd799c93fe2e0fa97c673c778493a09e8b501d6ec31cfa5b00b4a731b4b78795c8399ebaac248d9ee2766a4f693be05a5c067b65abad836984f596b173536979b8c6f69ba63ae8e921335fb4d8caf34fef66bb78a675e9585a62821941b858c2e47b56872b7e7ed43795d493a94ffe8630ee25ebe55f3a7e20be8211e593168ad74ce3b414da3b47bc4f405df48264b066e80e26cf2fbbd038e1e525e7b0cafd150c8e6b2ca7559f60e04f384cd90c5949002c89c6e41fc60e75322b1ac2170bd59d843fa7fb5688abe09ebfa87a9b9a3069a9c435b386269f2638046688da0df9ae52f38aa272c169c83e84ebc4b7a20d81f4c9b3e63997177d52a6f2c051b319652c5604928f1f1bb4d451f180867e32a3ecd1b714b658fe9b041db441bd7770fc21fe370ab6c65b7fa0c1578092af6c7b2e7603491a68c6bc58fb82da9b562c930f68d7a72393d44ee8ae065c8d2b9a59017b02e7e689b6bdd6f394f933ff089123b022f9beb4b714917578f8e25e871cf65d6deb902c0172359d7c105081813ce08e55f55fdf42f4e22c15429cd8d8e0baf7a8f75d378b9c1a01f97f01a7059851ea17f7ba2ff513f03c087f146d1a4e7a218ec6aaf9500e0477c73b05f2fc785ca950379dc20ca747820f109bf3625502a677ebd9f48297a2292273d557936ebba29eb924ac61d756b2e162ab2505d1b14b986df8f79d469a33967a6bd39f96261495e0bbd13dad8fd7762785f9fe6d5a40859a66946dd6c22c6d4ec657140e236f8762d134fe33fbb5a7ee7ffb74745e5a4b7b74e737ce63d8a00e0e457a9c04ddd4b3c3b3b37537991dc26be672f2ae5ba73512bd55db69e53e42cf9ac5714d7ee324f305810888e50b0e27763eed75c646ee1f63b7cc3ec3ebb83314bf6b58f052b3b6977290a6434fa5407525ac4bd22db758435304912c5192f017a60431f73149d642a684c153068777ef2f515b368243a3c1dd0e3a5e1727946ee76c9f29bc3774f4ab1b8681bd6d859a704237e010305a5933b44f1925cb080da482f0d2e5a87b1cc208517e09034bc1cfa4b90509a088fb18906463aaf8b84c8e5ef8125ba;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h475ef5f6bfcfbf21f90fb77a07ab5cdcd8ddfe682c34c927ee8022a35b8543c7ec0d708acfce4891d0bb10cf6200c589f7ff86915c92af40af94f7453c9b089d8b233d9bca5bde6baad711670a65d21e0a4f338b0679a48fe9f271d4d8b9e6e10dd961d145d49c229221d9410d7c7aa98e1222fffae9532076c0d4ff213b359880a83963ee068ed4bc96c22c93e3bfcceccafe1d01e5294df44dbe842ea960becdc8fac6dc4713f8a0a05a7d20b811b38487fed41a7bb6ffce440c1751108e42aad1cc3fd513f76d38ddc26ef716e80acb1fca78ee6f6b42bc4a35ae85d7ac7bfff1ac452b471e3e8b24576c2296118b57daca0042c6a1a707d70f9304126563cdda73d91a70ad61533bef184cb11f01ecf246b1b4e088f5f50deda42e99e10e64c311dc906dcd5bf6d682bdf71db7c508aed7992118d13129c67539adfd5f4995a4adeddd72dd5857c26ded2b664de361dde034dc7462728629a2fd93ed0bfab777e0782d3b34d1abb62d41bf3e27f34a9b8ccb25fc880ca3795bc9a666e16048c492c15d3e1e3ff589bed000f5ab69f53fa3b2400cff48ff0e1fae3a89c0cfec2fc9a67beffb83de0231a61762f882fb58d8475700a8ae84f92dd0436998c22bfb975501155345919d42232b17acdbd25c7f8335935b11e67e0de7085c028b55ccefbc4017dced79213e1bf5430e2f80cb9c00a0abcd352efd6e5252e06d157e070f1ce2eeac681bd8aa9a87ee1903e602303e880fed4034d7f1e47829998eb5c4f1de23e0baf58d107fcb0a5e88b3b1677d960ad29fc49bd7d1a672c97730d74ea8710d29d7a86db546d4771a3b7b74cdfc94ba960b177a1e99f8f20118d9065832043524335791ac08ab656da2dc4edf1e5338e7c044a209ad88afdf578b40261aa7d91808bf8b0d2c384021a30721b85d6f9dc8d1c307ed028d4e6433508d04f16c4d37a7ae9ebd08be6333eb7fba64a9cb25b4a22716bfed4f3e285a73aad7a89d9ea6b1a9dc95c2bd188772e9ec9272278459f682f795a7d4d3bc16f8580e2d099532755c8207ee4d12a4e5ca27a7f65ae837e51b8bcef966e445d8ce7bb65f61fc8cda82a24d8c178cf21b4743f7626c4fdea965c10c5c1eb6868f38199155ce24d4ee98f1930534a6414dbe42e6fc5614d4da95ce155da50732e2670591c3d8a9f8045db625d8e6fec4a17562da54f24e17c8ef370f27dc348dd1cf79f7f9a2b9bd5818e3ebd06256ad9f770d1dfffcdad9e0623f8d598abf3d6c5c01d28dafc9ef03efdce404f0e9e4ab79771d5b07ff38e9cad7e8a259fc10559bbf2670b299caeaee815de536e73a8911597139f9aa9256189998155977c1ed9b8b10fbacde076fd2e1981f92d7aa4e0b1fad132b355e002960e26407d470781d0ea13f8de7ccf983ae7d491e3e4bc0757e6fafdc01156a102777f641fd5818a535079c088c726f1982eb3f1597e70ae422c42b658e65ab3bc9683de71427e1d260a2b508f5dce7e37b509b31dc4c1445a8deb148017f095a106e4d7d9eab1ef4e55e52cd5e44a89e0d9e45355f6e81963bfec42467034487b69bcf7ff70037589f721bdae4379ab8654472d3ddb13afc9326c06d52973cc55b5d6d6936b0ace34bba6858e94c087a3c2c8e3f6eb93a7fd30590e7f91396c250b50082b69fb803b4ffb6325fe08c14888451d4fb39d13e93fb7452606a56d1cb584133d5eb8fdef22f85397d4bd7299ce7b9bc821ee365dc830e413a820d6821036589e986700e52a7ee6a4ee72db37cbe7dfde6f9707cba6abbf91bf26ce352bf5115ab96eb4af7052c6e6ad76a53c34334fd573d8617;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h64b05331b4d661733fe80bb248070c72f92a5bb5cfb0c5a4dad093ccf5d5cefcac4eaa76a116474dd9cccce44842a00e20c29f5fe71795dc9da9a12af82b37658a53952d3633a98b4abb3c18555f799878c6c592af8e037bf52d8222fd230533dbdc0b746de72634935c0e66246296e88881779f335a71cbb5cedcea4a7c8a8486acff63598693c504718eb867c03746c980e2cbc41554919b4438e0607a4a11670d1a6c364ca3eb4acb4a2151f4e9e41ad3260d3541d1d33987bf1d14477c97a5157464a779083943eeba39d21ccdbc4f1cddde442396d260fababda3623762639e9db1a0a65d9919705655a36d046d11f731908c692ecdb3b35b42ed772d1af1565ec71058acf9542271fac3fc82b999ee4ce74a2302ebce473a68fe7721c5eeeadbfc75fe5d831128b36cbfd882866db2d78d4f653a9c9f713f9067d692aa8ed0c0b73bee283f286064a60babb09f97c41616daa35d722ddd8c64501e2e8db3bd77468ad3eb39417640eefe0177514ec85c04e35a529447b0e8bbc3493bb0d65bd7544eaf1d86180ee3f76e411c01e42d9dd9e0b1385fcc7641897c4ab1501060bc0aafdc9615d6495d36dde9737fe82fced403bc60949bfde1de836d8a9e355e3e6ffc1e10c603d97b379284166ab79e92c53f9fd2f5647db10cce251edcab8daa32c61b0304de88f8d00a278f4c717a5372cee380c0c523e54b3a8ac21e4209edcd2805d31340af655b4b02f13edff8c5ef54bae3dc134bb101222173cac5f50fb9a16d6c68a22387f417505f0d9a708693f785b142f211de4e20ba3a37d43bc4d80f33418d8103d5d85c31b93daf318cbf2f861327c68e9c3a51b78f481e4a2af76ece012ee6f80544036e810f42c4fe181378e89693fb97e32de91765af211b6b0078a47ecc8de5adef6d680ce1e8f716e01579de7010cdda83effdfdb07c0543a5486cceefbe3791c576fb92c2c8f0de4331960c5ade296e4b985c93cbed4606eb567b1d1a3a146165729a99a879f7bff9bd9688c28a8d371ba76fe606ff250a18bcfd611c16b5cd9fb10bd9167b24e126c232cae1882d58809faafcc77970eb329dcb810fb100d40f88cbcf1cf2c1ad00ef18f8d8a0ce6513ed8dff9272d28d2d0bed8b1854b37a1f1455963f1f3d8dba3f2a2b84dfbb92bd21d7e57718bf853ba3f51e07b7590924e0ca5f046d51917e0bc7863a4782fb4e37c7932b154872bf8d166298c677de2a65ac494ea37e5d8a4c725baacb98035c5039b9b7a6d4814863477a5e8b3272d6b871c08546cef410101acb9b7cd4f0230dfaae4ef83bf0302758ab3d652537b3faafbcf0cf0c3974f2794e24dc76d100ca4f0d0afce0765b6266e1687d7525c9a733fe897d87f8e61c1db5d454eea547b2485ec4ce9d5c11fadfd0042de576015280c54e3baf12ea55be038a65e739dcb29e7ae86befdb7953d99f11e298c5c6c686ec8d94ca809ce24b8fc86b2c618cb596b7bce8c09e986636ecac6efd23b278bf4a618cf04b63628f56b9bb289e6961d1dfbe43cf339173a9ead173441fda1ddd6e9fbd9e95a2eb7bdff61ea966a916027ed1bec8582cbc3d9e7728ab449c1ba554493aa7d0be1a94e4cb2b6298fdd6f03bab8831f109edf54f3ef312ac09a3b96071a4e5c484fe600eec8855f74ff2261d74e9d47ad2aba194e83c43a4f1673c6f4630fa7a04542ff94d7f98e32e0cdb7f60b2364cca2311e33111a3cd19cc8c159be3f52bdf60de612dc0e9d07419681f760005c867c20ebdb8a3d39091acb780d3f363c22b2184c1338ab8ed23f74ff52d00e96963f34efd4b83660413b530c0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h51578fbd5572f667f192eb9d2fd92a7305710654fe627bddd5758c27d9376656953b20dbabfcca82e5410944a8649f5b0ff6ce3a4f2112cf3900b9ec6e467805b59d1cb12cfae20bcae3d123e15e7d691b3a545ca6292d1aaf554f98149aac48a20558d8f4aefcd65b167f478d93531022a3dd1c7b236db7efbc202bee6c0d05d0d46418d95d0cb596afc8ef22eaa057eb071106c77d2e793ec65ce8a50b40a8b530ae2256833daa30b29d2859cd4306b97d600bd828acaba99e32188be3cbc65b042642ff2aa86ec9f7ad812a9102673c9fcf9b120d4a9c2f66658e8ecc5a96010a9af1dd85c653797c5ea3d1b8f58c409f3ec4286de32c22b2f5935ffb5cdc3294709336e0610f7fc3ddde8827c255becc285bc653a73ded5c2a0809f3b8acfb366f5209864c59ed7b5b05a4ba63a7c8c098aa6bb40b56b7970c46530dcb16d81523ecfdf8e813e82ff50e580e6b3c79e0e999d7b502fc5989008490536e4f52a5b359878a15094c1f2314a7510bf22573e1bf8f70e4621f7e50be0ae0838661868fa2951a3c895e84a5860b190072ae56b3bf605845c6f5b26559adb1494e560e5d65a42c6c34798877f891b55e49115ea086dc91e080942174e4e0d56167b9f6e4e7d68f498dc1e61eec9ef5f6c130e39a7fef1bb9450d66d6f4eb2a23487d942b6c5b1d040e642003e86743afbe4c4f8ef275b2088cc0b8f0d4dabfb81852dc4cd5b1cb1a17fc65f8cd497f779bb30a85e19b60644b96ea6f884153224d908a5d65815731173d467d60c1e1ce7a31d019b2db3900df72c776f0d87f43fcbb345716d85f0c2bf5338828eace4bd07ae04ddcf3e31731cef94ce2c4df742f18006bbce2d5a0b2006d7a02fb214616e26bdc2ac1700057a3c5804275bd97c96033d5cfb03407a82677bdfb8c052bda7c49038a0c522dd2cfe05142342b664fee5e2b205dbb452c1a216e7c35dad5e5ce17a19b6ec5688bc91383fe6b1cd3ed2250b66b3b1fc89390d89875059f2f501dc78d911bdd94e0d3d637ef4b2d4d65367b00f2b13319e7cc7ef1f69198ad96ac87818226405379731b19934375733cc3226952510c5ddceb3c0d7597e2e4ba0aa076080bce780b60b887a25aa0ed9f6d34c7478f4c355ff953ebd64f7faf58cd9c795ec2415c50a1085b42922db0500519d28bf07b1d358b1935aca9c17b07b7c62946053ac50fef53c70c93dd42063aaa1a6bf0655580ff7f5c124a81c5f587c097e34423871a3753a0d4b20aade1e897c6c4b479cd874c12ee44f4a4079dc29b8b4ff7c5e2739057feafface442c1ffec38d1c31640f2161647fcb2e75937b79a2106afb42ca3bca832c4316845274be17ad76956364223e11fd874282da1e64ff993e50df59f4fc9f45f199c07aa9d51828586afe4ae7e31bd679f2381ecbf2951e0272a618b996bf083fc684129073cbdab4ef64c4fbf3ac4c67a123ec032696df4188058565172913345d92fa98eeecb3a0c3b057ff0e95d32f995d77e7c74555e7a5421dba9dd23fc99546dd46a39f72ff85c2d1329c1bf230986cbd05bb609ec59cc9bf26e68b5decbd9b44b175c3251a2a5569bb5ca0af2341f20fb8492ab5bd30c12f4a37c76c39fe84212b68de1fa13a46481caa7e77b8f95e49c2ee86d17a1e4aaf0e7add338bef2f3ca45ddab992df22e8e8d92b844b0beed4846cfa5805d9e4b7f2e4fe9204d03a2cf2a37050c422fd98738c4b0c3928527de59ff4323064c9ad01d355b43d691f1fb1c55984da3fac5693d1c5bbf63670dd0a381504a8d0784a6c705db15e8a2028b380784bf7ea07182735b71579a3a91f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h644e94676d9d1155a1e7a6e2d53023263f3d8d2c1ebd6a0af0485065d9092d121183d3bd8e8bd23384f1d9a6a4fe2b50f32658fda443c278cffeaa5a40dc8a06a4293eca975a3e9aaa38419f096457a3d004de643fddc6c37f117818fa9bbdb434a78fbf96a80bf90a0f8f6bf439e247abf813c4f55a996618b76fa54263a75bf5eb785c67c821f9bf91c745ca55d39785ece0bcf96bdf9b29ea7bc35ff3aa2ac877267efce890b2fa74e064cd13268414d21ede8bfb370670f3a620aedef0007c6d53bdc9d5f8dc5374812020f14d9c59a8459ca229d543fa2f0d44a66f178a8abcf66a697c571f533963a4b50df66a1dc35bf93f214a9d8101ca87e2236a833b548e52f31e3d1f0e0278507a669ec4d4adadb2044b1c5077bab664528d25ffb9d0fba1d0c41a1f2f5937ba599fe2735b2c3305c74e2289e2c2ee06eae492e5a3193812044985a8fc4b77ff2905cc74a18d85b5269b2d4289ca96b8bb7f1ac629a4d992e2843fa14914b57b7063f70fe31a03bc02c23ad8f5e6d6933e9ea1b832693d1b0a27a06af3e23c3c5e69404b95c8eff50d2c30dd2db306dc7db6f051784397c18c8cee1ee3b0d85f04fcf003fb0f2cb51aa47c7d3401f1f49f3db3b232b77a6c8dd4e7a804680d092c81d2c83f1949dba8869ecf119b3395c8bda9ad9d2266a4062da18e7ee3b2d08d4b234e39d2c9a0d88e9ce48930e53966fe59606d27693dd1fa1eaafd1b28cac803506b1d84191dae7acb6887f2897975bfed6653cb9e1f89ddc04d582aa44f4e37bb528280234dad13939122574f64d7926d1dfa3059b35f34db73de09e4eb37e04e744c95e051803cc6bcbb90acb38e230301812c1ee9002a66a71ac8d75f48e26c6de7970459847306467a4ce94689b59612b6bc42204e0d03c16a415ecee8b62db1e83176fb0706be6a2d523590961ac2e83e4b05150b2cacb79e609e02bfc139ea4cf5374f33200dc42be65b3ba2cf43383eaf13eb735b04c6907595267dd972a01cefc030d19bbeed91c2e67ba9cd627656076543261bff13a891f352487ab664269ca6cd7bc9235a932fe54a93b7dde50108a30e253a4056048a39e278234669790debaa899eee259136c8c0f692cc0b76a563b567783050e8cd68afef780c963483345e07416b43f5f15c463fbf7edbc62b789c008097b109e61da460c22e4d8254f76efcf1526db62c009617f36a0028c99ea27eaa40355a8a264f5aacc9b8c81f82f481975b975fa8c75d97c88253082d5e5020cccbe26909c7a234566438ed701fac75245bfadb535757c427fa3f64db2d1f01b7f666bc96763d823c8565c350c29e0e9968d6c9c93fc7c96f8c8f66ee4bb15eb6bcfbc8d2a460cca8a58dac4897bf20c3dd2d68c6ae3d0f9a16dc57f772c563a15da17c0b6ca836236472b61b70e7da4f7dec106edb1c794010c94f397093766ac7eb9d03ffbc810b0e408513c2ba45fc9513e5cbe182526a77900bda9bbcaab1d2d3f66bb23b3042ea3f381c72afaab209229d29705fbdad120bf159937589a73fd26267e63f761c616d50717941af331fcc257512fc265f60ce21a1ecb97d17ca3b855af85807095b803398a8631be6cc17fb51ba993806ac13e49d07e9c501341587bb1370cce4b13d563de2463bf67dea79895628dcade48e36d0b87fe256a993ecdf433e7022275ceea29038e1060c27bb1f1c0396661c2d5af4b54f72aada419844cd01004372e0406b1068f193c29d3527dc5724ed277c2d2b27eaa894f07dedb2198a42ff106f68231a16a47e34c2972cdb152f7d7d12d6a0d4707fee69fbd1595f4ee1376c74;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hcfffebeadd8597488eadfa4983b2e2a0ed13afc5567c4aa0d50591b1b41c02f2445c7a034b42ddb860952a3ffceddfd863ecd7f33a47bde38105d9cda99e9b4c04762a39b1c6bbfc77adee0792f7c7c45379c74be47d0bae5ee3701442b62d7ecad696ed3ff7ac40d754b8863854634eae7e41659e2ebdea6b9dbec75d0b568f4721b918ff52ffbf0b1206468b02de1153addc90c58af6df0472df3c75256f665ad7a902c28114ccf001fba09f0fffdf3565bcc6757a80b75caf5e021325ee4e4a1bd5f9ee5569e0fb4fc6a5b7d06d2206789ddadd03d348337c055fee6504f915b5b1e4c2fc6c148e5c5c7a0cbbe459effc38640af1e2e5310735d44bd236647f02f5cf8068658c03fa10abd90c7495c55dfec2be330a79e539c557727593be1b7e4ce50ebe071d0aba275a975130a6ea34be34e1ca7693d5e87dd4acc7478c214db6b185e09836f5b0d0b6ac7780994f959477994d59c1617b082aa3ebb63d4d5eaeb104e5c1412c5970fa69acc9b14e90c531b6b8e2d390c800ab5067e495d49570feb4483b725fbea6bab4fb4a034a2d624566498b15554d67fd8a1ceba677fe3595bd2aec0b2c85b31f5ea1348dd124de2566429d3d62ee2fd0d23c291e73afafcfccfeceb498517570718b7d9f3a1d67235e282bf02372af63feb61a2889e44bfa1aa4d64bba25744999a3131ac6f6343b289570f606d6419cf793dd416d2afd636f3dad56bd6bd3edc02c15f3215d7ae09eff96f0abb28a700edf7117d93c106d425da9fe904bc8588d42185c3477b13a274f0e198f0258dd0d73ec4755be6ef2a26b05f2380a2ee5c3901540e6da356f4fd36324c57f7557ea8c51da46d985c037e0ba5d0bbbc9f9ce404a619d45f249f03a71cd8eddbcdc4b5e6bd3a0523213ea88413086691c51ce987f1d4ff66545ef41aed53f2768d136d26b95aaa5eb2295f344091888e48fd6bfa6e51ef9abcc83a7574f498377df6cb0ad8dbf913cf66b8f58115f7534cc6466c67d65cd69149caaad1a987a0227cd2ac9f6f622b18762dbf436c7290ee201d0641c51b23a89cc2ecee604e17fa64047557ccca32b68800a93c01ffff29c427262ad05efb81e1656db3e58fbb430eecac4ab0a1a2f621c7c8937022070055fe3987ae78a2f7b237d424b3317a46824425bfd6a9a0a997a851a98b44a9d84ee6220f32511d7426cb16eb908c37cd5da908a929a812467233ab1eff53740580352e89c4d8d0a4d3a3eac87e04c1aaf6b69770463e60bb966b177b53b106ceb8e8db2bb7a8c2369866ac9b036f8cc419bbacf444d67e8f5592b9fc3009954662648530e99c76c6124fb72d47825c89f4d827167c4fdf1e7ce2274541e7d1ad1dec9e12c9d0504a44079667d2f67b30edba0af9299656b876828ac030e46d00b8a64774de377c875e3c6bd4d47f21c1a2d237cefcd7b9e83a8cf8ad8102453093091b796a68e69f54dd24e72313a37154476941895b8aa901dbf06270a0d478fa381a35d5d8fd49078878d4b882bc234f2204184d540c8fd704aef6de6c30bb7f7ac899539f6df6e2b7e2ad7cc412ae316b2a4569c6a97532328a4702726643a2576ace28919020f371f4ce5a0d0ce157bbf6dcc8d8ab1d0a4f95d9d342538f34050c901b78f3599f595e1456cf541dc58419849c0c31c47e4da12d522d435bcdeffeddc53ae21a6a3b4b40661bb159d19af754990390d58a75520934a9a660cfd04036c6e0b756e664274d187a31ebc1a2335033bd66c19df78ea922dd1cf4b4990e3902b53d9f3227e9e62502e2103889fcf29b437dfaec666f02e633193b488a371ae;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'ha3085a9181397c4f91b633742f796478e9429019846bc11eb028639c149f03bc3e32453b1396d07153b8fb3affb7361d3e67f5c4de12823d343899ad53f04f70639e1418e76d76c98c3c87ce1ac78256fa87d04c2671eea316cefac0f7d39f09cb99535b447927e2715027129efa61838ca11c43220e7bfc43485f2bcaff8c5b9a8fc5bee331d53926c7f42e65732e76dedfa2d69543733d7bbf8ba39614e437e8500a19aad718e85a23bab07e57dfdd68a6663f5455aeacc63b5f1de3b121912faeca568f0814d912bd5adee92bb3d2322f73a2589081df5957a807a51ef65914437366eadc556a7cb8f45080d1724340d45d62eee4e201277e2ccb73e1449ec9b7e8630f1e968e2c74889eebcc6bb0ef8b11906ce86f068e62e8ab50558a34cf742111ef5484026f34b7ce4f2c593de425882e972ed591f08a618f9c82a38863d8810abdc2e0febf0a77afcd1ffe8b31d85c413ea81bc417a5cf6d113dfd051b0d13a678717040fdabe228a63531228a9c8aae72d52baa54ee6c672d66a5cedbe159ac02428bb0c0bc259447ef5b31f984f914461d54fd1a616d133704e4d032f1202893b84dc0620132baba6489d2a1edf4bc9e7b7a4bdcdce32c1ed617ac786699aea8abf1e4c355a5bd8b40806023e7b8959e18dae0fe30a91b0fa9a52f4b08705a7510f8ab9c66f18e707cb26b8187648389147e7c05e941614391ee0668e1171a3a6ca58e3ad249b328f55afe3a7301c0728e9ceb0771297035c85e74090fd409282abb5f23e39578586299541661605fb6f202204b2f37a0016cceb526aaf63d2b0c277d1a1f6cb931f2d2b64df7cf003a03c0e2abc7e6f27b6fec39f367a4b3284ffec004a05547e3f2c06d5d819dae3d10d7bca6aa768db5a30a46b4ff595185a850f823e2effa610681e1f3f7047c4b37ed308f1ef8b4c0524d571ca8e750207dadcd80968f6a747492b9e46f5730f9e26fb780e5e44634b5e7765aaa219d01e5cd663ff4211b5b0c985c381cd9cb2095475e54fc4d8ed131b800ee193996d34751f5b566a2090a5761a3c617d2c8694eab6f70e1712a7140bddfd41ed3c23be2055fea6155742c8699c2639036c6e90ab07bbe16058f6fe0d28f6ddc285fa40fb8431d63da37d060bc3042a6209f6cef8c432030f4424ad5155d627e3f385b3d4a9b5bddf5d85a82b68385c98c1c24230c87b75bdf869293c2a28e3ba7ac94b1a029411a1008bd01ff04a2b1c7a90e541a872765982fb603f5e7e274db5ccc0c71e9bbbaf9d077efc4255a3b4a376267b12f997eca055ce6b200336c1dcea3e4730d3b7edd672a0087ab2407eac3641e78a59783bfb9e6a6dc17ace34784fb72a209947f4135341bce26df37a86c3d742bcfb9ea29eafe108bed27528ca585052fa3dfa26d47a8b00764d8561de315c6ea705672481b42be7314313bbcbca49075680c29645f877de81922cd3bf4dbdac788c427b88db70e042a31e257917511b0ffb21ad22e1ccb9a8b6fa32c27d0ec2c122ae4e458df801750bc4fc5623ced37d51d985269527f7cb8ad3a0ff24f14c8bd5e3aaf94382552c9e40d100c9f61066e48a49d2acaddcf904b25a9d001d6b563e062543555fdb1a4c4a9c1cb51b3543030d9b03af90d91a458c022acd8cdcb92962fc6398572e9a34ec414b12cccefa908593c0b273dedff8f824439cc8cbf3bdbee269797dd79c4aa0e182e56d282c9e6ac3c31a849c80374341aa4883414610558b7b8ef741d4a6464ee423e0940d20d6e5415400f07c543354f7b61ed99b500418c75713815e2547a6be9f36830e8aaa1997ae40e8876;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hd26bc94809ce4e8fcb5e192876481077eedc258741c13992f132279778352afb09e6a33c8b1e59ba9f7a09c34d19cb1ebfe2fe70c499425a4624a72f1c8fcbdb81efa203c1c3439d7f66442c3d6eaefba1e81b73b473d72a0b53179046b0079143bbd5fcde52fc4c43f1a1752d2b440851979bf99c2060584a1f0f594b327ae9f8a96023d4983f4d9503add17f424441a967f683e0af68410ad5319f637d2ea4f9f8d83e5d674060997e626f48938f371aeeefec5935a31ec91b06087277c4e577a469c2876b3dced121e91f650cc51ec6f6dd0b6fb939b7e9b11505774e659be3d147f7b6fe7efd4e98274af96ae438b4c62c90d021fe42cec88e6d512ccd7af029519232fa83d7416b8646f12785f0374544860e8b822946be08497bc4eadd90aade1af47422bf2e1f76f4c9414ab8f32315c08169ffd30bbfd009f1d2639032eccf40df4e2660886662fd4d492bc70b467222fad73ce55f56d8461b4e9c3b18ef0852243861352b0d29fedc97379a896d6c3b1ab1f08412d2cb80fea013be799b6541ddf4e0de8f1a3c580e7ee54154c011128d896e6b2f77f7d6cb45508df9a1004ccb5843978de53ed5f4ec0b9901d4e1a6200ca3bc167d11ecba32e10d2fd40b9a94eb1b5eda750761b5151ab0e3466f82bfb68a85873b2c5feabbb3ffb812ca8eb39d7b55b4c44420e3cd6b506250a2d731e409b2dcbd05efb0942b2ea2f7bc800a35716f1458b826ab3f151a4f43d10858bf8ba67135be0e5bd900ee2a1983b66f1550595a828e8fa5554e9ba3f0777c3eb8b71c90809a8fe1439cb8cf67f4b6de8de719cff6e753ea895921a103101e8229a896a5e86555b7dc928f5db8e78ed8f9319745a491d64829f8d6fff076c2c27fb362208b908b98b0955c26c173c0638746b8a13808851ca378f0be2cea0b790b7835ac2bc200ff4d031ddf6985523f0e66145e92aa6596becdc6c7f716135255c20157380bb3b0bd04d3e7ae75c13e596c0d9f631b83155f09bed24d84ab074579f87430fefdb8abef2527aa2863f2059e5cf7318328b0b3f69d28a689a3ddd8e7e12823bdd9b3b250b7bacc5e9872d57dc51e57cb399af0a95a3b586cf6ae04943193c115d276c96529fa622bee9624bbfd44b8459ef8846f56ce4bc965ceb0aaca1755d68e9b1fe5e135c447c4e5bf437e643a15c76578362c305cc46f99b90e62e84af476d6adbadac1fcd1912027fbc9ccb06f1619a1bfc0739f526b9cbf51cc4689d946c1a6f408b62aa3111b0eb712eb295adc84198fed004436c95c9860c467f64bdec571d72914dde5c2c815edcbedadf51f7f2106140e9d1957d2e25d39ca0188d527e7e1b942e77a4c2f66eb702464b75e6a72113f9aadade9cc4758cec8119cbd260b6a2ef5ecace26fd487c711e0b069e40043331ea4fa25356d30a6f8d63b7508fc29a4f1a893690e1feffce3f81206d998ecd443adfe3c3fbbbfa338dd088ac4fc8ddb2d1d75853c0bb3ad63cc7cfdf1abf3e2d820482acdb56fa203ec3286646080d10852d5410a4819743687622ad27e654796871abede107daf8a93271cb6ec26e3910fc42326b0c32f57e29aee168929c20f58ab5099a8613a0e3ec19e55407bc63b6bf46d902b3c101c54b12682236a7325937c620c77440842b7bd7c28ac8597fc0b0bd1d67e7aac5a7b4e99c2e2d34bb3321f6e9260060bdd605655975aec95d4e19d3b0b07dce3980d84a942afe0835b927dc53618f90a2b7fcd6f0ed259a59199315dfd0dbf6d50e42cf8f6d2aa8b6e621f9221b7b06647668d8bd363c067c4ef839998342f2c1766e6c6267757c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h82a0a56da08000cbef6ef91b6bd7fe6a3170ac9fa058d033bfb84cec65d03625678de804b6249a6e2813dc320bed4aa7cf13a7d0481206e73237d6cb0a30c1e12b17f8ce7d5032211200fcffbfc1e835e5d192335050c2c15da03c8f967300d5405c8680b39a6c1868867012b7c4473f88c4306058721806bee0a0b0a86751f8e7eb0bd5bf012c706e9cb885d68a25e47d5ed526d13d4401311bc259d033c00cd07cf945e1253be6b0e598ac1670b9d9c95a5e4220ff3ea3cdb6a640076cc5c513eed050496774f8d42bcf10fa6750cb11e53ef9e260a4d4314663d4c7d0b7dbc1ab5e3759cd1a64f63eb8a364c9ecdd9a5f8f5653afccae7c5f52830f637099f115d442fe9bf2bb4f4fe1189ef6eabd170bf4c34e7897d341f0eacc3dc61d97cb2a6268316aa9b72537e7848794632b008dd8514039659f6256733ab1f431cf339e87492f774728e2af6041745ce3286ac765ea581d6d0d29886bf2c7e7a815812766357cee3bbc5cb4d3e18a5439bb21da1754d7533f63bd83e27f90a44995419a709d3f71b2483234ae5a430c5510d6de03e8d82e09c38ce3186a6b95700b8bac564cde33c4a35538f3b88e1beeb85ed036a11e32ab5a120b5c49fd54751ed7ec860f40472c940250243a8d7e94b7d713ae233f670ccf31e08c48d93f2359c742505e3284c857cc812e2c7029ed35eb1b7e705d9ccd0b9d187203436abc6e4f28213eab260b71a7c148c649a703d630ae97a34107c3bf7b6c5864c87148089d6c1d91f5b86ad721f345fc957edbf602ea90363f703bdafa32668fd26dfe226685c2f6b6ccefc9ba89b8fa87a077dd077c766061e16263fed896b014a867d304a71cd66e9e2fae8c00a16d07c5cbeda726e234e0f2e5261f160ae379efc4202793df41a486a8ebe0de381f041b5fb93ebefb8fe6b010befe467b370ef8cbded5653d1cd475eb184067c10f7d04f30616eac380681408ae14b6014c32f4e1f3f9bd9aafe9bd2047fa3805cd111b861fceda26a64f220332a09ea5b9ead9d0c353f0bca97bcba4dab7fe6615b071a5756f63df8739d5cd1df74588c0736485340594b9543749a921e729b07448633c6ecec5def28b6d1b02575ab9014ac8af4a04b2caed9f5d451f122783efd21c87fd6d7ae1c77c8da1657755a56790ce050f8567afd7d3e41fcafbf6be24e51eccb64f060546d1ff478abf142dcc14f08eef0f65cfcd15e445fbae33fcd8f8d3d96cb0936089c27529b41807c34e7ddfd4f72907ad023dd4c3442a240e53b508353ea8c5fca7d3ce81e3ef33a24ceba431d366d3712474f4de586b2db6a77d96e0fc732843eb3c0aafcf753bfb89c32a63ffaf0bedca5de9bc06fe7a57cdd1349c61dcdee878efa724c6660105c43c97fc29bd51ecc991867edc119fdbfd2669cef9d2935e32628e5e47fe4f8aba82db41409be01f34ff0fd524ed4bf682cc9223c4eeb834c929967f205f5021987b5b72bc0f4caead73ed8e2fe9df55b2e22d538aea5b8545adc73b0a6701331f848cc86143669613a9a3d6c84e52195bd93ae6bd4ba578ab2ace08d833c48acb7030a592d766ad50d8ba34d173f5ffa79ddf6450b6809c199608d426e30338963b379d96bb2df08a2116cc045f04dc6fa97c2a1247913be042bf6c17490ddc38b7b153dde1c4ab9483900cfc0e8c6d4f9a6cb6d3549ef121fac0ea333a6ee03db234f85fc41d033c95f0b23865ac6a358dc78bc40bc5f4ffb21c6caf9b74391abbcfe032fd971b01f705a24bf88a560a161d64a97802fb60257c20d3f3ccb9b85d0f30d37477e813a5fe916dfebca8509655c42b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h8306461e7c3a230c8b0b9ebf5b7602a2355f3b87340b126158486c83f6ec4747cd015559f9f5cf7ce388d228a79b71db329c08f46a25b661ec7bdd37a6db03c9290986a27c9761b7430f32ff747237f6680f65bea9438f8244153424a9f2f8f06896dc9f946842298e945c08f16b596a0271dc2983f937f207661428cd3af8264045a71a4ca09f0dc3e4e0daf457bdbfe23a7db8b28eb5e076aaf218815f9181ac53b359ca57cf5a80f9f779c462a46c932decf8dbd564cd1f5c39d42deabc4611f841408c237a651171128c2ab085bd43ac1b48d9a58ae409414d70c42ce5fcfac1862295371603cdcfbebd5a8914fff746b7aebe24002e4443e125a62f9e6d13448c467cc47315317bf00dfe6c54b05e06ef7045e8ea44da79cdda27385e7e7ee8802904a8524a99b2b2d3b94d6573b12be92ded74ba1e6d14ec368d96f746ffcb174cf9a52d4994a3b99438ebaf8932e69393405aecf886d455c92b807c6f5960344b1a70fa26cede59d62eb75d1d9da07ee61eedcfc459dbd485f8ab742261af7a1de91643825ed4c681180a0371d9bde6510085bb41a67a8ed374cff5459f4bee3652d9a4ce1d724e7b1be229a34f30c7b17ff7bf9a3a3cef0d5c35002a4cf2c404d525e7cc498682f8d5c09479af97a90a26f41187d9b1985546e6e89f38b455231526f6e17123e36f59c49f6a2e74d4963fe25bd0ff1db2296b05667cb1ba0d4cc51c65d198c82ec434ffad921fde813cad68b0f736dd92501f89a3a2b97b5fdb160d06090c4f655b3a83b68aed4add1d166768590e228f7000984b50280f80ed971b63b0c97aeacb248244b380d991a4c5ddb57240ef0fb94d5d1443a89da44772dc218aea005941015589243902968a54fe3def55c94f49e92793a902e6361f3068709229cab0a3936655feffb97d473edc7302164e08636201ceba39b195e3b777a2d651e9bfbb003c4df2de26fed1ca463c5a94004991b0d74acdc2a7d0176eb7d54ae25836a8d97aacf7556aa0920574d74ec5516694a01045cc7f0bb5361178816f7443f0731c652d865f1f863c49d4aefa2ed9b98bab27b7569f61ba94486d6c77a35c742290d72a0f2e2dbc5ee50ff472113bdbb8a70d86c36a4ae428f1fb281eabf754d90394cb4e054b2c7b8f4854b0c23aa2337b6efaf5fbc98c809d735c69f1ae4098621d37a145e3193917e285549b2cc175fb43196e70675c723674a52af8b5aeb011cfb521c73eadf385da6114bef8508d30f179dafed53a50cc59dececec221a1456379f113b3b5837eb5d053cad199038a349fc79ac2b273cc8529247caaaa3d0d8a0954b79105ff968ce0a72e8d7b8ad14d6e23ed50609c11316957ee0bbeb87741786d4fc894774dbe1be3336086bd6b99573e44e7966a2a4041ff61e3927dab8dfa66a30fd2af62293bc39911c7eb8bc0210941a16a11c9b76de466ba01e8ff975859116bcadb0fb77ed21fec05783810454bc1ba32c818c0d26ae6c3c6e59bebe1f8a1adba3e3221cc9ae944f37db778b120757e78d45ffed1f6230f3a215e9ee2ab20d2598fa37663472621c6229ebd4df6f8ed097acb8db9e2bfd548bf62c095c52e5aa372ae074e6356c1ac166390d1d12d1b33a9ccbc88beb735da8a798ef759b21f1ac872cabf0c142d6cde24118104f01ac72ae1678179d4f4b8b36f59f9898525ff7a68a083d8032a628ab0263fefebf5b5df991551d2edb5cc032f75ccb66422c2ad421d14fdabd834cb6380f8191ff195634efdf8fe1c8808cc198139b5ef0105577faf1566a5301d90f45f794b7406f7608c96b2bffb8773ecbabef997;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h95e9465debe2bd3ed2018af221a2d2b8aa9a16e99185a6b9db4f80e2612b93adf74df13296d1b4a949f5c8dd89ea1dace28142be09c7b93e225958846b1b65ae6aa9edc038aaba85acfc06423a325e04264bdc595b3a6ebaec654bd888dcd969977dede265bce404e448891fb002068b907f2246c46827cdb181bb771ea880ff72e47e166d71264060c85c2550f81b380594c2832ef52843f08e5d92ef3076e387215c72a63820543143db11cf8e6269b94afe25e32264732d71e9fe2133628e10038086a4b07d090759f5aab712aca596e7f0abdd9ac1a7c18785663aaeae1fab8c22280687724ee833bb1cef913588ad4a976a533dc1223a291f0da6743fc5cf06e58074d2e5b27085e66662096cf3aff47efb22093aa1ff840e1917ef67f0c6d0c4103a73bb850de37d102ca6dcabb2e53e04877128036e3015884a0c17540d68679315c359efb78f28d3a43ffe4770dde561e98c058b5aae63f87a6b37f68db05d394fa7714d55b2b1511c6aa15b1fb3dab6a7f49b07e09aa74174a329ee0d20487823c445f8d0a8e9fa9584174305db23144e77161f5de3dc5a21fc860b2cf95182e8d8546c421699422440673864f9f9736c072dfcb4986f526b0656d81168bc4531e5fbd8b303a5417d1bfad9b3df625265eb40883c7c63fe80c4b61b20af9a1b17e29b949812c16eab928bf399702f219d15bbb3f2696c67a0f4dad4f3035387e8318e7db035d4645120d7d3931c94cf1ba7df7ca667c21de127507a528e14fc669dbb5a17f3057bd378153a074c110c70286240cb24f6d81b5a33480c23e2f18ea6cd798c9647ed25bac55fc12af139d67aa20b26c27a146d59b217ae50fc46cdf5f6ad9a2890ddc3e1ea7043544a430daf8943355bbcb2f3a0f3a91d6d9dec7efca6c0e2044ea5d66e3c45be71f16ca9f25f5d26aaf345b68184bc8349c4db745524c891e2ad0fa3ba880165608710b81bdef69bcf8cfe6c4a129773deb4a3242778917a4d9d9bf79a7f527a00d496dc216fff2087583f913e14e6ddc04d5ff47a240650c3318bac6891316fc81a0a8c18234947ff4e0a9feb18dbc79e9ec983bf8a6e596fadb1dca0f7839935f61ce83793b72a150737dc2b6d7e9d41c2471c5b2b685a22c92b94c2a52bd21199bf421d1a34372a5be5030f9d060b41a9db2ba3ff11aeb2f36355226a6010a4068fe3e4d01c06151dbe2743a07e2506c39b6922985bbcf94b35e90f8f0e0efbde44ae09c2d6980fd3dde2d61aef719a8f20c0b1deceb11563c9208da7fa4bbf65e8b1d3d04c53913ac94fc483c0082fa0e4f5e77b2f8b99baf18ee2fb7442a5db39bae6933cfaa6199ada7101d49600c2818081c7ce77c5b1f7ae40a9bc07ee7adc92217489f027366c345c9cdd61e4e231149ccd985fcaf8d4c6ba261f62899aed22a6b867897117afb237f12a18e848c77e0a45dbbc805cbcd623ff35cb6218e4f5a88e91342ce7d442d547cc09d2b5891e420ccdc13a750221c625d93462dadca2c1c3c6ebb0e623b1dbd21a694304567f7e6d281a7c866a0c2f3db167a10e21905ccf9462e0cb70219f349ad3754ebdccfc913e0a77e41a9842bf5fd32f781ebf23209c131732e0f0b82107b5a69f713e9fb80676a01792e42a8b2daecddc2e9afdfbf30f3be56031fdd973399e6e359180739d368a8782d75e9ce64a688b76df0d99a24476a93789f97043b33bc9d8822908f3f0d9e756dbd6da2d8e71d4da470ea040fa17874df81dcb9fb3e4a39fc4298313a5a7913a03cc25a5d6a38e65b1eca7a25d4fb7218ada8f8d9eca6d4d4d29fd78addff97648ddecea;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h39c044f5a773a64d4754ce034421f40ebdb1969cf54b692c4530a84fe7306bf98621848aba4691ec1a7ac959c66aaccf424477f55ed3e5a3dfee9a2abdcb93bb29e59716d69d4d0365295d23bcc5f4d5d203f3ccbd1e77e49e96a28b2a00485a996a2be85cc7fa848f649d0c1a98c72090f737d4e2c72ee54211e9065d581985e83203911f1f159cc3623f5c5fa13dbe86514e1045a4b295338c68cb2faed24ba265630113001fba767a4930892bb7311ae7263111bef36b9a22406c52d54e53a14042464598fd5cad699401ed3797d4f3cd2e2c63f0aafe06f7feca1bfdbc7dc31a05e1930a920f38d8eee0128f82a3258080e28a797a30967c4fb53972085b97c9f4c179b465e1dc75bb2fc19d5f453751c98ddde4e99030cde03683868d1b93a29650da906d10f2b07a9cd91b7009fa6e32ed7bc97d7e331cf94829e02fd69d8e03fcf0dc701962c5d2947f76435c36a0f8f548c9b27e65464954566d3c68d1db824df31bb9e73c363c44d23b4f046ed60b0da5d72797b283b32d1b0e7e9fdec12ca3e8c88807d16febaec306caace37fc4eabe3460c29f2b2a19c5305191ac1cbfacf61ac4754d42c6f9874a0bec20b5a660a8642f7ea017e98d3f51704f268956dbb56fd80ef169d06435f767777a1b70aa6acc32821f4da355e69e18e61cdf7d11591c386f931cc0c75082fee91e7749825a6eee603cbcb74c39e2145dd3f108aa4ed872e21b8867c29e172dc992b7a7072e711bc68970e6ee97bf96daa843d02b8524c1e4ef0425ea970f16d8bd5080d9431485c0301a6d875da2afa449f6f59fab44a76ca7b9c0372c15371740b5d3d6cdcde9dd364fbeba52e8aa6ffb5325359cf6d82209c22c30787b33bee68bcb4c999afd172c016bfd2b584d34a60f56af18515e3cbb552560858d2b8ec13e9ace110a68a846567dfa2a364b174a30e2773f5fac95089b1fc5d853aaf6cec1b57fd37127f61e4e8dc0bb60acc0de68600a5ae1765a7f061f1f18afff830884c490b25046fed6194856b28b3b4c16a1ed687557c3a0599a9c0fc39ef9a8b09d956ee412252fe9eac4add8a0329879a7276458ef649d75910e435f317f3e2ea7dc2b9440f4670c30f560c6f221c6ce4aea93915741a85c3a81106f731b877c48374b9746565a44e872ec24c96387df65440af331d7940d8bd19f8947c89c20e24144a8c3a88447b3eaf2d32a4acc5fddaf8ea2d16f0d00c9fec067b3cf4907f05d94eabd249d614ee0a27d6b4cf5e03b872772dcb5245f2c91fe9db8f5b20cf5613db6ec12d26b9510934260fdfd74b2cd0c2058061e6432e345917f34edfebc17f701acb0c6982da35f08ddc9b77646a4033c77bcff2e7c9f53fbc84b74dca9ddec02641d1fcd35f905d1d7eac9f81a89b14b0caf526d7d77550e25c77b2fbe0c74f3b51a42833a783b8e8043c304c0884f9860a7a9361c0e329c5b49ac4472b6b35dd98e2b86afabbe727d4ece8a930b201b0abed8cff385f991ff8de3eafbcae3f2a8e4037e5dfe93c83542aa55e894e5ae9755686e84a738136a17241cfb15f1309fc44ca317140903cf64df43c98f7f01ec987c0f487aa56dad8d3c20867ca6e38adb7796e6b1ad035d8e7e5a4d56a39f76cbfb8066d2c0f6f52d86c9281b52b731d7f57e4fd32cfc73210e5e6da86b919b05153604cdfcc491c8434dc0158d7af09ba3320d7f95e2b20c08b212ddc5cf4c3ac6d250dda638564b210bc25af18fbcc3cca54d00283e24f1d198f1c1a61f9d8deda6c9cc5eb43ee516d99039b5222194666ab77c7eaae4f1bc93fa43c765de8d9f87551c1a0abc80e7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'hd7ad4bc350417bfc7d112c27c52ff163495c445b57f06b85f4428412c2fe34ec4637a9351a6004dc4ce651c571ed9cb3bdc77adae7488b04aac2a7ec7c28803a906473bf24f21029d0581c20e75f73743a4e34a067250788a0cc931c1e14bef46c1b331d25a6b9fcfe06d6841be17aa06233fe94aaafaeba51d4b4a9034f3440a0c6988b04ff9e3074ffb76381e7fce7ac0b6beeffc15c0459bb42c63d1f8c973b6f123efcea0427465a680a7673a5390346c176e43f50e22dcee814bc7c2f866fbce25ad715f4a4fda0d0fc297b9760b34665600019b83ed0b4f07f815d0da1f1d2135dba3bc6899392878f7c1876c6139bdb5dd653c9b5e249cfc725d52abe361b40a8e94bf04a05e6557a869f8fe59f9a9c1e0a2ec73c7e5e380f005c6adb7bcd0259001fbe3a46a41c6045eebc75677867ea4a927604211f96aff48a63c674cc387b0168cded136761cdd894569b90ce20d31f877f946ef349de8f90af55b72184cbcd7b973fd793f5f0873f56142664f4e66f2a907e52371b8d2c5f74bbde04de230fb042d278ffc57f38129247a3d149ee064a43a076b57a55548b100b2cef6317ebb4bb935a42e4b9d5557d45c06c54533a295d4728ebd6fac0ca6b0e1c12cd219dc70098e45369cd8542539e33c40583e13e49bc8a86868df4a60aee0f38e31df1b648c48b5d51cfd5de641301132d1cd9caed1c937526a5ca75783184da3af5d05397d6a6eb4a1d27db4eba775031fd7cf6f5011e635708b4f14fa6972ac7dcafffce65046048cc3b54b929690f28341fbfc35dcdb7a4ea18ea5f2cafae483fd8d142e28fdddf3d94630c3afe33d6e1d2ceb31ff666cf4429c014c5122208048563fbad39ef8f21db40467e346bdefd5fbf559b2e44a71e0bdf025dc1a7268028554d997b94570f62b98384bd3e6f43b01a17ee3edca21c6eb80da1621c0e6e0faf3d10b1fae1897d15e84d73651981216f9939bb1d68e91f27ad75803b0e42822055f4268f5c959bb875a9ff3b63030a80e5837fcdf2a3839b5d2858a45e716e519395d52194937de25ac288a0e5573e2046105281a03e5b7e1e0ccaf2ffe13017c5a711395b9aa64c49e20a6a14c10897147a676bac5852ae04c0bd3533afedfb7aacfd92ee4d5b52ae0d496ace76f2d3424767426e8e3c8cbf86ffe79a833fc7dde5b4b66240e9530e9f79d2bac68eed42e5c8cafc82f6146948288f4a0bf9d6ed8e52274c36e9afdf1d32d6e8fc217092a977773b57b147dd8bb5792d60189ef65b5aec4f9e6e1ded98c762db47e843c2040b22e5af6b07b0c6808fb841657c7df46bd8aa26c669b13b5d49afc5b412b6f151c4192166a8713557f3194f1df61d6c0e138c787201c0d0eb436389bd29819d6e14a6d18ce9bea0aaebed7006bde55c226bc39fc8d2d508aed0ca0505daea10bd5c8b5c3f13dbbf7a568c748883db9412d11fc0488f82bcb4e4456e873ec2e9a6530b3a9656c8b731ae7f86042eea81ee9fd5b1f2e05973d50d779e7bda5597345f168780dab2067fc1c8aac9e80c10ec1654f02d21068e0880be285eb9d015df7db6f632fa437aef0cfabdaac02e2e95febfe56714fd0e38119d01ca647251e18cbc7d1d2c037ee27ac374bd7e9e0936c9e3434114b1143ab8b82ec43d2a5bab6156c730f8c7ab3c27515e83e69a6d54142a32723df7f14ce774d5d3dfbcdf67a1826cdbbe9ec032945a72aab159fde4921c801e9149cc30cdaf8e6f3ad6c9a8a78b7b337ce808893adeb329af1376c59befcb74a6079ca00e4561223a02ffc58bc890bd595aa3c503761789a87e5b626bd97cffcfb2c9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h2c160315509430031af9c58b63784c0eec9888fd718b9d69b6d735ef05ba43c3f9c94d139e9c70eb3cf005297849cf0094e61c1cab37e3f203ce82d4123f655fc65f432bc7752291219c8c8dd7f007fb5a2f276ae9e7ac87ef224667742326821238f0dc60ce037d52dff2c682f65e7f5e75b2289dcdf663d6accbf0d0ed58918f5b66bcf0584eb91900011d5f05611564d6000f92e5ee27ed9e5461d643cc0b01490f6281684e74b85d6c5d25f63558e915fa96f3c08fe9c6e6fad39170afa160028abfaa32bb6c02a725cf9e2ecfe63b4f15675fc32a1d60bc5598297f9b42b8a0017cc9c0d63bb20b360b94d52019f283d2c2c2505b260e9ebedc78544dabe4bdfcf8e913d240ea59a475891e441ee31e67820e6e04932bd01d60159518506db3b07ae2da4dcb041f772132dd946f0df59fb4fcbaeaa1ad3e33c9c512b387ab27fa9305afa1be0a148af44f2d3ac1095312afddb388bdd8b23ba24fb1b89140bbea1a910b3efb4bff6d2f7078d8d3408453d70c953e6affbc0ff2ce026e5b1ac9f74be6b05bb267b84dbbfc93f0dd73766f64e863d528048f1081700879c0b28f45677329239e7dbedc808c4a36d935d3601ffc33a6df54c66e9ab7aa459be710a0f70d0a95301d3c98d055ebfbb2f3f26b53a54bdf5c3fb1e89a16fa3fa34242c107cb41d06e4c94c75945079dd4525789ca8bc9ec10961b87e869289848f385ca5a4fa3201b416385cc80b9fdb494bb7a02284921517161442baaa8af3836d0226f7303ca9d58b1f1c4d7a0dd09bb48d8a400b84314d067403b7b3e1c7d3c29017c7c8bec7881fc6c6397a1501aa2b30d653bcde1cde50ac09ef67ad220ec559ffa99796f590627dfbb0684620d2a7419158dc432212f8c9537134784ecd6aa8b1bb52940582eee2706891beccac96d1f4ef44fb484045e92eb3c8ddc12467ac88df2e926f60787702d532ca187b6012bd708bbdac543a3211c4294c9386e2d94fd951dca779abf49cd556b0d5d0e6ca989c9f755e37bd6318c119469aedf98747c5cad36a4dae5c4cb1f708062dfa953eabeb290ed031eb4c72ba801175e581663b220899a13647c7fadf40efeea2fb5a3f922a17338b54c8f16fc406354da6692f9c59ff858e4ee50b2ace21de15a428e8abc8a1967b9e972bf771308b799dc93cce0a2ecc431dc17179de66e406fb2f8213507f7a9e8366f984afb05f855bcec138c598f4dc308b2a6fea0d0f8c3ddfbf5d0590aafed8e5ad7c6b09737301acfd9541ecf46f0cb8b6c4b6159e46a604aca233b4b1f359f09ac5b340fd1afc8b762e03e495e794d928fa6fe1375592067740c5ec13c37d95c6751a4d8dd434c8d7d5b2b06657f9141989e67c4111ec258fbd60167c97b39219d2496d17de1bb75c9f14cf1a1f911acdbc45bd0ecc7aa62897ce9e24f254909ee4a1daffcbf211dc8cd7f6bf92bf218c6bc1633fdb27182c20ae6cc347de9caf4d5d3b8e40bc5bf0f838245aeef6ddba2c5fb4a0a196e00a23aa4e0f2e062a38878779fe2c3c4949e18ad5781c0192b46e872ddc398aa112254ed570bfa5583edbb9b409c7650dab52eb4f6773b882e6ed17f83078a79e851c91d5262fc91540d47859738cdd60a9c96cfbc38c85e07cce50f59e8c5e8219f04bdf2919556b9ba4ff5a222b20c73bc265ba9505eb966dcd5a6a153fdbeb98b89157eed2a93194bd821ebe6e792127ab4016e4c0ed826fe20631adaa4c14e352fadb2fae6b1a9515f4e8a1192fe5e5255da1b2c238434e97b90f4176f22f7839f7df4dff8776ad37d2beff6c9ca64ddbf2d2ada86bd16ad21ad85;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h3f970592e3143b498142a1739ff36beeac918fd575b8c5f3a26327a544e3e7f2f4d893d8450658f967a9f9b169c939876d33a3574b6f71a3246cf309ae2966de5d729e7ea8a642e28c6a22e2de43197ebd835f58df6eaa999a6187e81eeaadb0dd1b5eebba020d7e5cdbcd54189830237f665494fd557b6a27646a7ca67edf52ad334ad828c718f756300d13f39be7c540e4aff480a828bad84c33c85ca024313eedf97c04b1f0835b43222026271c2b5b3f0bd2e1857905a0546599766606fc09cc3c6e23dec6ef51f3538af525a0329792adc464f0fff6837ebdbc38e8cb03829bf34db4ecc69b790ffbb21ae237554b28715b8cd3e99ea5175c4cb7d7ce071c81773fd59811c9be1188daad158208dd396ad8bc44093ea214f8cf240216ba45d114ff409738eb65bed0ceab4a826fbfdabd6dbc2906198346c8e5e9c263c7e06d8a1efb0702109d419e307b54b87b483fd3c3123189a3382131da1dd968d79d76aec3bae068be6c2e7e171f266eff7ad050c175e73a3689cc587e6a08d939f7d184d5366cb74f0598980fe3a4919cde3abcd42424871d51cb15eb0cff5a1f817ea8b90c54da77ea6eeac14f693b15e9296b4437b91030cd130c634f19ae587b22785e17464448b792818338d1af936ccf419dfb5660cf006d0e6450b5f761ed090635ad2a57adbc644cfe57ab0d3512d7d647e09d8857387e1a8a0fc5f0c2710010cbbed2af917281315744980ba4a644a27ffa4dc6b42f5811cd67254884a1cf14ee84d35ea82154fc13dc45892b037e8e05d2b5808ef09a47c6b713a51769b09f4d6053a2cd6d5d3565a45cb190c8b38787bb8ba8d499d9e370752365e63a95b13f85235edd8a19f5f06c42ea4b48f6cbc0f3b84e7637199766d4f14ade41328dc8d7db039d1c14fd5b16557c46ffe4563e3a63ff53f3b103079616d0eb9148e500e91542322c0900807690a5f9f3bb31c36a0650e7075f7ca59a9fa9487232b18d56cf061b8cc345986ffeb97ce90d4b76e42365033099264b375e945e34be5ab6951451916be679ee014bcb497bcc4f888c7310363c1ee23a3a6e8a9bd5746d5e8fba0165a8b7e7d658d4cbcd20f34d25cb6a79cf5ef62d70ec558f8a019c8547e2dbbb1459633ddc6949e0f946081a40ef77c104caea6b3e7fa0bdb0504833ee98026bfa89ad925ae73eace3fe390364650e8ebefd7c7f9a5b4073dd43a7e1c56b0a000abe4cf711f8bb9f9e7657fc510ec0c435655f1571381997b913e9fcf37c43b3dcde9166c125c82fbfd4640a23787340989fae77526710e2611363c431481a27f2c6af2d21f4559f14cfd661b144bca11ecf57dee62b94435d1db12405af103ee702d071e51423dd96e5f2431f1a7edbfe66dfe6fbf82d8acf058c44da0332651d8c3794f7c5095622a965b996f8c712c93282efe4186556c7d60cfd6608f47ff0e776c23dc89126bc6e6291f3515c24deed7f218cf3b3f987b758d045388b72b9d4dfa6b5da99493e90a7bd55896f070a99a5a795bc133ff69784cb3991f551322cd9d0e3f3eaf418822b4ccc95109ff7aa4dd941de36e38aca331b3eea707d5740409ffa15d6af5f8cd483787284b2cc4a000c1152ea92f551d97d7bf12712633672ae73fc2b5a93e71bbe23adee34285ebf757a95de467654ad57e892e316e91bdcede4850d1904481e07fc8509f05d8886ce032ccc7c119ab3c48c59fab33cea4d56b7ef2f4e7817b1876fbf433b7ebe941ee8edb7b844e109ed20bed50eb80df55624bbaf2b651c59636da26909d9042ddf16a97544630b81f21e2750a1fc670c849af8f911d2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h15e2a088f4e9b007f91db53f99cb8e5d287a0f086af42e368be532e9ed75037fb2908917d08e11b52e958827596af6980eac0826cb359e1878669971a500dfadd48065568953e2a4d9d158b804806d4e110442f595d80aa555f5ba79ae808e4eeda0db57ae94eb6fe505c3bed91577a6f05a9e9b022fee953f9903215932ea2fc2e652688edf9cb5d65202821f69eaeab6efff16d79801b2ab682cc48366ef6bd4f0c7d435defbfdded3d618f4aa41e05f0fd7645a0831b8e70d47b8691965583dc1081d5de00f207c3b58ae9fed6940fd1fb31d2c2bc47780779226f4f11715569378272c475c2c4c7f213d97527c7cb660f87c5cd3874d5f44d4f84907b162c525cde7f08a2b3758a1aa3af7e0c6ac797853cccd45ea3db40904560dec416fc1d012af36d9ccc420ef1029c60a73b59fb2b2ac292686e5596838759d9a676ccd867cd55b9950b1009a90852a33ddff5b8b2f8a791a81a0ec3534a2f6ac81aeba80e1e3da88f0e0865bffc26a32424fc56fc713e617b36dcfed8b5767e5884f8ecec7e17ea5a5c5b57994cba598f99d76c98deefc3e0fe3f8b707ed292363a79ecebfc7058e521b2093eae1dc9bbc170ae51c498e895654df0db753d05c0ebe9a9a9623eadb77a43e73fe2dd8d403cbeaf676120bd6c3b447dba1c39f4c54cf17582efa8d0fc5ccd14448d14163e4a0d7d5ab08e00a33da9ca30f66d4eb816f708fa081e276c9a114b68d78c788c8cc17e74066499ce0ad6d2d7a036632a7f05d982730d9c8e0b79db6648b5d386d6d529a75791e7d4a23f160de631e642c13a148595409fbc7a57beb7d7137fe77d9254b1f9aaa3d89a0dc33c77288a8879be698e0792a05120d8bae803306a4953151e0b856e6e1b0eb50ad71c9f505ba7619cb6fc6bbb945557a16231e35aaefe476ca8163653d4c09ad3cd390f3ce5fb2a2892e4c798d003243585e996ab05c395bd97339a99568c72c26895c694228f406f37110443f2ebc2b4f7dd6f6e16ad259e41610e966c9481ff2a212784fefc15ecd15954bf02fcea28d9c8d696043dbe2d4b12fb3827f765ce0765a6b284bdfe281db6a73b1619a7eeb828bef73a5d06205551a4df39df170591305f514ce81cdb392d33ca1122d441ed66837d003f18426f290fac7d502513713a0eeaec592b832b97fe7da5981d84e89e3c59fe0831fc42b66af49b57f517862ced97e0e5803a838dda390c705149eb7d6a2eea2f4652082537f5f456847c3e512b8c8dfa4b3f3e026c9719a304e6d296fb5d8630cebb11aa8667964fba91149e28aa18feafb74556502a141b498439e06f3d180436a13be59ab8b5bfb26f1f44ee7427078dfd05bd8fb3b080c5d0dd686f13e1d9345d65721452bc469aa65e09fb887981ef2f1f051ec524e7ae6474995834e01047767447ef2a0057f0e01fa984b7e05ddb076ea52f3b692a39b761486c0b2eeba55ee95eee7ebc509dbc1607e31ca9603cbb7171dc33e2f227909293d2d44c14c6d969466ca4ff5dc6df16ba734313c47b7817626744818d7ec4cf011ae9c32eb5a6b57332dac194e27446fb5ef7c0eb3c9bc08a37ab5439d9c568c936874f841fa53c472f546b01c11f95d55adfa4679d93b7af1156343200e76ae189447f9f7ca5fa6e6e17a2cc9c350f46ad271c81922507780ac7d355343e4b9230e03d8e9ad4f78ae19d8bfdf6764b4e94febe5b6bd3a7d99cc8caf712f66d28a2eb607fc1e4ba2fdbbcab08d44ae776dc768c02b260938dcba7ab5ce7b04d74c94bcf2f00814cbcaec74683007a011adf6c2d06f1a720a5b385c135d6e164178ceb5ed28;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'he7e7941d4252353e2d366e10751f794490defe214c6df3a63d8647754880c9cb6333f485caf06c7fae6d4ec783dfb9368b5951a9e207e6c0a20ba9b3fb3a90a871c8f91a7a25a9ccb429920b4f87b616b67381bc2beb9b5dd5c61a99b0967a26c116f02906b5b3e59b703cf0a9d3645a83c12792dd51d4e8306da6affa4676c9dd4d9bc4fed0baa71c57d62f5ea9c53ba3a0a2e202e0d8e74630a3af6e244af0d1c4112edb1e0dd0abc4e507e9bedc9fce0ceba60495d94efdd845a2288f5b61c58ad65efb28b95dbf2086e1858b057dd0699714926ce23b09be3a786fa1a0e3452310fee573173ae46c7dfef908035002ad2101c07e6c754867751b08dd81ac3c7118cee664726c8ec069e2e4598a9749389f53e27fbd3b10c2fa5fa47824314dc98ee9a4be2807f45f0e5f567350370450496adff29529151b529bfe5666e583e57a312f34b26d88a162f9150bfd2c4f5e6d3343a30817eb742f4dd8c3ac96c15aeedd2c90047cb2388e117f61947f55eb509a76cf2ad346cc46ce52ba7fccdd7b694aa4f5d3d41569c53af6c109d363d10e0a2cb6edb3d53d654dd68d460ae59b2027e6fc260f4f239b8e03cf35c5131b8dde6ca9d1f4167fe407cf7bde43b60253deddbf8c53fdcd1bb464b28f57046c64b7a7303c1c1d0e2acf0f70186a29ec32e42fbb9d9aaa2368fb7de8d47a7613548416473a42213f6e24efa20ec11872005203dc3cbf613148038de37e326640a3a4ec847e770095f33bc7717813ef776a1692fedf1fdf18036e4cd5b44c1547a3c91ed92d26a7e0e0e5be78e9a7003154ca43339c6e3d278ab2ef80882da80295835034ba79ddc6a447e5fd4f20a1ad557da3438f5c852b8e6ca24deb37b01fd199cc6f4b791b6611838cd854968852f0a5e5ba7e07440ec4a661bc682e2bedef8d50036d4d4b00a21fd2190bd840343bb766709708505dd7d8e3e44503f236a973bd649cf675a4a6bcb8f2369b945bc597d64574c1f391c6276318d838ad631b16b5ab7a9467b7673324f3e9686e66c6b07fb63c4abc8c31c9b5b1e2ee920ddbe2f70c20da508213ba3faf276442ae570a1edb1979771e19e2862d6cf69a6b99165535a8326c04d207f991424b8325b530949dbd3749fea77a32444d3d960c88aedba4ce18d61f3f3f45e9822feb445389d504a41d33c9b377b15c1778bed8079d94f90a606d36d151c916eb93f854a03d7c9a850ab2c8e97ff3e072228d47b5668fc56793b873cec3374e807b4053adaaa95efab501e91b65dbdc6e373df9bf20fdbb7bc417f97569df42f75e94b6faff69ee6ec41e3f5384e6f918d7173d696494b1eb073c5a31613edf5e6b8b380d7e964a698cd9a981a4d7c620561a2e8fe1a7e77696d9b4d34c052d4140265dbb1fd11c0c0c51f21c5a833505d659639f5b81941e246c9e086d4e5bbaef4d12f3ac24a77f0e357215a2b87cc794171d998a654b1090cba9815d34b917146168f1c46e480092c627f95aebb1a130b60738b636f9f8fc4d725afc7f848e714b9d3b3765a4fc53e0d85e87802fb0e0c3e0764332bb870ea434609c3fd94b418fa8012536c7633028bbdcff32ff4c18c4d407aacba41a30109e9e1768b1f64c0ad75ac1ce5c308221e6351ce742f97f0cdfc11e85eb8baad97571c8eedb223b7f0ef6eac33c6e4772beabb941e535e833cd75170562de668c05bb359b7dd74f0653ddd8cc6f0be52e0728bdfa72cc704d22fddb827810e87abbbd40d7bc68e814862260576ca39b9ac030c788bebea966503e92802ba4ca5765cbe487a7ed80a5638213246017fa2dc82531b1f649db;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 10368'h4a7aadc2293bb60238c88cfdb26247b834b971a7b392fa2b1cd96b6998d15015a102ed4ec28849872d2bfc424970208dad476f74edda7b3ed9a459b14ac33095d885bda361ee08ba41bd61d07c0b260614d89518efe7d6244a00d60262599a73e5c26bf0d0aa0d690a414e274ac8fa690f62840f9cf96e2a26275bad0c9810bd1a3c02bf5c2a7e601e823afbfc4617e559aa0a0b875bec84b6c5053e31422fb88e818441ffab4c7035e2a316b0963cc732a0801c191ab9a4033706174b420ad4dea4cae6c82fe8347fb34d67e694111f5b76219c9e5df0dd22a87d0acdb5f543491344c24013dfead5ad91f5bfcb6a39d96424021fd26995a5ac31bb4e13c54bd9ea1c2ee9db6e6a2e89abf9ca01597f0523c0b3f72aff7d1e350ca3eaac7beda27e33f1c5ac817896546e7e732fc3ff4f48ced2596df7613745ca621992fe27cc5b14d218d57bbcf7c68fc98e64999d322af4b057d1799f9cab7e7d58cc19e39db237ea82f886d2e9bc0f2f8ee160e253191d5faf151e189d64cd84c13de5f39ef038624f40820ade936b03df41c29e22b10481b7aec1619f812464a914d058fe8618e3c6f801cbbe2ee3474c9c073ee17b1ea05552cc04de3306c353d7db492155bf1744d4a40dc2a5aa835e07b7a5c715fd65471d4e1a360f484bb37b8314b95ffccb62e46ea591b941593ab10f041b960db65860c1bc9c5954c9078fea38a65c771c30afa89315b891872d10df6da60c8d050e79312d6a5b3944f33b82a01b8ea6f26a297af2b2c81cf90eda61a37b773322768c9a8280139f5e2215ff79d1935e50d7df91ef5aae5850c887e920737e47718d9ccc71e7545ca73681193e850568badfacdc0ebdebc1a6c7e6e94e8175846fbdec6303e58df89747ef7fd79276df33085b6129f358bc734ae554e700aae5133ffc314478ee86f76acffa385244f469d1a4649b551628d2a2d485d773e94cd6eee95a5d917458b084e7388892eb1e79c3ba8c213db54b3dc8b867e8ce90de33fed777fea28fed4275385a2699ed56cbab6aaf446432bc95a14d2b98fb05b00a011b04a5fe68fff4862c4cc34d03bf1e3de4d8fdc7142e31d25fa1c0a3b953e6a7b1de2190b414d908bcd2df3c08039831b4dee7998b0f71782c90edaf45a5c73fe1e00cfbac918f5a43e43acf68cf8ae353fe3e3de1fd4f190fe0a5a77b5f00fb9d7b0b43ae19468b9bc2325eb5a323f9cf98bd94e285244124d2119e3b538f49bcaefe570192c6faa4363ec34d90bed84f353a3b6ed53e5cc0b667587aa993ad9ab912522c5db44a0b7a5805204b4f514b872b058e03f45a8c0f332e3032dffafb6f76a296ca86df5c0ecc724f13980ce8da4bcac28efc0bb0bf95f16a43587043eae5dc11292906da868f779e2e4e16dcb119078461bc9eeb879233b06efc7fd3a96320adce08b9bed72f75ce18928ca6599356f794649fb1ec10364b3db93472a4d6994210bd328fb2c09fd69eaf08b86a40fba08ccf8783906203afbd8c227bc4c604832479ae857b6ddb4eda1ea9bbd64af872fd0b712ea22d9afe6a026535b5f8f3be9cc37aebac57d517d7f9655a94c700864340ab645b997e23928ca8d6c85a779ba84c26e184e2f2a1d98b812e82033d62ecc87423387693bda335656b6711b17906d5030c9afd27ca5293248a0ce944f2b9e9a43e6d7ca3641b3726106d2956d6307739becb43f94fc1f06fc577df906cdbbc24e9b400821aa8d2693bc06bb240b5dc86841f4510b12c9f593fde85fffd23dd6c6fffe10b7aad66dc506e4ce138acc37356aecfb0b41630c3a3f29fb6786f221169ae32;
        #1
        $finish();
    end
endmodule
