module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3bd821f48209406557b24a33a79b4a56b52af03a8f848a7359e6f0ca0a1dd44c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4461c167fa801c774914e0871a06e94e1fbaf9275e5473f6f3170974f980793a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h166039d0b78e9f34d28d8817a10825bed38006618c31c20f8070fd88c1911234;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc875eb6f1ca302de550688381fcf7db713d69857c423c55eb908d59d2395ca03;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e566da2aa8b5b53290eb46e08f04a5c787a345078f35086fc1c45fb999ac125;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb85d5fa3e1b24b05ca140b70437e00285920fbc5b8b3e4cfd5c18a22ed24690;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c4230681616e26fb3d824125a8ffd5add05287a0952af6341d3b393be6a603b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ad438779ebb03b8c2f5ec98ff6d4856241a0245fb3aab04d231a44e38d880f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b3dbb94c1222fa1e8b4b7f94d10296065d339b9243b30075ccfc8f631fb093e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6140618f801e30c34d2f1371aaa09cb860aad305d483877290f8171f49d3918;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hceb036755bf1afd5d61eaf184eef52f7cba62656a665a16ce6866b61f0c762a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc579d75b8622b76f52534779f76c29cb8f3e8ab74151d94f900abca6491d9396;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0049218544408168098bc1d03153d59e5ec761082aa43117d41efc119554530;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61817f86e205c6781757fbc8bf19e9821b7994141d554b26ecd613310ce209e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9822a6e81e68706b4d952306ebb909c2b8fcd684073acf8cb35236797f75a03;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb2c6be9c390a734c71c84abb2eaa9220f00fb2acc32f2bf535d777fac037b631;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3a239211a8a19fa08cdad4cae28cab9363c2d03786a73557f7d8aaccc1cdb04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h117105c29fd416927dc7a091aade2bb1a66b79b80f5cf4fdacd5ddff8edea9e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb842071e8fa4aa7940d0b14a471464dda300166809fd707306148e30cb564c6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63dcac02597bdca31569fecd304760812403aa8d0ec165582d3832f2eedf35f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h201988e4232b2767a61531b1392589a5ec9e8a90776c48e862a69cb4b3d2a69e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h840046a1c5bcba5e16a631e08b356d04b309b2bfdb45d50d0ed547fbe1decd68;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc66baf4241fd59414a7b314943aefb767957c477824ef822dcf823463667e498;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5809686c6cc67b4abbf54a09a280901ae0196a0c6c4c49e2fb3f40b31d45e2e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h766b1056f29488ba7d0b1378340076f2f123986fca740af84a92c0c9af7f6985;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5f1fc19dc4d9c9b0b8ce59d3afbb6b3599fb2e0e0ad77dc87efdb0a53fd8eda;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7e0bf69c4e9e8fc3df45dfabcd4459f0ff4539fa9411907e56027f910f01e5f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h79d4c26c946d6cefe0a001e6149951b7dce589669a46266bf8522cee610c5a18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8871bfe660eaf366ec6e6583ad8e8b427564b48b120672087387d32ed97441e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h540dfd7acd1cad243b354ed9815ee70f02978d58337ebe2b021b496c8992ad02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b91d7529558ce3c5306cc0b20c3bb1945cd43f6616c9bb029a624b975ac20c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96fcb26ff2c7237dc9dcb412f9cf74c3e99b982416559d5241fd211c22d4824;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55a2b88dbe13fa89c115ecd05b509964a5875c677723c2ad5abd1d9135f25d40;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7e05b363c1e4ce838ced5e0741490f36b2994a99ca03fdb5d6f032a3e49d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc852cd745ab316a046c3ac974a936fc9853a2da089b3e51e70d075bdb7a81e4c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71c83fa7c23376103f7b2d89e23f38ed555b976af1e4284f14129391741d09bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b253471dc52b92792b387ac8d7be1bf79c67d1930311edfbca439d9133bad54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72a54359f972968030123377486da0a96247f54671f0442bd11ed233d44c1cb0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcbf51c70464b992c2763d9cefe0b31d2a9c38afcaed0bf22464e848c85b726fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6ffd9bc34325a20d481db7f13fd84ff966f1abc50314431fd99af4450d957f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8255d73a4b49b4b65c4d8d5f2ba754f440d71200bc4c59777737786122da1cd2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd029ff962199b0ced24cd3b7da5e2ff84ae507034b1ee737d3e8fd59c667aa2b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb54b12ca452f056a752cf5421f939e9eaf60a2f70cb081a6726a7008f2a953d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5392fffc8d598e279ec398fd3d432ba03820da3a3aec89d5ff315f695a8d6a9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a07eb11f396f4eb98df81dde95bcba3e004aab5e1e2d8d7d017b28d5e51bee1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44ba4d5db0fc24eb1fcb349910d95f8844d9b7b1773245e126b769fbc5278875;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9acfc8e8e39ce1ca8b023c5924c02564ed5685534947c2ea8dc62a92d1deb4ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d8844282d145a6d926133a8f77ceffb71c0c97e571ee87f3d017001dd28cf2b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he77e157bb8f8f55a072012505112b9ccdd1ca24dfcb376f168e1147a01889f54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46def21bb6c8cbb7d8315454afe12ca19c3fc8ccbb3ce0d8a144781d34b0f051;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5af7be72569a8b2e059f0d9d29f442cc741f67f0a2c833c17237839b0e8fbcd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6885dbf421159d5c24b0098fe982044a8e5cef8579c71d949e317a6f23a6cc4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef2a379fb1fa09507bc7a2082225f33477effe568a10be1c33242552c5898d9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb8b8792787b60eec96c06bbbbe09d197d61c1cc1cf8fbb7f966d5949d1b08bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd9d5dfaa9d90b2258077303d2ed2f7c8e79a570cda190d6617f11bf8709ec630;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h405f5b28d9d3a63753257ca85c9d6769ae064b22bfb7f820b8fe5222ccb386bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c15d0e75726c19912afd1a821727c6c2ec1760c462ce6f5869e70b7829f9247;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7de52b75a582febb9b0579caeabd5c9dd543d5b80d0f66b265f1336fe875c6df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h931498d4dfc71c9265851663a6bf91f3b0203b298d06f1a87dc9edea127cbf94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2cb1c1013972adc4231c3198ebb3bc755d1e1cb667e3016d4f0f22980720f91;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78b92e881b9902bd1a506b11adf9d4b7dea7df725084a5e3c79132cdf0ced09b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h67d55391e863cb59b1d6ca4976f147f78ad2834eb80202fb98b46e2a01e55ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb6127916b0675a88d6f331c69671e42a188361216ea45dabffdd990392cb2fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h22a0e6d33f14d986fcc009d892390dc4d89858a9b1ed38f151306a5b710e52ff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcddf4851c3aac412a3e813b3fd0ea655799add9d637230481063904cf8ba6003;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcdf716a900b593cc2b230f714ad74beb4dae3549c69bdae4c6ec301a0b011d7d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h980eebe5f138b9f164f870523c231f357d5060b33c4a674e03a4cb0422508a3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c3840a0d2b7d8bf98e86ebc4286fb02a1667aaa5ac3463a6338a78e6fa55661;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e687e97a37bb688c2354a2d1bddfd54216c02523984959daac8897d793de5d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h284d3bb597a454dd2ba0e46eea78db0accef158bc5feb8118aa3054ce9e8b62a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb56613fe7ad7abc05c727ea9f62036467dfa9c1db237e35c44c81520acd30de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1a0ea28920c54779ea05fff5fd3c763aad19d07d6ff766e82896e181f505edc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3e24243fdc94a085b4dcb24be0b5700bee8f35c21e8bc826b119c8c73a853a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24c874bdbc9759ed2ebc22de82fcd5d4146ea129e658052d2c0ae53c68022b67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98d5d803a45263230ae26fe9aafcdc5e9f1597513a68566289b4b5d90d1461ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf29723b2db05864f51b7af0d6cb9e45fe10340540b80d9c8122413a730204490;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ef4f490b3a211761856712d8f510d61dfdbaa8738267f5906c0f47f7be9ef67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a112c11cd387ccc0ea759e4fe29ee94abbc37ebd753530b78519a0ffdecd0b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h963560075e453acaa98f5cf69a64363443fbf53a8e6ff12a6ba4e51137b1857;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h79caf2bb47004b1102693381724425540e02794af8148ee58d03c69603f87ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h555b6fbfa212a5a248beb7b3a9e40ae7a52aa7a909d420ecd542f8967085506e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf8894c88d05786682ee9f3e571f0616c8a44afe8d2af96f3fbcd9a1b4097a96d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h851b8b84965b83df3cf684488f89890e451585dc7c64cb592c9ce1b9f1a0f4c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2fcb038a6a5705986188eaf2b04d9a4774093a975d8c40e5dfae5b7fa707ed8c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41d440af110ed60d0e711b938dc8d98d3e9c6647ea7c7215813897aaa7df5213;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h889002b9aac2ab20a4e8aec78ffb449946b0717769d1407e15d04a79fdce8bc6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffd06abccc36c9414efb91ccea4835c64be8c393bd5dc03f5b988219cc951f58;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45d35c67dd780657f8d0d56c9e89b1d5d8af47804e5089df4e958f80fb955370;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85bcab5f78702428b7108c6d76d82d6d3a49e76f79d34a36802c7feacc8e1a30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfbb13e9a038948c69725f1210f3952db25513a853f96b85687c14216d6d6c0c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb907af92902bd59e18b9cfa3a6e74a265e0629decb1d98fe08d761eb6a940477;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5755aecf56fd05a5ee8f84de58635c5a5fc8e24aa6eaab9d3373d9e8957563d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23903a72a9ee265a66404b78c516087cf10314290fae4d12518f079f35e57526;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44170376b8f2e814da31f9b8b0c00df2e1851e05eda668a7419fe17f13bb56c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28303c50ee4976f231c402a29a84ba64cead422241eddbb31883d35a3adaa872;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8b74355403c77f257f5a3083ee13da17cfd0e1f468121273d2e70679c6f60c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68fb238016a9b5d0d914231708849ee7b4eab54c5afcc747c342f4e9a71f92b3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5046893179c1b85422b8cf0cfe4186da004b4e08042c38715daf9366e7d08ae5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6177d44291cb64be359282aa23617db4107ab2005ebe57e84f0f8c3e849d8bde;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6a539cbfe3786c05481c60141172f3369e0a377c42e02b89167b7f765788c1d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h803490b72afdf54dd370acbf44626fdefca1f1a2051c1c3c1eef201e71f8ed44;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6152b14f838bb89ea222d90d23cc918f4bd7c79e4dd028716d7c374dd5af1e82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h960c557167c7ba53601b66d503e0c9eace973105c6ac7914ac7d7606f333a045;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36da0ddd487b2bf8141cc037a78b6efb1425acceff122b6e5cfe577c47a444d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcac4f140c7ef8eed31e000ddc7bd9d07aced7b385133a80c4d76055f702caee3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb931e00b119ba0aa2c1572b56f834bceb58363022b8475c993726b0f309ee843;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb79d21823c5ef9791fcbe8ba1d4b089044608ed3a88f188a83763ca1180d569c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93081ed2a20013cc5a4fb52a70ec405f23eab4d0dbaafa8f4efd16ce4ac39293;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h865179014c3184b749851c069223b273c8cf30b89f404d612c93ff550d874ef0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3225ee21dfe18425d2c0a810e8838b7b5d0ba1920ecaeb368d697070602e168;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd57deef4d61ba637f0bad6119e745d97d7c1ac3c5b0b1d6814b15e875a4c17e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb729d70d762a7098c1fdb5d3c865a2bc7991a1d5e68e827b390d5bb82962b0d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35a50cab40f2418df785cee54b188fd0534537625b6087d21722e7413f647184;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee7908b2d4753503b0b9f591ce37191b9854cb383e982ae7425686dde9ef89bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h713a1e518e1b76c59ebf42cdb8015d4524926c0283d93ffac6ff515ae6b8c0b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68fbc5d6291ceb5e10baf4504ef4273d547a2cd999bfa95b07baecd66fbfe56c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he921e2fd8fa9c3545218c0be7a36d2e4c2525d0ae48808430b3f72e7b47d40a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32e20061ab5a47ce3fe369804e69d55208526cb36fe59a589457f3265ccd6d98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h656e605e1e4bb30a506e74bc8bf51efd60ff206a30617b7f9364e7019f32a700;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e6be60af11760cd2ce32d1ea9faed4afce758c70472cedea58ec301af8e0d1e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8626b32fc2660a3e368c9e32c64e3b68a810645f7ae000a501ea436f19344bd6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53d66d592a2b1f28163fe1328539d724fba2752c11a45d20735ae476746483b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5fc7acb0e946c823b1a89f2282b87229fcd8bb1a4c8fcb0ff141cba82bc47d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58cafd85b507dc9c8557289c183f5a69eb581c795e9e5c4c68bfc8085681ba3f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h241341a955d278cc5f3d37840d474998a24f08dbe82c0e79110581d8a91d3cad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0bd37fbdbea8dfe3f1b54eccae54c397b74be630e369b8c306cb2e48e76f9d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5da3205e8dcd8325de8ba88c6f3d3c0e02714340c9d17e79d363144d2283bf6a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5f6a855ce0115f225f42a06c2bb1fe9f524c690f35acae3441298a62ccaca9a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42d8b3e60c590e12d602faa7347930114fd3595aba9fb7bb49d5a9892a4dc57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d530eff3671ab353f99eb73cd403fdf0e24693687c9fbca912db059239b0942;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h813b9189e7f0c0c0927eb9c340a986836968ee0f0db60775efda6de767716bdb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h13e64e1c4ad0b176507b95c7d349a1ab7e4c1d79497bcf61dd7e4abfac40282c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8852d2c1a4b1fe8c554bbbdd7ce0f77e9dca2e69202ea999beede3c88ef55506;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed254346f7eb852dff7d099ad100ef7e0583a55ee2314b82bd93d663785a1f6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf90f73ca4f0c951decebd6eca32fa3a2571360de96e855e9067c4220687efb99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf02deed1cf07f35492ede4b91fa59a0a97cd9aa4dbbbb4340e6911dcd0455d0b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcae0d696b4e6846d63bf506e317ce866c786f95b4b3fea07fe98e41d4cea0b1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b028ab117728210554af438f54e04c5b0fef1c3b99e60acc4d142113684ceb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h27ffe8dd0d0783ffb9fa8b01a348e979dcf646548fea7b9f488bdf10bc136527;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39ce6f10b65b77d2665dd8dee8bea315d5aefdff1cc713f3b7db8a1f3da4c7e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92597a3dabc940322c235759329ac4021aaa9cb6bc9122832d54a09c2a943fa2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h713909201bda3376ce9189daded9fd473d3ab780c9d1086161886caf50e68d24;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6294438d23b588b3bb2fe381ad8692bd5d39b6a243740d12adce63423b7c30e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ea0ad47ff0d1843293f77275fda3f1c602a650931ca2563e6b93d2b3b42d117;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h926ffcf46c06036787629232ad973609d90a62359fbcd6bbf2330e940b44b270;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h133e964b0f04eaf23d5f7f71d1f29113c03afe20f6f0b8bb0fb7387c2c9cb901;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8187f529f5b72fd2d4a7618b6af80b4447523a648542cb49dbe6ddd65aec476;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e88c51334e4f386f512295b57b63b614136cd182caefe29f7bc41a1d9e9d8c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc61fae30aa81dfe891dfe79f4283abb9d9e9390869a89804ac3fb16a61a4391b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15ac051c14c101d0750102e3ce7dc6d0df98c9cc71cc839f81a2e4c3d2aa36e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46dc5c112eef7948b070ff69751688b8fc75d4e77256c8bb21d89efc89f28082;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49e07847118abc1ab77bbe5be37a590b847aab404b9fff384a781833b70d98be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd70227db2bd492409ce8d68eb86cf23c90f2a51209cf9daab29789875c4cf516;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54132f49d023a2d8bffb33e4165abd8836531649f0520701ea94e0c79679a216;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53b51373220ebf7449c79a350138c3c98306ec8b565827d092fa5a389f494d2a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f488d7322e4b4404a09820f0a5216916713329e16a37bde4f6343ca5c812a94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha66eb829402aa6e0bc5d2e370db3e80e5107052853dd6f1f24a4c70ddbb4fe20;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39f9b33a9c23b21f21bc05282064a8a92d837b2a1ee121d4f1696f39e031de4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h201b79af1d801f93a5c1602c781dea4aed13f160795a561c300db140db6adaa6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90dfe159bd00af304852550edbb9f81aed1cafc38a4304f51f6fcda4b4a69bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1028ff5288298eb24a3b9f484937f35f6409122baebd4fdee09cfdc77e4f973;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc20f5618e0d798b569f35bb721e20599d55601a5905bf2802d4567a91371efa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h828e96e7d99a385b24d1532bdcfab3e956b9094755cd52bdc32477c38893cdd5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3aaaced60af68936c36c55902bfa6c9a32d1882e303de5b2ed6d2d4b683afde6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h494ee7eea95b8af52890fd4c5531a4f3a1a000d0995d8dbefda8fa594abdade3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5d5cb8de1fcbfc921617ee33e9fb4229fa3011454e8a8938f20acb8472a0533;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57ebe30027e4e8db35ea073ae130afe834634f1db382d23b931f5014532ca329;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d28691c0d817cc88bffb095f035f7d448542ae731a16582cdb8e04cd10b7af6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23e9cd100aefb42128d568a897c7cca41b5cbd43360ec661be64b574e825b080;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b58242635e7c2a223e14956bf5c44328ecddde306b490a57e47ccff3ec73b3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he43beaa5320f15ded570fdb441c6190826ad53653269ec04071cf3f4867ce009;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff079d2ecc85a5655e48f5443eb5f87ff7c788758b323b1995901643d25fd4ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8fb6b78af1769fc92745c204f0c0beb6a5516e76158328c7dd4d54562547d7f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h796ab61cd81755d3c1cfae0ef98f2eecabdf3c9711b4308ec0e01a5a566d6d0a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbaa1cbdd8ef9d00d06ca347809c3a12dc5f8915cd799e41825147ecc05f16d5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11b8554649c2cd618563edb317c98bd03c8af10f0ae06c643f114aa4017878bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3261ea62a1af902814aaf865054fdbae77a9a01f48baf58e67cc8039342809a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b3a59135a7f98a665a3d22dea802eec922ba995efb65f1bc960ef6804786f0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4851437061ded2293df86a95b37384b477f6d78c241a46191964cefacc3128b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d941efc8a0af4cdd00ea4a1667875914895a30edfb608d3c20acb087532424f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf604597e3c2c636f38e49c0665f17ec640e2cf99604dae651f7a952564f75a2b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7cd649704b0617c10d12dfb45032b27c32a41a1bc02ea85625042fd71c9bdee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h973c03ec3c935b80a6c6616e8e6e5480be315b5d8f6d4244ac7381c5f3420c68;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe3dfbeb9b739bae5a558fec25eeec20d960efb02efb0ca7d3ff5dcf3c135649;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b4dabde49adb08b20ecc9fcf3842dbea0092113418351ca64b109c5011c15a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4bd4f53493fc55765b85e8faa412df851865442a556e14e479ab58e61fb3999;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfcaa88f0f0d579a0344d86d3a866973f0d393bbd7cc1f66e2849f667f0905ae3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h592f19658c0b23606cee235f20956910477f6186e48feaae496296a6f9d651bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6bd2fc548910f5aee7daca81cc01bf1c43d16f63212510c5be8c30cc7f5b4f9a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h651a63fb2f6a5a40d8ebb91264538759956f3ddedc87de16ddbbad9c6bd52c83;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b10043559e536bc5d2a82c7648180ccb4ecde509622b2df0b9b0de6d008584;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46e042f29bc92464ba204cf82287d1e887a5f1c5aaa69ebce9ef85fb1d79db3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2121e6d042d8cc7237a57e82f4ab624852caf8975a40e06eadcdd4aaa27ccc9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6f7947ae5f12ff9d4d8ea4f8ed7b199783ec8b552095c9c9aeffeae89d826698;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4622fa93c1b591e701abcd3e4b6ec3594ac4d90ecca721da762d53d93b5102a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf1e43db4200a8e29f4d71f5d4afd9c53295abd0b654d9cee0726d80d292adc8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h581c49672c9d42e8a0284c1dce60ba5edf8949fbf22579d0c361555436d3eff5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf485ca30913f3cd6c9b42a57a87248f2a97c672b4c0ee295f804ed4c2f71f4cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50d743ef53145be4a42506f79bec92087278dfbe98d5577f5ee46448ea032a21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd113147b519a48db8323fbbfabbfdd0430e7b9954d80a9bf460ccfec57e5f236;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5b3744d811b20d629f69961eab3c4b0f25c7f68c50a4b14c8a138c7cde81e48;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf68a1342fc213ea77a6992a8a7ea781fb546c698aae2d1013e1dfef2ad417281;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77f8911e00f4fcc289c91eae63392eab93886aecb58c0c50bf519b73a0cc0b4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7cd045f44fd85bb378e1929aea2f3a67ae46923e097e39ce6b21c8e21e6e549;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hddec461df39158388423409c92974264e881f15ee432f9c6a111e5992dabd5c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h590d8afaf99af6e6f584162144a400697eacbdea0a1e5265a41e64981e43f39;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h289edceff4bd6f063eb4073df6dc0fe64de9b25752787b3f0177f647d3844c67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72e7efc929f27295d79e258b623c5580b2f148f1fe09a226953d516720837c41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68fa3481458a43490786f60a9ba386401325958b46e06bb0443aab6efb4de020;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42b51edfbd3402651f8af4234a3b17e13fdb11fe81ff88a4c710ee087b904fd8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ed613f8e141c9fd6f0b578bd8a23b3d6c7cf396efd0f2d4c6cb812b39c171b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1dfd2f8b6f480c22d9a104425c62fc0dd941e9878f7c51c38cb83475045bb33;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h680b4e386368a13c0179a0cd0c739e9011b045e605b18169038856e18b49b557;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce46453f58156d0991e6eed5f822c36353df905bd4ae9892b4210807ed534f71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd740a9abf5833342c618248a7740a91fa88ac9e1bd1bfdec91bd06a34f452ea1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h43ed5e0539b7d0f4e7148a0029a6dcc4fb37650b482c4d194ff0f9626b3f9bc8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54131028dfca593f07a0c1e1352cd5832793380399691b77a8490a97d3ad6220;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7caa6161251f651927a6703f621642955af97949c0e8003500e8bcd7ed5f0ab9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80db99c3b740905a9cd016ad4a3fda88dd0a1d00b3111056a160bd52554f901;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h735cb1e46aaf0932d93f2c0c5034f0351b51def24da6f510eed7bb1e4106fcdd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7a60d1be6342f2b8338c98cb49ec5d9d9dd1769c45c8e2d08ec6feaa34b57bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6a10f5a813aa8370614f936b1e224dd0138ee97f8cb7732c5f82228c6e9052b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19caa97515f2018066b653a62d2d0646bb671dfd73e5bc997e4882cb8576be1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha74e62d5a1118fe6b99337771b41cd8630af520a6887aafcd52b150c3e77a0ad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf17762b0e5678a696e6ed14d5bc155919e072ac401f84bde72727fbd33cb05b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37099bb678201d0a95f6fac8631e57d0c479164a5f1a9b1cb9834d9a208d4e2d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb381e9062469004fa21935c75f0c3a1ca88ddc3b4507a778d9a2118a492dc64;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7314247891613e770f16031a4e85334d35faf916c7c969e7372a1541895ac56;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac59e3e884b41bc5ef05669aed47e9a40d6f28f8843c3e3ab7c55251fc84896;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e18857b43475a98e8dc80e7ea55cf84ad0aab559437a6310b50c0db0805664f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24ebb1265566b36d6da6baeb701aae203283011d71987ad862366914755affc4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4304b292335e0f38703da16ab0d015ff41920bd2a48eeafd25a151e0e012a59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c4b7dfa007ddd1f302e43746659c5465823762872c31ec97d4b4d054c556af3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h853424035fbea7bac96b03624d7ab998544500d118fc6316b762ed17f939c420;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1edc95496abb99f2221c09be06df745b858f929eb1954b102536fa20a0f86553;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0fb9ae6faf37d331f041442214a4d1d9d0956957c7876103cb7344dedd0a04e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h636c6e6e2f9052e70d8319c7fff2c714173e11a688e94edf420a768144f8eb65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfef4e9b5944040c08b2b19e10fe29573e6bb8b49704758aa956e15522ab43cd6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64e06d2ba681d83a73445ac67f95b564893e69cf3d28a01300ac6e65a8da1fb9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92b20002c529b59aff25d4d519565192f63cddc5e8c31900144569c6f48cb60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78f0185b9440f34722f621aaa44adf232468e66a91b6c65b72afa337ec5a6d61;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb517dc9c0d3fea0dcf58787aec211f29e96004131117e41e5a2d0818d9cd6db4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf659ec81c1d93440c398a2240f2e7b72ff54a369e88330344c3e4a5e571ae58d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd3cbcbb9459b700e1b9e50dd47e4e3fd0ecdee0c6cc9ca940a45f9dde85d6f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbbed5e0e2a5c4e018b851e31bb4825a6f6a39c9e3b7702ab0f86071aa8aab297;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha084a4e2743c862d3a1a6eeb5c3b577bd07c5b592b231e3169f3fa67cca781c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h196b5a67e0aad0cc8ed4325dc3086243e391e97b3a100988e65108dbb03ba5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf14931c37de32b177fa375495af2ad7920d41354f976c96a7931642d8136e492;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6dc4d9d37334b4bcd74546cacb7a7eb1c0cacc573e97079e4850083c08d77c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8395c35946093c9ac843352796bc210325d61bf30eee68ac4366d9f7c8bb7fb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h183f692603fae09f2d915d7dafaf121442aa5291f0c5df95f26d6bcae0b71818;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3ccd6c00034f09840d54b07a0eec80027fb6637a7e218d42d2c159285844925;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50cb4a5b35e40fb5c4e7df944df41dafbcde49cef0318656bc1bf22c841ebe49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15dce32725dd310ac138b66288e547bce49620046cfa24b5c22eecacf5bec6c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5599cd52005f50d19f92307d6053ac787e92b9e59168fb0bf511ccecae91bd33;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1fa83e4ad8ed85a459d84c8d59fbd43d7003cdc5cd19746d5aa847a403c6aa5c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2340c339c21498f8c7e569763dd0fc1adb586797381d268f760930be3f0d4e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h13b1142179d2aef75b6e7279d2317e3d1e06df33741ae7e1ef04224409726;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7915bc39183ddef8a6c6f3a27dd48663dbe79ce5d3b7ad2f886216862eb8535;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19b2ee7f08db2e77d5a9aa29333fd63858446c7e32bf602ef2bc356d84a0c445;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72c584799f0cb0f718b9ccdc523da1301657a40ed249f25efc0b4fc8c0ad2881;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a53840c97dca2787a7c41ad987e6720c2706539cd401561023db33a0727305d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfdd7dd4ae0586c29f6a731f887d881771ac1b3126ed203e15a7ed90fe340df8d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6a7f952bb438faf98c3815c3cb115e19781afee53aa01f1612c958a74484b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hedbc525eca288356fd6d0ff61e85bea1bf97efa1c6a0b5a3a1df957749066e45;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc8b2ab606d7cf0db1e47307ba26431efd358d4e5a060d54262dd85242a9a7dc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39d2c15937893b004c67e713b89d64ab8668ed44b530d7f78b32d2a6a5d55ac8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65807aaa1daf4cadea6ddf29fbda78f20e8b88915ad92596297f676247852a86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5dcb32fd74f87e1e142b258c4029f91109a703bb70457270150213a6e76691;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2b442133e5928ba3c417d461e4bd1f59264d230ddf78dd3cf7ecd4fc2a62f97;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32d5cf856af008393fb7dbeb613bcee012b9c7f41844533d3b701c40906fe2c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he74a780f9065cd2e40d1d4b6f6e2db0cd3a00ba43ec92dc466f3ad6068083c75;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1167c86ec09e5996d22a30733b7e4b7fed1106e861755f266d74d47d59a9170b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4920a656db696c2ad4e7a84239118feb0749f113e48fc04a9c5fc8d60ccebb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h397ffdc528c8ae58c45ad2a4041172769aaccdf687dd8dcffec1d658ccda0752;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8271b0673ed5f4b81a00cb41e72d899ec705f73f499c04ee833f7bd588f2c80;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h533c6aae51de9b6509fbee73d6a608850d91e50d433f8b8c42b5c773ebbae6d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haeaaa012c7cd73d55993f4dbe2e76b8e5e25a9910fc067be2f02d788f83e3373;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c3c684c1a022666899f3d6254a00e3edf8e24aedd56e907dd3b7bb80e7eeae2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha02fe0394c52e5af88abcca297514d2b87f8d398910d3853a6d400bf4d431fa9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8dd4e0760997fd40dee76185d1b3eb3a4336b1c81ef509f524d26310871d7284;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b5ff9505484e5c3c67ff51f131c63a0d750b4174d9e77d9a4d9757ef1703c01;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h731981850a203ad8be267e8aba21b2875e852d1a6347b2ea2d7f7d556b1b18d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ad1eb40b8ea78aa4c14a1b3fc985377a9d74e8b75471db23d39782744b0d487;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f460c62f16df93b4dc5f4fcf5667916f8842a0b7b8d988710c173dbab139b0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5af84a24e51800990da819024785ddfa1546ee4e54873b8fe58bb38c62fda;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77711ceeea16f99bf1e2cae69353588f17db4a335569a479e12391ef02b76679;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc1757c3aa63a2114da037a96e2d708255f9a05ee8462b011a31d38cae54f217;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b77d1065e41443482bd35987f45538bf8067f3a7bf2d209b16ed0689fe71e20;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73fa4c774bbf1f86dae093dcc05320e770241562c97315aa8e6db1cdbbfe560c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee7d5c1e73a6125e15ae1dcc77a60dbd3cdf0c1409750d0841626dec5cc18c2a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h255f27c511794393dacc5b03c8735556aadb74f63abeaf65c19e2d573932b99f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc513a30bd194bf7d5d5d5f91aaad7dfdefc99894d9962efe83d65ef4bf37b61f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ec82b197968db734c219ffafc1ef995da32b20e41f7974da65f429108c99963;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfaabce70627f299fc8dc06a92ee3029a0069154c4735f721bae2a6bbb7c719cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff1be7889f5cfdc16d67f69ab7a87444d81e502d80b15488656fb7b2aa233551;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36b6c8c067fd3d4b4bf2b936e1da744d3f141b1c2161d3221d61fffe59f3e883;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h994ba8a3788d112713d9698db3516fd92ccf8c5f924bcbeb4b8386872d36fda;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e511154ebcca6ba60b8227a55e2ce78a25bd54a2e3732818deb58775f08efa9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a0617635d22fb4d38370e230f9aaa2367c461faedb187f635b9d242e28bd92;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4aefca5b03f88bd27e1e334bb3768758ef7e5c73175cdc093cfbe3fb0da9a3a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe2e2bd989b797d44166e844a709a9968238b3bf853901cb7fb14b5bf948b4c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdfd5f84f34dcb9976d99a473a0e41852e01212223ff3205d22541886d36a0897;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf7fc01683cce064acd5839157ceb9a88b38e89e9bcc827fc5c229d02b1aeff8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa90ac6a54019942d489467699017e0d36d74923b69a9b4e31d713f6f59c0fcf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h353734ef2b91014076d9797382d0aa3a41283b4120c21107bd5ea24e7c0b393b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6ed7f5cd8dec4e0dd3de9f1d87151729de7c5d4730b745d1f90db6df2de256e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he87ec8a662895e40eaa1915adca263d00ccbc94d1c46602914f01e5725b0b292;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f489a5637aba31b9b3ec27f441028687387fae52e9240f6aae36e8f59da2ad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d09f442cd39d1bb2772f039b32e10167fa572acc785087dfdd545187208a31d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5a036ba2b5583e6fa59ece856ead7f7af719c759f3441a4c0b872a474de17a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37dfa73701713b824bb5f4c2cc8e7b4386293f83702f76a42ae7f83f562ae29c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdbcb3564a330d3068f9217c461f689d7c5aa67171e372daa33251d6c42e4dc9d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4b93079789af8a0093c90255ae30412df26d19f36dc9dd2d2036dc9d40682ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h501989f967907f7817655b78515f7de64c6390aa8b616198fed07f7d70a5379;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbde2d87b5ccf11955b6b26956bb33edaa36390c33f86a1f62b6c4ef2f74e86c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8383b73012d3471b4a068b8a4b59c5fa1608db41e9a5ad5a8e9d6b907a6e681;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hecce2d9eff9c2683d564fb21f2951a0b525af768a074b9cc2798ea44d953946e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h50f22eebf46e18f8e4e752e580b34739ef61d6d2eb3aba2c82f6917acc05f405;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2977459f5f9097a857ade0b77447a71023955afb8d92065163b3423f83a5c743;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4cdd95f221e78679d2909f7ff5a22852e7ece851a83c49be2174869eb8d89b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d31efb693a0a8682a1db5abda053b0556a4829f58ea5313c14a061bb6009569;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3fde22a2fe971a813a7ae35f7f147f49964bdb751aba8170f16f466b6d523e0b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba5302a22c8985974b6ba8d9a9e9d445a0c8ea4f95b1ffe031c301d06a679295;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h81d735d4164a5a93a8531fc86e6aca6eb274f20cce71a5e34dac979c4c939944;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a30819f4041540b27989e55477677387211cc8b12c70eab94c3fe3fc9b98d7a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc1c19b0ba6397383fa50f685ef7553003e7e7bd16af9b97586e4745e807b74b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d02812e160464e0d3b4b7638968ca565c519c09a0669dea3c2e72857a5c7a55;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb2402c9bf9a3f1b15ae45e9b01f301f5d15f58e13c162ea43bb03dc7db355b88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc913a16e7b0b0c6d0951e44d13a34d6f1c33f5ba6956a6bbe45da59f8e21c344;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf584103e2d0390e914faae07cee3d5c361927676e58a1932f2db36e0016a2a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hded89ec40c822f6094ea49073ecb8ed8296fa242503c9bcd5cdd453addef2b63;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28c2c2bba964b015c136e4762ed77322b951417c6ba0de1a952bbb410728349d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcbbfa46db3b014d030ab7220b3d0edd907de0750fdb926e806edf53adf28036c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc003d469e3f613d573318741dd08bce5c36916c78a8c19ad51cc7d5f058fab53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc4dee7a596755cca4708db30dfcf920e70977ff6324189ccd69bd2868677355;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffc144e9d5fdcefc7a9f4963648da504aac23ebe17d05efda2f7ebdc0dfa1b2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6056b2fb7de02d887e71c6957dddcc3d1738d9d503ef8b5066c2adba0ebd4c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h180308611ec7477c9a6fe4e6835ffe0a84d6121d45ec397238fa807fee39356a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h294f5c69ab2ee162c508eb7a5b8aa6991e78e619c0099d3278323ff8136578ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h353587b0b40513f67fa25e0177f3589bccf5bb5b8df41694bf04cfb141c5ac2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8edaed2e863d870f394661d24b2de3b35562376271cc61a6b32b9849b2f15b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4880547cce3629d9f828bfa4082d9281686d42a1fe0476942a13276d7c5171ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4850a690147d63486a3b7a07def6e2daa5b2fbec44453f99a1cde73c844b62bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b61e11e3a119ff333f13e7984dbf218b7d0cc1bca816967eba7b392cbcecce5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h761ff49961392d0b8ae66e54a3a976eb155ddd9ac60542aefa82b4cda988c34a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfba720d7afbb74ecdb705910c032e25f415a207f9aeba8d4818b955cad5f1c8b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b4e1bdc9b046162727d7d1932d17a0c5a18331d694d949799c814209f362b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heeb2769d70cb3444d12a8fe6250c255dd698c6ece45d109b0beb1409b9a77f5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h237690fbd4dcb612c6143b1a5f55378f562158d07e6607d1c317b257dde04dff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52345d3d40652be1404b8d31648489d7e6fb0f37c2da4041e7f35a6d503bffd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d9de69829abebe6540ca9bfa521def3454ca0bbb1359a5ea2814f582a316b5d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h556dfffcb53538f5732a967bb97443561133fab17de3d00b23cb24292b0b9eb9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8780f04192d4604ec07670f08cccf46155c3ae193df120aa6aa62bf0e0c97ff9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3d0f3d3c4f0cc52e42d47041086803a2775aa72154608e002c6ff5bd4d3f92e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd6067dc5fea7898ca2f4690bbb73011955725696309c3097a04cefad75b6265;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a5ef9411291c6477cd754c314cd0b42368ff5a243cad433e0a9d2d9ec7cce20;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89bb85ee4ede5f65624864f1be04d815b88a05585942a9d828fc2d8792d74808;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h18c467b9c8cd0fd04dc5b7bb1ecb51df187c49ef6d3e9653b0a865d738325fac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7001db51f2065256903dc3a3f8385ac12e7921f395ffc5d7f3d53089747b8664;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc812270f464831dc717004d2352d97e7e9fa74e513a95ef4ded37104d7fccb57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4f47f5616e382c62adc353afafd3f9c9ac96f6567a0be9b1b60f633b269e20;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he877347d78149ed6ad905c3abaa8c03f28efea9b96bf5b1fde30d2078d6fc1c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha10d6812f9c418f7b987edd0e8b2b20d4c0c64da7d04b121362d0f3c7be2d810;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a35124e2a47875cdfec4b8e9ee1c74ae63fe92cdba91c6aeabd5679e93ff1d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5217527cd11200b9bffc91ad0b1738faebb2d018540d898f305344a0b948dffd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb626318057c127958aedc232ebe090aff444912f5643988f5779db2b093b5272;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ba81882d0b9065c7295b173c09958b680070e61f1997aaa1f4cad490c045b49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89c1e563a0302788afdc5b14cd4cf1bcecbc1eb7454841aeeee1a32149004ae0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5d28969a03425b7b8fe81989a317809d1a4b1f878f8ccf18dd0118cc336854e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h81e830e58c6dc4c2d7869e5b5c83d5ed0293f1ea4958154402f8ccb58a283a7a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h805cbf0fe90885fed268c344c9ba453b3d636f1cbb718b00d1dd5e0db6203ed4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9966264188d2b9a4941d35758e57eda949a23feb002fa2fd1638da67fe7dfc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfbad2cb217ef2efafb8b096b2029b303cca10d1b3af1a98df3d2f2aa58524f79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4bddba7d33bf85308734f35f422e28981bc1036e1effc4c8759c72763a5cf2a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45a1593fedcd4bc13291986d47ecd13b5896a234cf344dca92749bc68ad30690;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h14c93200bc5b4a6960ac7872fc3f8bcdbbb27eaa9a723e902c43e70dcdc42001;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8535dcb9f9eb8267d1777ba1954dc4456cd03f51eef37db16a39f4ceeb41227c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha428afe1270328accd5e95167dbf4881109e838d7a6eac6f2fdbe8a69511fe07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87fdad49a26d069b638ebead7d4a18f2d133a26870a3e8760b35505e88ef4f44;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd9fcde38d95bada88a9a589438ce741358c2bc84fe963afdc783526443224911;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb8b0a8a824c1a10beb89bc4e2af5d1f234bce74016a14456099ec0371453483;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58068b4175c6dfca0fd18773628b724fd673fc0b2da1336f421ec7c79e544430;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha192aff28a524bd320ac15756934298ad7194aaff247a7df29f5e09209a88705;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf09e8d00e9616dc393a6c98ad543378c251df9962349a7934d620b52abc4b818;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he497e1c1e5474c810225d1332221251ac803e4be7904e219a8830ed32b032f3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h571a296b3ac870a1f6816ef2f2a23ef20bcbf4266be5f36b3d3f997bb623f430;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heaff60dd33a94c6c45249828bf0d4d7a62441fc10b24944c04f2ce08ec417e40;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha861664db206a71698a56ee930fa85d17baaa3c756cb0b0ad9bc0a379ad6f229;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52e5e94ebc5a674c7c4e84cf6ece669ef57307b46e5a67cd12c0a456cbf12a1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h289bef94881762628adb14c0cab276860dd49cffcef6e50e6f0a76d4324d9bad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he730e4c581fa360d47158ffe5f159b5a1f9a317063fe230cee764d27a0342b7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h22c592a38cd3f8898356bc145e3e6fcc9593b2d54912f2c3556f772f11904d8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3154504e6a55243de229ed1341d4480f2f1aaeab2aea5a8a4c0745070b595c37;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf06834c4926d4dbe825e92dccb550f465f8d98e946ff0cdd884545d6334a1a05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7aeb104ec30209016d36706a1a1c2521afd5f734b008ce3a51f912db29158dea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7fa201318c6e0bb0116d319865df310f2a7abfb65af099fc753d7c8f7787b85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf41acbaed8cdfc5f1f718a9340d585f474f4b2dd7c81bb97aa1d0efdb6fb209;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ad1c81a05142edf7710bc1ee39836c60925c47af338b54280d1c6a82fa60a3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea18ac7942cc95b09fb14186d58ce454e5ce633d619703135c764a71c054876b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb87b0ae748ee1cd2e276506109130eb80881418f0e301da862c571320a3845d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9557737da26a5ea8cb07831077220d1ee74fbe36ab9a646d7ac56abe1bf972;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h348b4a44fff3ed699b48048c6d936c3119bff6a9b1cd799ff0db47ca6dced344;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heccb85a12c7e574523900f50259c28a56fc17425e380882c6f75904d83d43bdd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd223b6c4bc91104885a0e3a44d1b061fe7b9aa2d1dd4862589440a4a8825ef79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97e36139897aa78745059c303a2330aa92461160ba12c4212176d6e58fd10e46;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf434d1c9620cb0dfd9a23a224095d255f586f8eb97734b45f4af8c5f7f150d59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5b293ab97195e3642442884e62a6cfc6e4ac41d6f0f4f9fa96f20d00c5287c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had539bf7263a97ec42d37fac954478b166ef6db1932023d861fad3426b1b05b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d5f448bed94d12b183a76138535adc2019bb5b2d8eef6739f35d0fb73be7a3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h487c7257bc834a0463aadd674a66dfaf8fc33b20ca4bbbddfd8b6605c7d90597;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7bd83048c09ab591e3b08c1565c099965f54ef19bf39b0dd3f9a8fea3d77a63;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h755866a81b6e589bd64d58a14ee984f546020938ced97c3ed6fb65de20dcd66d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9fd5534505778ab68f072e17cc08352fa746577c134070d5c9e4c98e2a7ac06;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h931549355118a81939f133408aba7f0cebd4fad67d747f7bf24e620b98e6813a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h315083dc7acd55f3acb665127a39eda0c9d624399eb1767f6df01e9cca13760e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7293bdde7b2348f606bbcda6253c116d1cb3137ca3d68b00f81202ace0bfc4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfd45831dbc5a3892551cd590e036a06ab986a64cbde82f73fcfd408508e856fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72670a6da4682b390572206e78eba8ddf3bf2a636b87cabd85f189ffb8c10009;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h29a1ed2872615e4ac11440c43fd865a6ba669bed6d76d6f2bc5308152cce765e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80637d466afb2a87a8d5fc298458f0eaf40202cd65f730d5e248273d7acabe69;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4d8aa4d719a3ead21f1f2897001a464e26ebbbf2e1de22e898deffb98f72bc2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf114deadf42fa39a25612ee990874674d8c8c3c171c32e5cec727620e0167cfc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c0c98037a92940055dba51e94255370f1417032213e345136de96d5988c517e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h839e06bf24f60550f506c940641ada240ce2d42ae818f69857b93397c8475b9e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ef017ba18eb8a90599bdf811c0c29b7affab3e139be0d10305f92d94373dceb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7aa6725d67b4af4f0c7052f158b9b1acbac8b10638fd54989b2ce57048870bd2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ef8fe9a0d653c6c97551fd59b2d590ee8929cd29b0673908836ddd5f27c654;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ed512a5f9fc60cad90d733301afc0f91372cda1d6ea5e4e0e60dbf04f6af495;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h913640da00ebf3e82a6d8bef98b4863b5bc6790d4b3cafc51e93187d7651a93a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbfe2ca8f8efb867801ba4d7a7d59d6aa219b3b84e4be992421b11c0f8d7d3e17;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he080470ccc50566604ff3815256d772131eda1be72eb46fdf1c2ea5e04ff04c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee6ae27a8f326f3fdd02c9e48e483464a25eda4e343560e3934cb84c54c91d1d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c5509c9d985c00d250500f03534e2806db60eb3b3fdd66d89f1ec75c10009a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1cf393a98ca23c899ee149bb03808d12858de3ebbb4283eacc1b24c5eb753240;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6128a7c9b891fc1fcbc58a25c632741551ca5fd5699f3df8275022ef9dc75a21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha78f20272da10eb76155bb77a6b47a0188382a0e5461fc98df06a66a3ddee3de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d4591ba89aaad05b37d8c2b2b32305d3921b63595a4cf44986676c5eb282bc4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3ad5d65a8fe47e542c0407803f1ef14c48bbff7161bee495ef7ff9c27a6dd0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee6c7409bf3359c68c3516b574566da43c825dd878a7323286a2150daa985b95;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbdbf7d9c1ca115bc154045e34b55edaf6dc6abf3f4b15409922b39624a2d0f01;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a7ca60eb79145a3ff6d4c6cf5c1854c8b1775710c0797cf2b0897af4c130506;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h752d9719bc49a33b9c582059adb18f314cd604da44bcecc505d428e406756371;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3aec3b73568dea886f8129945ce14108e40d9b19705589905947fc029922fb49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17f9a5b260c426f54a1dd7e4fcbfe1765779ff998a078a1bc942e554d9763ca6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65189c17d0f1e73e743b2780f9bd1a6fa7790926055729cc297b5cda77f6d70d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4949e4ebb40a3d1abdffc30955d7553c8b3cd1a48bcca55fda11566a39f7d596;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5924b9cd0a317871af6068d64a0e3aa4cd124736e0b5d57a9ec0ee6412747b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12b31e0024a95c4b812de0af17a23f81f0c43f6c310babcd69a52b962275e84d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa432cb094a23f47c33a648dc0e07ddf044af9b2a1b3a18a262daa2c3831844d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10d5dd44b06b1a8a3a7a6e7392c4d654a5c24ed4691b7a0e733b9882755f433a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb96874ee3e46130087b699a85dceb0332b7715caeacf250eaf6767215c17c5e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54aec07413d24b962251ddbfdc48fd7ba1e97eb2337407b316e1f7434a6e7f33;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf72d1420e624eec97b2f932dcc4f139c818bffa9a37d4bd3b6a82b9300cc45fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb71ec471d46970426bf2a3ff1bf2181b3b43098d80dcb3f34a4e34ac3f9368c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5ee9564f8633aad1404d5e971961aa22878e0c3489116bbc9c6be53094b8c0d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4df7e802f3b92da1f1e8280896799804db97dc3036884676b639cebcc2c0a84;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6cc7e455621223bd71903468c0973683fe7b079c8a17bea77e4013224e757f74;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93712e0431dc4208e2318b814fd7561e70e6f778f3d0c3867f3cff81fa6e647d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0d5c6114396db42654c68fbe9d1bb731e0596921f409ccf687fae5ae0de0c7f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2818a3564218ed9252a63a2e36246f482dbbc83ac859e6abd0655b0ded8d2be5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5b0d9d68990982be3457b8b4b9a102ea1a8db0d6ce7612f9c3fa0e0df399d0b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83317e5e25b915aa22e503697a4cd22ab08be41b048eb55e22da77997ba33939;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd3f32f1d9734f5b598bd22063952b7c21617a6015368b760f75252ba2e861c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h14a385b712e6e7becf24f627c55d05e4c0b6a4591e756fbdc1977052df363bd8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h85f329eb82fde800de5fecb5a586e01f5c50b8f6ef967b1a9ee4cf70795da4e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9de8b73882a362aac028948a4a05f7e18ce52d6b19f21fc602cd22e32b96c2d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ab927b7a0d46eb2876f09832970cdc319622d7c60f6588078e098a033060eba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82f4922680d8bce81e86917ee75f782f14db4d87a1be1745d21faf0d0d412cbb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1bdf91a3e6aa5c67010c482aaec621a38202dd5d5bbe5e9c0794eea44624aa76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac2a46e427c28ba6f76689e3e30ccc250cef0c964112193c3ff05c6f845f17e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25ec7674ccf06873ce5efa41345763622bde68c1373facb38f8e499321e7ecc2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e55891bc1761df9cebc1c70e2ec258998646eb6ec03ee64e3f6d9110004b26;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hedec3eb575e314246844c568b5e07786192b81bc01da84344f8e5e37aba9e205;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdcf192817e393d3460f00e8d5569c7ef6bf81965b2d3128a34690a93a86d2fb8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32f7e31eb355015357b6b0d8eec8c73f353e4fd1714b79ae9b765d3d5219497d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8725aea30361b15ec3457fd1e1f7b48b3e3e405347a02f874623a14701e3e48a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc78724b130c75d2796cc57c010a7ec3b95e8d205cd9a1164d642d4a5641cdaec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h432039f0d135cb95ffc6acb7c4c7e35c5be32d60b2352cf2d3c491ad94d5d223;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc8708e68de0513c255bd66c2463e50963b23ce3c08a0895443fde8f151d65d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he6eee66cbd257ec02f9be02540b56e3514266ed8ab97e1e203c681f80d31082d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3fd2faecb3fe3b1504af8654563a9e67b1b0e4ce7799b9c542368e2bfbaf791;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h565e37fa963cdb9c62b7aea7d2c0bf1a1f703112c0ce61bd52b54eb98805ac4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba5c574b8031658d42c53a1bb2a2a972d1c5ff2e535180723d2cb91326cb54e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfac04054416e1af42309e0f683bc09fb98f44be448deeca2eaa63246b4b7f874;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea7f644fcccde7b73fb3106f67444deaf448ca1414088c8af83e784aeaee8a71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17f81f741a22f149a98f5d16119fa85eb6d6ef032a5bcb5d97019f81c651475a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11e54203020389725e5c367f10adb572b1128d95d5da2f20946c1aa4a5c1928a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6f9b2a11f87624a57a577f5dbc5a954a49001631df77c0a43e18ab8ad68dc59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3febf7f78b594f6db7e833651cab8781e11df9f2540911f766934bd2fe90e433;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2cfdc2776f7caf44a840c629051e0ea030fe9c6f29cdd2ab02ac386908f7195d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb2825df2df596615f79a72357033870876173d11a7a004d7e3680318a83c040;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f8632f218565c45d63f957390c47879b577b8f5f6d7413e4837a1ad71fddec1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80af0c4fdf656a59cc59105444444bf924a650a3701f66e344576df3690df95d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d670abc9f160d0cd2d7c86524496d398ab3ab6a6f869a84cd6ed8f0050fc5b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4578b5b254d262dc5da595a011b5f9df3a1a6fecf42555c96f21340d9e1beb1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hadc1a741fcbd1983ea0588ecac2ccb40716def07385c413d67e991ed0588cae8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd45fd469ab375a10ad098a98945b75a4cc9ac585ff45c72403f6722c27591ae2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6adbb0f2b8dcafa0954311595bafe823a4645e1fae8b880957cf98064400f89;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h764b3821a49fc08bf66fe987a4bc901073672f7bf1314057bbbee66e42c42359;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a07d2322786477ca48b76a168ec182935a48f5b1dd78bdd31f0ccd98fb256b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9637cfd1c9394d4aa79afd25447c7163513b3f63fcd0697e396871f0dfacc6a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23ac022576407c6789ef3c1e69f536508ff20f93e4cb7503029e3339d9e3c1f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c2e73d11aae81f995b924eeaf3febc65c20ab36ae90335ffdbce009595fee1f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3515986339b4436892577d2c8591f02be06428ba5bcc36bf840009121b05c70a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha03d44f008b208f58f9c54080dc0068c4c5465837de0b5c06a28bb15ada19b3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb6c5dc6eb637c10d55384573e693a552aa69b6e15ce098e52c006561082e574;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffe8a02b4a287132da8128bff6ad2d74d4dc64015bc5cccf1c22001c699f352e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0c47b2736d50ad9eb7d9ef90695d90d0e16a06430eb12924009bc5af1afe001;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88d0d3ed5106175aea208efa8dc432e69e0bf46c19a75408b2cd2205e7efbe6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda6895f499368fe3179c00ffee4eb920bb33356686c52a1b5e8640d388f1a276;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a194b51e549adf1bec562ff0abe2e62f9c829da56dc910060bd542435edd1d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c23ec6ab5c9a92c5ee3b51a07da0a723eba2f00d2f009f1c921159462a9b6a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4026450afaff77a118dab025924e1701bea47ef10aa214e40d1117ab5387114b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he636f30b2e4815d3fe3ded8f30cba77f7ab1e4628bbc29982e9e1aeaecd483aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc510a87256e4d21d3d7be65ebd4524113a989de928a2578c0c65e65b80bc2823;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h34a068cc09d34f1f6620e3f876aec99947d3d6d840d086095db6fdc9759e482a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3fbf77e7c4f78c435cd1a07914c06505e6aac7e4e260303274a45c4e88e9303e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h314ae56bac35bcf5a06503e8dc7dbf5458fc65e007c938772be45d1d02d2135b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7ff8ad8e0fe741257d41a8b35cd7e080a611b1d9cec78ef4a582f05b3709d44;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha94b72f3d2152390fc82bfb264975e1ba13a3458a86004b5840d636ca97ef470;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c25bcacd11eb66b45f01ce9783065f6ecbebcca44e0b2ad4945c0564b2c6ee8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb31adc5ddb44428c2ebc2c1b409271698ae3c2cb1e351afab66b69209b89b73;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c6267cc39e63f8ab105de78a2898487cf4cd278e335870beba3dc589b637f29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h855dc9a8a54f223c3b62493e353cd4b91ab7fa9ee3cc408b9ddbc21d79deaf3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he11fdd7a78d066d85f5b91f754c6c2e3ab9d71d30bcff1598912b6290b0ed88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6bdfe9bfc8a33fb5d25a489310b47d4d556c3732f11b5caff82c9e6cb4e23485;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha93eb8cba2538503add6e8f131fa82e87ee7a702ffb71e94b8995699ca663cc7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa3a9c5c7e28a8d59497350ed7f0d83033a7f2b472f1e02879666eb066797d66;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f819dd6014773fb004b819ec12e9909d578dd045fdaa13a3a4b6bbb0a7cfa90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c115e8037658175475166f31086feaff93b843b035b5fcd23efe289797f51a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6228ead9557855d5313a6cfd8ccbaeb78fb0de34412b70f84bb914e3c9c6552;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6bc1043e229c154038e80402feb5693db3f84f98665c0f3da0728c73691fc007;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e9b5dfcab04dd6326fc63abb15992b8a080edd22a4eaad8daa24c440803d428;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8cd814eba79d82ddb700e7bcf706a5497d337110bd293d44b0b0a028f18a20cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62de4accac61eff79ae00de8e05b88da09815b1cb2778acf89a7dc755a514b27;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha34d5f96722d830b3a16aff82548a9c4f8f0056c44ed54e9995610e3c92bd4c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h786ac0a8aec46cba4517671430d260d22a3e69479ad3beb04c232d442f0fad4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb35fa416e62c4a81cd680f60aeb08e8aa3ed880802e31a85531d299a103c7454;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d8764a431309cb4947d84877eff25f89d886f2ef09a17d27c12874f0308b530;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6df2f4615b02cf4472ce62692a1aa2163d37f78ffcb78f644fda4427d4cd565;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5940cef91efb17f2992ecdf419e1735a9e1ea87c5df0ab66eec0866a9fc82183;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf66caf6bbe32a428cdb4edbf5517b70ffa8237536546d3c1677e660514997641;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h29d4b1437368386c3ced98936b8928b88da78ee3729f2dc921e26b2a54e06b63;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h460f6f7f91a66941b799ae9448d347e8ad65d035c848fef4d0f7842d9be9bb91;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8059bf370ef8d5ebb7460b72852ae146edff99312280dbbcb81edb38d22f373b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b55ce0e7f904d314ee25b7c287736027bba462b41f0d165086a88aae030f4cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28958d542157ee02f5411eab480c986a9f0215bc2bfd5f9f2c684b0df059e04c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9dcdfd501f546c2ca1fcb8791e70c118b0e5f5fe2a6b894a202fbb3e077c774;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6fe858f1def7e01b2238a46dab90959cd24d880aec6cc7b3b641c32cc880a2db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e5034302bd87d7a3292cb117ffe4d4aef6a471a7bc75c13be05dee95b6515cf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he93a1849923a7000ba82183d773f7c570613eeac8dd7a07ae3ac784aaca0e339;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc16661b40261013bfcaf2e2949df7afae95b06131747103644cf8180357b3bbe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h692aa5d5604b4f4a12f6041a73b051d065f511329eacb15be681ccea834bb2ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57b1dde47df3370495815f320b7139d33a62b4170a8c3f312439b4bdd40d0cc0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3cb5e6c4a0458ccfc9aa487fc5779e22b2c484e9f5ad97b3633e2e32110ab98f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h34efb848f0656d10f0244f5f9dc0d3db6be1077c7c59effe92bb1ffce05a6232;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53aa8f35c50e1dc16192c888519da3e8fab44f61b4d115b9b0d0322fedcf3962;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc29a4337591ea5f9f232fee6c19ca8d3f297118a1ec864a2a6fd6b4d8e60263;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94240368e2974f2b9d425583c358da7f92b2b545a8d33b2b24dc3e8a82f70d01;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70fe0e81200244699d934ca42f9180d746479f309c218d3f38b4e329a43cd070;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66c91bfe93a3ee9f438bf7ece1f5d52c9f30995aaf73d393adf9d5736fd57601;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae6ca33cf4b14fa852b27d41f2ae7e4c594554c4469b7cc972385fc9536262db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd98b6b09146b6c056166c29525a551e1ac94c16cf36ad218c4de6ade835e7557;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5cde77f3c0e86f736771fc5f44b82b0fbcf77afb006df633845bb65cac3662a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28a9dd0f63604f9368f3d7d4d151814187dd0e0f00f5eaa35e42dd0479342506;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f862a386d8806169a489c174e11986b21479b2f9cece26849d5516e886f71f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8d927d04d02c93e78bcc0c306869ffe1e1ecaec589a790b4a362b22b1c901e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e5a2168a87c37d26ba923994819f00ef5482947fa0486bcdf4d369864c75d92;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93ffb53b257cbbc29b1ca2f302dcb095f7ef05b29e2605033f4d6361f73d33d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb68f4abaca487b5d6915d98d9a87bf07e49ea67090ad9f75dae89227a419de5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff60f9c79663b69bfcfa4eb8e329412fd0277f5109b8dce20aa0c63870a8b54d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4408056e1ee3332e60d34408789b5814b33a71a399f6f6f2d4d573d276cb0238;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd12206ebb9860d4749d33ca1dcd7a00b8b023826af017386efdb7d60f73164e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f615012b140a2319e27aff3689a86aaf613bd575980062ef83511a61e7b61c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1fb07741bf325f51f788dab557aeb9bc5d44ea709b6567d7b23d43c5f0a1497;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78394acf8a9c90e4a03100e088ceea3418e3d7c20454c8c19cde1cf01ff30c34;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5a51543ecc7003a5086b76bb749c20a8771537013b58ecd0957f50b63296b6b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb770cc77e6e78dd78bcd9c8040c56b24def84d31cd6b7316b42120e8fe1b6cc8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39c4f02b256c182f97e1e419d6398ca98120d54b04f2d3b64868b3f53a16a455;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb3c187a1b2e10c68e6609446531b33d50c3f6aa40ea4e5369cbdfdf4b4e393c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77c5484bc91341faadf063e8b7a27d7d625d66f19ae2455066af55730a0957d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28d5ac8f66d9266858a63de983c423c4c9191483eb086419867a09ac723afccc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h175f7f6593d95416fc91a099e79b32d8530e21180fb5c0c62289d03c0d564ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3007b4c8fc75890ea565f513aad574ea2a5a83a59e0beca2d24e39fc37c9195d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h795bf264add42078b3977c3dbd2a771ac0a5796831726eed1a3cdf6a7bc96110;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5bd00ebb3c50fac5ba073e1702c96629d7da21769fa6dc3319e57ea793090da6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hde1af042b1e2bcbf951aa227ca556107a96563a90dcf48447ccf1409dcc6e17f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c849fbff548ca9c215734654c1c8b2e4e038e4989c77f1c21d6f90ebbc0a51c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd18a5a8eb4418e57037c6b2b483fe0c487b5de77aae58303070152c021d93e84;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef82ff34c1365233890cb909580b4f6749042c7bfc03cb8ff2da4adb1a8fe971;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h208b77b28019710996473793ff6017c9496f4f20b779baa03fea0a91dea4c797;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9fe3e97a84360984edee627da7cda6e6f690f294af8bb225b03ac6af8160d734;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca70c4f4ec68f78a6cb37867412258f49ae27cb797c3703ee33605419878cbf2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc092832f48dff4faab7b47de31b272680c36c069518f08b596df5755afe30656;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e63788294988e16d5e39854db57c61f2e313120b01217a2fe35a1c95e488f4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9abc8b595612aa9126a37105ab76cb2fa7cec75069b60f7d820077e4c8d8f35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb729ab5b66f73b392d24177cc2807a7a027d5fd70702eb9d397d21deba193b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e5f26478303fe4dcfdc18c5c19faa7b5f14c4cd4b0cac985caeeeab48a547f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5787a829739694a29f24a943e5c15c2fd9da3d602936755e40bbd4ab6b471e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd171df1a3dc1819e332aa5c53f70b1d0915368fdaecc6a0b28c1b614d244f127;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1be633c40b9630b6680f5e79030d0bdbc1598d84d775ff31931c678548257552;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6626b9f49b7b57e20c9c3dedfb9838e45ff6ac69beefc5e3cb043a6949f0ce2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heeaa57346a4c4e2473b467e691026cd7840ba1a0300c3a1602784b46a052deb3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b7d4156de543ddcccbfa665570452999c8da2acd5510fef5fc0beb01b1e55f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcadb2787b5408908564203b95c93eadee645841eed57fc17ffed7d47f8dc59f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb375a6774d7fb2d9cbe610425251209e8971fba289d0006102eaac3bacc5a1aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ed176c263a721bbce0c553c2dfe812f2f2ecba4241454294083f3669b5e6390;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28fa575a3b7bef96ccd66217a631ce350734c66456efdf52bbe45cb16d2f43f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd3500363315973b8b4c98eda1371413124dbea03e8e1bcc1d3f13fa0474e7b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf025eeb873484dcf0bd193c16201c3caacaf6b517297bddd945d9739d3f51361;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6f2db929897ea720e1238903d29b7918638be60dcf240e8315d9289e43626d2d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf5949ae781e5557bf6cf23e3835e7b4df0be80c3579d34a15ad0f26c53206beb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc31b91f28878c877d5812b232f5f1f6518c84e0bca1ac3ee098026ff0b48ef8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab92cf4696b600fe901f6f0f3af1054e492f8ad4f9d0f5ab39d5d5ef984ce050;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6486cf600586122d8ab6432ff9bef8fa6cfedc8c7dea3ca815e007053086f18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4e61ca373f27b3ef7fc020f1218208ecbe7692223c00f0ac8bf1ab0fcef202f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a8b3d1c4e77064f5cd46d06f7446510c91038680b71b56ad1c5c84b87d8eb16;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5249a6a52f96eca0e1c9a9df3f94cc81b24dbbb6a0744f2749b51cb9e13233d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc681110144d4f751c839df552b8d8a0f6b9b1386dfcf92349ed4ac5503d9469;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfcac9301612a4106564d62a233f1530707321a027dae9c8031e794e73b6f9928;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9876458b0d67afb2624fa37e3c5138925e8f95d7ad58cd5ec310763a75b181e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfadd12026b13e7f89e7c715cc95f1cdb3c3f2d8fe9d32a4e71a0bda47a597c92;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f8d3fe87aa383939f7ff2216697559f09e1b1099b93f43e2514f6c38045fedb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5691f495c477cfedfb2b14ba6e4f3b2c91596793900a5498040c157c65532459;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb49c0112cc0ab736f27e4c3b57412c7d8e19a62ddcfc5be48de376ae373187b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa1b7baa43672c5b545e6a4a245bda2927836cab9b18c83bec7ec83959840128;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae21584671e9ee4c136578b9c4d2e413704d3303df9fe694b95ff5dbc0dcd2a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47b655986931a696efb2f36967dc9be531691d30bba0e85b4c3806c250871778;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcad5a51eccea7c22e48e176942c035792f51daec62c26b91563177fe71e8b389;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfbb22fe884f57d479be2b4bc050f48bee21820700b176b58a00ad83725eadd9b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61225c9edaf80ed0d3744700745b4a2dfbe918a0f0b4ac0b50325db5a9a462ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h381060902d7c37271340304c49ffc258ac9766cf87febfd6876e0e23b64eedce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d666a739458bf325123d1a093dd0a7f8b65396b62ec4efe80434f888724ea21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6757e0007c51b70b258b76e717042ad5bae89c1f89a98b98b681aed1ce2e9f21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ffabf0c837ac93bb20ba8c429d850f69c69d4313104e90e118d939e655a06e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h944cc77d4bb655fd35314ea7488190411c98044f7c96e0d6227282f8af11ca62;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h836a70621fdfd7495e709f54c5d13ea51ac6d9c3f00251e04b5d57c5dfe94a4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h91f50558753b3cab5c070589761b27f6fada619fb2bb69e731677985a72ac0d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0605137c361a7b0bfb354aa0df5c9927dfb34f852a45ce0f4aca8f7d19b5467;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca3cb1f6076ff392b933eb20fa15b4b061671ecb8a85b60988f265ce18f611dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h79e4ffbbad4c174756f7d328e0d0a11307a169ae74976e4a1ec8d24cbbc975a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h250bf588fb47eb67511fb21b0e2203eedb22474a7705ff507c3c4355259f8ddd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb9721e06c7b9bada7b809ef024b0ffcfbf2b949920774d1dd3e5334a1d00e26;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdff4d059adc8807a73db8dbac61bffa36e40e46d9882d45e23f5a91c73772acf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2c60fad7f03e9a1839a13843df29bd5c57f3d07ec559ba3d45ce07f39ad79ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d8dc81986eda381c9459e10345ee9e48494848515b1e8d066fd29b5c8d10c74;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h649588633812b64f601ce950da192413e9b6104b71812af3c726451783004c5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7cdda7f3987fc3c806e429f598a3eb01d40a6127d12a9c183fe56496431e9b4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f4e6bb7c56ce1bebe1dc9acb1c4a22d08f00923675af437ffb7d00e453750df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2237e4b6db5072e0334c56d0d19951734ce4802c349834641bd80f5299176901;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h303b7f284618bfd7955f3af8be21e054b541fb302857b8520b0134383266fcd5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h267886e54024706177214d6165d15f983cacf2ac451ca3ffc6c791d0d5d21802;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b9ab42e05c22da8b61a199b16fecbf223bfb3dbb265838b3aa59adfcbb60888;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49881a76cae590e04ca33784cd113a1ea4b545c58ad54c1cfe0986e4a446aa46;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbbaee51de56812b3adaaa0e77cc3dd3815c684191abe844ccabf8270bb6d5979;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h533d654b6da4e83226400475f11ac7e2db8f563f6f73dd16febd0695bb92d0a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf850aaf86f71f2f9f2f8ad347b6dd2f171eefeb8029559cf939a044528a07d3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a907199a1997775c8c4d266218e25c5b34a96f5288281ce56b88b71cde8728;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4644638b582072020cff6c11618d8237532c60d7679a17d385395b07c3f1ba1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc9f3427303b0e58c96a36e2cc72f099231f630fe742b52423d3f4a6c96864e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h901cfeec42f9bcd33d2f6601510240a57cf85bb93237a18a293c29be10768af6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b848e80bb85d1d6c75ede35114230b758412c292a681d153968780b89762b5c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd313c9b4bbb57540b8c143f2309baa5c320eafa9828e1524c372a57fe7ac372e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hade3e6870cd0403b971539bd99b7ddda1f7261535bf521dd8ec6510233158385;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb306d4276d31f59db44aa59e17ef2a6208a398249032eeee2d24dddf99815af3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b91f4ac8d84d6b4918fb20a6d1c4d9cba628993e55756b483edc7471e8a3254;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4b359a677938172b080f4986fff63010f361bec89f7625c3ed7aad27b35532f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h660abd739f740ede3e561104c275dcc9a5851f21830d965ad4e34cb96ea1a49f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc06536ffef64d52639bdbefc4e15b5a13c883fee0d97d3be2436b0dd74893f98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcdb7e21c2e917cec5b5e84d0d2328fd79981c3fb679d7f4f66b7c29c24f68b49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51e03c15208c0354e3c188d7fba62610a1a2b51e02d687e8ef0aefa85fe5a90e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce94c1d2954419b72cf9046c9bcf0c32efd21ff7e0c508f186b6b632b8bb7860;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc11524f450e2a4a26956872385280b7fbfd31a7cf5ce6a6b5ee41afdf625f15;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71a880f34627fb9becd091f075a4a50f7443ac4b4fde16848242aa2742e56e75;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc97f99df33ddaf0c3fdb5811cdfe8fc94fd65481d65bd628a04c1ae9a434bdf4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64f183cbfe4874615a49d8a037f7cecf19752b818b1ae8ce969bdac764a87671;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc921a6bfe074b25eebcd35642084cbd649e0dbe924f24be32875d0b11872e176;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc303550ab359908bdf13d62896d77a05ec01ebd0a4f18ed6e413695be3db7878;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h831a8fc5f0bd964315fb837f55076ec47d3912555650656b3c6010fa415ca6fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7299b1cc663655b7e50bdc154e6dba27402f825d8335753551bb5c97397d6409;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36f9e645507b9cfaa72241037dea4a6588fe90278dc7973b69bbd184e80ae107;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40bb548754e816c2e96812c1e781e5d1f6a9f0d8e2ffcd876f340e49f9094aa9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h123f49d23839a46a540bf5fd19367c8c052222301426327ccca9aa6c9920ea36;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47d4c7616f21d69436cc33842dbfd74741aef20b7fb98341009c4878151c8066;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9cea97d48c2b139a2675a7624011583baabb70ce8870bf60ab7140963ca6dd1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he278087b2148ac683654f8c4961d70b5e1db3ffccd04883bf35261b5840c6890;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32f38083548469fdbd8acaa09939963b9db6a68b67710b9b5687a8be655273d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4948814e2e74f6fd0dcfa1de801e03c89cdb405be8758369842d761fd36a5b08;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf25eb264c8311ba710f845e4b5eafa9f33a18c1076f52d04cd6c5da14d68ecb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99c2a513d5b8106170ffb6a7051040c2af60c1d743687117ecd98a0ed14efb10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5284fcbfe3564634ec41b87f4c00dceb9e90683c688a98e5fe54576f5da97378;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4804603fd3ff6a746b33c31fdbdb04515373a1c69045ae0d69201ffa9c465c51;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3de3b67c78a47f7bc22a4f6f9d58caad9e2921cfcedc3be369ee43a8c26ecca1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6a69a5c1010f4307dd0535df661580b0dde278423d25a5b0f60fffc670e27e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdef72f012ffb9035894e317ac172f674e015526de6db89ecd2e9221f5c97b4e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71d92f1b98267ac9e36daf46eda2639ac97a99cf454dfe80ae8933867e12376a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he81d66f0b2960cc6ad344a6eb135df2dde05cac7895cb2f93db58899cbf29d2a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd24be3d1907973c80a218a39e743c6e967151c8a7c7b5c48a8b7f1df95d97383;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8330d6bf146c334c97d8a2a30ec42d7a9f9781ebf6abf54f3d9af6001d81a53f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf405faca55f821fc24291979c490cf1875abc2ee2bca5f463ab652fbf65fcb7a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf13dcb96e5072340bc71dd8b99d8a1faa73cff366867276bc53a8e2aa413424a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2fed9eeea509c04c122f7676cfd414ddfb3c479ec5341ffc1813c01ac6fad93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb127a8d978ec025978124a2cec646ddd7fded63d1645d8713024f6dad2b5a587;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf30e645d0d9483fea0b51a2b237aa309759cff4374f38ddd58c6b62f8a9d2cd3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86eae3e53b4e03b9ec3ed3a208a7cfc6b46abdde45eaf7117b32585dcf025471;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he866ba0246620e90309caabc25ca34054165a207039742ac2c2bce1069d68158;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9ffd203152110d92b4191dce5c6f55072999531cf50044263b9c575f6d70ef2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41b5ccf94cb5cf6fdb529c65207d630157601eb6cdcef973124a9d98cc6eb8d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6b9fcd3e4efff54f05c34feb5dc0e37a02819a724dccfe4f0c74bcf1b143707;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5dd92a9b01aaee3c31ec93a2c7b0a62f9478bf9b3426595c298f07eb296c2112;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6457ae7d56c36abfe51c12c0948708373df15797f80add7ef9431823cc089ae9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd86714924394796a8b21af9c53afe7df66f207297569b19b639bc56c93f7f706;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d5a926fe8056bf8b6ebda86fbe753741aa847c9ea910079f3440926d2ebc630;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h14c13af9aaaa051a9c950e5aef06a475e18d4f11f16e7c7f7906b92b944d0311;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e652997af21969045508b125568b1610835a13e0bfcca06da6818c3560c0ec2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc490f77766b1bbd597bfd282fa880a11e17e422899734a7ba6906361bcc7b9fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d81662f89a06520ae798d7923a860c757e5d8ec4389ec8c8c70b05b9e3341f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3701a87f50ee210ad345b8c128843107970d6dfadae4fa226622619ebe58125;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f771ba011bf8552fd3d65226a0eb2cbe612c4a032c1f6d4080f2f3de5928a69;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd98f963dd145dd2d1c1334f0f526d78ca072248ec8f9689d6f3a8ea6458989c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha70098d501afdd48f2c6b0c33af6d0f96ce7f6a33594b18813313035b7ca5a4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd638d3cb32f5274ba7775a5cfa910cbb518ed14b53e5c608865f09afc087b9e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4dfcfd32ace0d2ddfd023118431e105db76f89046a27848308e599ee0b6014fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39e58032cea4de772947eee282a04f8d3f381030debe85bc7c2fbec762bb89f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he94873488eb6379cc132430e893aed5c6b653b5cb4abd5365055707ab439294f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf5582704fff933e2fd3b450074f9500f8a3c493b4db2ba7868e289fee1964b7e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h26b4f9a1c759d79f98cd7d512d6dd8d09b3d43dc5597420e8ab466cbedb7316e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ce3be1c7550b5628cacb218bc8521681f82f840fbcb8442eb31c9f7a7ff71ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5533e9a8aa5056e4d57dce14ac2406144ed53e72601ce645056ad06cf15bf49e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33a7797e7ddd84838476613037b6b05255e426c2634c7507a4b10f7cabc1ee40;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8bdc8dd1dac6962703b44e59c1d5a40db1fb22b3e1f289fd6dddc6acf53893;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c7af9eeee73b4d8a438b75437b6f914583d57c4c1e19d56ba41f8f91db5cd86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f2f6c3c8741d4ca810c57f7dce9d3b6f0bab22a8d03697b759b05f55f6fe7ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdee0c5da50dda8c31e19ab048be19702b785fd992c181ad1439c23918e8b7246;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ecc76b3bbef03f16834b990df60104fba546bed662908a5fc0ea8d7283e5816;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5030e673b04faa0e99a586ce46bfd88f77b1b7c0c2d483f25961ecfa4676b13c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haec6e3c680eb5eea13007ef7e98cdb9dba6ebadd6b8b705bc3f021362b5b197;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e0257f53e58da6a0dcfa796e6fb2eaae7ee59eacf59d2250c8ad5b19aef6ab9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h299ace18d77887752e2b8ccab5754119435e904a9c2a489e15980ee4e57512b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5c30949c016302901b4545662fd3aa666058b5a5082b1c7240f9c0f27fc20c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7af466eb2ce33ce9f9b02b9a739e8ac39ec7f70728eace7952c7ee9ed879649;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11b5c91ce95577b624ba61ecd84b4638478e63d4befe8f8c3a272d2b8334ea7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94a27d725de2402b348ea7bb8405cbac8a310daa68a4e9270a8cfdaedb9b7314;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89bf6fefad541c395bcefd928efdfa1a89fa334ef90a4cf034867ab440c83961;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb441a3b7a071256b0d1a98f496cc2af873275e5d1cc1215539ab8453ab5bdffd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0b67d563bef164856bb38d4b87cbf50357395102ac36e61948069d84fbfaee4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf32b4725bedce83b54488084e85074ed81eeffa8a41d4adea50119a55a3657c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2008e5ad1872c4bc6d0651080653f0e28b801228738ba943020ac1c27f0a009;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2439f75cdd693b4e431e916ab25f8b4fab7ed6d67a94030a2143d95486777a88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h783a9a24a93752a2d64534d636b32c2dc20d18d60a9f7e6de20ad5b6f420a2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59a7e1431b1a79d479f9adb46508ee283e80530fb9b97f5042adbcb9ca6a1c00;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5eecc6ec437d67a56d6c41704acdbb752608dc7b529116fbb51496650539beb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb09db74db7b6b024c415a5488779a6a853f84d72f7d7236d8d24cc4b9a7e102c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74b85521b1849a918d30e001652f1e4caa8179d327999df7710ecfe122446f9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b5dda9fca8db9d01208e1dad51046ef21ce85a9ec8b7f4daf22eb8ed95a24e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h609b6eba476db246e276f13903729e0894fe69695407697def427beab590d42b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2832d7b3a65382c1b5b180466cfe02e741cc2552190befea1e5d21b46ec828c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa5a3d41a2d1a3f9261e652254cf65bf58d3f7725347c97667bcccebed177069;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10cce990e494a1c238c90f644436cb56978cf282a8e6948ea635b1ef0a9160f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7fa4cf191eeb3ce16d3b2092a3e5b2c16eb450caac186afa17f17b2957fa79c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1085367cf27f8cfc48ca5691ad7d9b5f016593efff24e1eefe39d9263ba68283;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc244935d310dfcac5ff03768c476f26706e23edc03957946fa930054ecff37eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9579762e5f3af44ae5ee3a3ae0764ef1c198b78be49dfab9c76de2ad4cebc60b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5e30adfc7311cd219ee2f82f82ef78286570f728baf0f62bf3530a97a9c4527;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33046953e0f5ab085619fb9bbbbad96da674a0f0dab5d85da366a0125dc2895a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d64dd7c009d08aec6f73368cd7f79b3d66cdf0500ee077d71c668d62fbc8e3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c91c34d084690ccbcc7043cd0863506812e6d600c484f9f5d53ceb22c2cd0b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3f1abdd97f277c91a937ffbc55ef87c44873dbdb9a46640c7d600b6281ff9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c1fd6d1ea52ca7dea6f1cb4465961e7d4271eece55ef3e762c3a7d11692387d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98c4e2e39c50a1367bc1df51f41bd98ad9a8cbe55a091325baa6335f6571fe76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e368707b4714d079deb12c39f8cd8ececeac79f6047c6723c521582d886986d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e6ae81870c98cf069ab2c133057f50dc33e5b50d2102f8e9536a6ec3d8e2d3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ac92e5c0eadbbc66e4ffb5d341af6f02bab646bcd0a6a64e29ac3f3d5c5cc69;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb881a90b914fb0c55db1d3e7953a2fe7771f6637d3315f15171712bdec76251d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1454a672d1c7fb7207900ff961c5b3f3a191d96cb5d65c1d78cd0c35d8b65f83;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha10947461b53f2e55c0dc664a0374482168944c57ad22957918cbeb238d40e72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e0b71a2a60ccbf38c1cbced9af4a3308f50db35df9a629999de31bfc18793ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f7dfb7a58877f94707948422ecd0f4a81892404d5522da4254430a88c12bee7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc3c637bd489a84c9e2c863322415ee2be52cc92802a553a68398c8b41223f87c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b28d8f4b986b5aaebcf518bf58f2f7b081299f1f5101e5d6fd6c18d2895f57e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h880683086fe75197c65a1529c900df97b1f8757aaa8cd1923d7c1aa9b6f533d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92dab0150c9263d4589251499030a21432707369d47436e9016114605a05d248;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6272786a932d47929689306d93ebf4a162faea3220f222823ebff93f8ed214e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5288f187262686ac96f2efa5bccd90f6f06de654ae052733a5046e45280b828d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8e3e0d9335cbc5388ebd43489c00553e2e521a4eb8101289e89ebab20008366;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf82c05501dd1ffdabc4db9bd3986b3d31bba3780ece1c39900882abb49df06;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21a9ec18de15d0e1df0815351248cc76abffa682942a49f0e637581e4aa3208b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64db75f1d3ed673907d87d24a5d552d3fa78baff04b3eddf7e4c78fdc352c9bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96e89659473eacf4caba9af0b61b78e8e3341b61843ed333e5ec55e1eae90b39;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba9e64b841f84427cb1f85a3dd8f66d669f4ea3aa0f61203592db183e49613ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf2366afc7088f8dc9bcc3109a9fc590157851e28f128457608a0b60a810fb7e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e9f0969b190d6a13adf6c9c4ff20181710a09a9efcf6bed64efcbf361084a38;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9da8d73bf2aba19376b02c291924db77cb893888ab7d26a5de94e34e50248e98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h925dd2fb763563432c9cd483713d751cfb6ef32ac992e8a0e1c1b57a351e32a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54be91e10830a6b834fc27956f159cee118ba415d7ef4fd33e38a3aac918355c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94b0010e39953c9c3850c2cf53720e5e83f91aa492ed638ffd545fc0aadc2578;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hafa0405213f1d7dc30408780e5122265cbf5c33a51a1a84a22976cf6b695a7da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3589ae7fbb33500c85a507bdcdcf10080fa57c3022b3839e554e6d8a882fd95;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe835fc593e8c67fe709df052258c27be3592cc75450091854329ce80dad2665;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec6c04c8dfcbb81ac8544c214ab1df1bc3a7b792e05893d13424435dbac5a6c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56d1a1052f2a4438801aa75362a0202ebc6c7551b7e9941c274cd19bd123d206;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d1e17334cbb6dff728791d83d262c264c58b8599ae05cb0222a2792f5cac8e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd557b5fb2f5ac1f62e2bdf99dafe5244c5e8340e41b94d145a68555c04ab20f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4bf899b174616ecf52344185f2305e6b43bdbc641ae11ce3c18ef4954e841aaf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h453e8338c1588d51b33bcb7892033fdce124b6acbb736fccd0f33d08a5817949;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7c97dc2254f8f587253bb3726ce1e0467e5d4eaa08f8e9abe8becc7eeeba67f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h969f72b58209deecd095f9660f84d9e3dc79565c8dece2684d4074205281de41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h844ebffb50596aec9b001298dbb88f33c95120af5e7d432c01ae0ca0c4beddb8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f12e8a140b09211f82bc48cd027098f1768138e621e3b154fabd6f393007c8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb2c3fc7e3cda8b12eb16a6b61568240d403607ac0b51c2b71f636bf2ba05a029;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe8989d003d8aa04e1ce70c733009261ed07179b00698cfb28c14b545c178328;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a0dbe38659429303d1d1538ab4303bbd69f9d51d57481d38144e95248c141d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74aed5cb8bda325caf7e8a72c3dc6f091bc2940280f6b676a0284e6be57c7ae3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab3090c6530ca4f98b1c68f47c467cd0948ec547fa26f7f3ae3fba4a1b577b4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h735a0f861ccdb117b3ae7f0ff49d2e1840d7aaff6d7aedde0a87562a7ff7a44e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8591a4d7d009580605647324f15969472f3ca960164e26e1d6375dec92f23e2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h673f96a6a252d3f4f1c597c50d2e889bd5d1c15f1408c0b36e6a50df46cac12f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb191ce98f6407bb3c3270134992f8764e4ac1148f4abed727f4d1ae8c27ecf17;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h931be412568b11d85ad7a3e43410653036ae60d566c6b39327b3d6803f5e0099;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h22c5ef2f70ea154ae67905fca4c72f8aeaab1afcb62c0aa85f8a0f14c39575d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h374e34c4cc466d1d1c20f09e5e837d28af73ac8ab40aeac95940ae171be6c71d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36b58b81322bbe7dfc6de5b0828e6ef608276121792fe65c1ad4ea62e67379ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e02c2024e2dd66f3913df948f7be5f52fa523e3578e1a16333197c463daca30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5079cf847dd38895d9c811115c0b4d5264dd3a86ab17c6f0ae3cf1950d57207e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda0fd1a7a9c8b02bbba956afcefb3f7a89362b6fccd9bf4a68255fb2164c8f4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2cd72ac824e64d42bb7de4204473069ef3ab3ea2f21adb31ae65fcbcca6a7400;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb81dc80dd729076d14b5beb040fa60108e014c7858ff63236beebb4d4fd13328;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha072e588b470d5b3cbde23dc693936258cbcbd038a16f545dd5586992b149ee5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffc1cb7334e211302bba7829787f71b9d5c7e52738180ddd417608de32f13958;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab57bd33a2f78f383399ccc404c0a8301672d3b32751354f6632da0563c928e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6683334523119ad4cfcd7fa00909042fe2d934a67c49412c4d18a10ff1feafc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f652677cf84d548374cace257a09777edd573077d7f447070c55c7d78bf91d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9f52f4817b413538ccb0a2c8829eac708c2878573710e3fd0ed6c7ef7f63de2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h732b1e7cb0ebb5e8f639bf859b87c5705f9eed12f6600a6290a0459598b097cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefc3ff68673352a16f179d6c614b4531682417002c23483cfdb08156e0c0a3ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h275cacd8e671e46c9cb908b759335e52464c27290233262cce6bff16e541788;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd20bb025886ea6cb5ca84262f8d9069db71eb759d094ed1d31cef28ddbea4846;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e3377bf3ddc14be5935cb615077036051a2e8e73aa45f0f7edf91e78f91e60f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1a8bdca3c641070cd291f78c508e044394dca2b043755f8689fdeadb1371143;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f2553f39d7c8e0547b554d7432fe6ef5e8e7d8f671e1c8f21adaa583f092bc3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6fd773373449a8cce9052b14a9a91f4506f8f4f90bce8fc568fec1505c1842e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5552afa10e4d571362e350f6d6956170292ea670bf5f22ec77e2c119331dbaba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbad02904ff03ed4702b8c2f7dc5d5bad5713defc8d8d039ba02f63f1a564d918;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b4ae17ec7e5e26c534d2a33e36fbd5aad890a04ba10d5c4099fed7fce95b9f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd635f12a221cc9803fc52357b08f847e057b86a25f6d86861e8abb99e2afe6b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8b2b82549b2c6ae2196683a4c43ebca58a3ae33cf49902658e8dd6697746f14;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h685f2dcac5e49a27ac8f17d8e94c33509bca5a5efbcf3c3073cd777f63008f2c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7de5046adaf1c5d4db3a52a0a64c06b92859822c2da59d5e8ad01de2d6f68f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc197a6e617f1bb2546cb62b4b45e87255f061adebb72464e99b49deba6e56200;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d762654b895b16caeab203c9e9f715af2fb1744c127dc5e04ee78ee974e0319;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9bf881feb3869ea68230294b7e021dfb1c6a50449643de54db42077ca3fb30c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hded6aec6b1d127695414ca8c258116bb9b0213b0f0c6d3a3c40739f918b2f33b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbce8c6fa9cecb916264bf415cce2aced9919e871b7028e24cb92183a81c773d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28790bf110c09b300921efbf10a086e076c7999dde39d910ee8c73b9772bd960;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e675ca20a0c0c124bdd4097b5c6d6b73049a9f5234ca9bee2ed0a0156ad1cf2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d2cdb52b0466f0d73260a1148bdbd69a89114cd167edc493fd54414f321b02a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a1da018c37328b8a9086a8a53996a75382d0ebc5265d36e727737bebabe9378;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h587d01c9e6ca6a0c7eb7cd003f162b8c5a6afa4444c0bbb51c47125e8119016c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d9d847f69835425f1a937d38fcd110fd7e05a4d2912c4c41ad7f8150a28ed3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0dcc58429c89a601b00e18ac142ca9ffbdf04d4727e168f851f876c9f479c52;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbbb872405d82b0962420e6fbafdbe79cfb76fcb777a2c8147ed3f552ffffea90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4aa82d41c19b03b66d364d93d38881ecda3541f95d3ec88772413b586c23d8f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd1f12f9df5206014e6f53f34177998618b20856f66febf9189cb1dbb7b13f21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h933a4a2867ac132081da25ae5dc5e8e2d7eba839cc40b2c2d55898b92576f576;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a3b0ec7ae32316ab8867743e71c4f8f3cea70eac3399f073d2961af25ea75a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54dfe0b54d54d0d4b10860529be85bd17bf2f5cb298938cfb33aea27a3a8636b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9234ca1a177eba75bcb78d0ef3ce95158e0c53fb7c23ae31b4b75957e65d01fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha332e180c9fcc66cc30366c28b1ca7bd4ec03929e7062393c835770e4b916f06;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h529f6dc11d6bc358cb7df7a4afb67177bd1e02cf22b05d2855f0284ebc094c7f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c4dbb8957bfc62393d235a2bbd893dc490fa3e49688946fcbf0483da54a2493;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h370371628855a7e9770da108574730255cfe780c3b7909fc56f3de6b7f14d18c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36fedb31e6a1399c93ee20e33bbd299587009d0b56ee56427cc43ea3b2795d22;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbacc6f7a81367a9f1218fafc7ca4525222f152ba2d3d14e569c004a178950545;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea81aebac410d909d1a7d89e07e640554e77e62924c5a8684043277e112771a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha507dca4544ad5273ef9976b57c9663c446bceb1fde88626ee06cadbb1daa353;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c88cb6f4ea0d5e7fd124deb5c0ab855e76d575aa62b7327de3cb40cd43995e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93801718faeca99d91c2e55ed6ba2789ba9a329ec75b86c67fa03b44c51e4d77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb2f6925b953c412aa12a2d443ea1f9d799733fbb78eb6fbac64ee6e1f9ebbdfa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfdbc6e8d4a5c896768e5c4d6ef14de498ec3fd197fdd71bef180003f07013416;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d9b3830dd898a9d4260fb68e37734b0b6da22a7b56ac09bf6661899c31e10ae;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6733856d1762dd5be35f19861d368427f6db6d46a1ce8cc42d62d7db5cf81f99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3401f0ed67e6145d71b7be87a5e04d5104cb06c43602e334eff4543d886b9bce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h660b4b857bb977e1c3507f9ff118827eef192daef720f17b558bb96440f17142;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ca036f91d1732948107bf1cee3c82df8dca8ea09cce60b8272c32c46d21cba3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h30f2c443afec2d0b142aabd1ed3ce6abb96c89300058903db318ab83e86ae76d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf55a265a71d16cfe7b49b925bd2a6b24ddd8213018497512f64ecf70a9005fe2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19fb05b69cb918704715b42d28f6f0a4e5cdd24bb0d9d7a4d4f0f087c529182d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a5a4a97d59530380f2f7404b1b0b1463586ec01e4394212a4372c6ba4ea8431;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1cfb539b1e83938bf96d424a189de0c8c6d80c8bcc63f3b316ee0edb9ba767c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heff913aa831cf8dd92adda1879e527158c4d49b15ed6f0bc2e5841888749455;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h287047b45d5da92c9aae6c003b32158fabc046f6835ec4e0066f80d7a943b234;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12b6a8d043269456905263a4c75a002259719fbf6b965e9243d00b3a50eaca63;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e7208972e184acb80676e5ccc3c483dde78ee82a7d4ab341ce6396c2fb513ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa08a79f51037cfd9f376a7ed2357b30a3d877fd777ca42d20595587e5ad9196;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h411c127a68cb11c160891fe121b1e743f38f0a42ce456db96df9fc31c2125e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f737d655c72d1c233a52ef63c08ea309cf783d425fa6638cb2bbed5e9d2aac4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb60ddaa6a4a4813a641d6c8ce06192999910015d5783db58ca0ac81a48db3590;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd03533b24b27996165daef502e4de0562a44903087e99ef732394d7176e47c2a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d24d0a32d6125ae98b33fb3d82d0c89b53a0a3a980a6504ea9413487660a101;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h30958ad7cd702f8acc1b8d3ad0c78ebc8920b504791730ed1c0275116d648483;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e8ed645a3b01f52f47633bd911d15897c49002ad347bf380b16a257440f2532;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf7551b48dd0a54994c0a5aad8eb566689ca251a0906721d6e0bd79a34a74674;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae2f37215ab7e62736450229de00cde612e0cb2dc00d36820ae2fe345208def7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hafb6527219193ee41058b1001397d8332a2e531b770cecea362dbd9f39f2dbbd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he15107a97df91bb1967ecbf9e936ab4fbd1282385c83f3b0a667448117e9840e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc83a5ef769c9c28be9e15cdae3abd339cbb98324df3ddc284c02b806db0a37a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2bcfe105b2548fd9fc256ed45a6d46a85bb4be6c1b4d38c253a1c90c15f5b2a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a6174dc0dcbfea2710a17f0f9ac88c0c4fb5de10fe334cbead715d1d70ef29c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9cf4f7f319567bd641fac6e8204999fac8b01189feb2dfa0e1c59040cfb05566;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8fb8b2fdb3f64ffb820a3f1c8ca59cbd12db92013d7439cdb532e1c5abd0c17;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66b443b7df86c68796680fc03ae9481be18f3bd93b2ed92f4d909fcb1dae5e05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc65b8ffe2db922e4917cb4ed6d50cfe44574ca3b620245622321a44f24576e16;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8c709f6927c44a63d0e611fde01d64bf7602c8571922578ce7d3dadb518230;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8fe313c659b66e90b7f430e8b2a66b8aabc0cd83882db9f179119455c6348da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7452a5b6f193ab1dbbb2d338d749bfa44792133494dc8f7966b5446a9edb4e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he41a58decd66757631566d353dc22317300eeb3549377ea5f4aa4449d40c8ed7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h79d1ded13ef3841e40744d0bc2af38de519bf613b274f3854cbee854d46a494d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd9a15ca5f4fbf2d0a216b51af1ea403478c2cd53873588c94a26e91e20ff8ce6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39794dff768b07fbbdd591f1b57f8e5b4eb288577498f2c5f3e65731697d3957;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7327fdba51527c68733a934cccf478a8f5414ee3b3046d3eb4976de9b0413985;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92452e1f094d8a64ded30eb03d3e610de70c3a5ab8fea258070715e2929eeaa7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e9cf329ad9646e3b3350e331f6c53ec53bbbd22a4b0103f97f39170f0ba510a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d0ef6092c7e29cb109377a0d74a0f8fd59aa4a61bf32c8c9a36ccc59161152b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc368651d20b5fc85d578caa8de3a207d4126627e8c60ddbe694620d9833c62b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2581d48d60d39c70fe5859bd2ebf5776e0913236269fedae7ef18c281580ecc5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h648494c5a30d829c008aec6d2011c4c137a5112089cfc3e13b5861a01194cd94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h401ddd5e71b251c4de6c51fda71086d68a9762b5cf5aa9de97f17eb492d2b8fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d62f5cdcdc1dfcdc26899bfbf1200916032dccfd9a88e0071ba8ef2a8d0ad67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heab0d80a5328d145069835ee91f20669d4e04f042efdb3840dac089a8760c570;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5e233418bab7d9727c513671d536f1ecbe686f5965b4440ab5c1e63fe329caf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf58eebae027e45f9bea0e2253bf4812ed1267badb9abd09dd214efaa1e98f35;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he33e6cca0a64dfc4438bbcfedfd427e3676fc12931a11cd00e2900a466b6b845;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3792295d915be72790dd0fb6d4af3d3d4d1b374858d3774b151cf3f4fa9531e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6437d3aca119e5f1afb30af397ba0fd291ee1fd63ccf02da473db128cce2d053;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75b13534e9c9d54524613fbbb25406e5c2fe8d4cced88763ca63631881133143;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h30ec19e971d313653aab6225a9a0c953be6ce5a19ca6e5a96d28ecffeec3bf43;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8381e659762a3241f7f9c981fbb0c20f7b724c8c3765d0acde8257bc4518eabb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf0086ff05ebbc761ee04a1d22bb450214a978771870fe26a6bcd6c25526e4942;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee71bc63ee6e8a00adc1ee03e820536feb742203f16e8910bcf314bd48a3cff1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5be0507ae7721972ef9e7bba6bf28458d88fa6a0add65491892a9e817de413d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha78352f28304acc22982f0805c107038d86022c48db02fbdbf773ba6934d67ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e2b6720a09f4ff54f4ede0101400529e99afe35b0e8fbff87a764cb0564aede;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h295e21ed1045967705f86d6dce8274f8dc5caaa3e1327b449937e5e36741d7cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8b00345a3ae88de8957e0ea50688b4e89a22659d8ca780bd9a22fb46354b6a1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h79b5de27b51ea28e91efbda7c6e7c36657d02dd8c6cf0dd17dccc1bb47db626b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb463f0b6c9ea1b068cc2f1d779780619dd9f809729ae6b6a7209c444feb77313;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2648cbc297601167537a0c331f9a72fe6b0b7488ca1dde09c6e3b4eece74c8d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he47f76b304c9230fd55fd00de29d364fff906d8fad0b75d31be0812a0ddcff47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5875a4f050af5ca422df5d4e47b0f0690d15ff9c83cf625c6a1344906b512b47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h562fdaff481c11abc0c672e1b8504eca4656cfa06f83f226f6ae4271a7c4c9d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb12653e14c27cd5307c124373fd5f73c983ad5268eec81a2c9e0d5195eb9c90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8baeeec9ecbe2ee4130404c75b182b99bed383df0692eab7bc199dbe39abe9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h242aaa707b7b94597f806baf7bcd0787f4a4a3b152a33107dec61cc4cb82060b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7882e1bdcd9d14fb3470b3b74574216f204a6cdc6d44f4f2dd1b88b8afb45668;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4467e61ed2e906152545acdb81823daa03e7d96c84bca85e1f313d5dc9dacefc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ae2629336edf2780e60f9d0d7d16c454e3012dfdd7db0321ee346c8f3cc67ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4bc6f0ae1034c719fea5e4173ed6b51133392f25aea6d3edd2d3555aa715fcca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdfab85bf76ac75544cdd9ff2301c0fc4ee6415758525ec37a49c4a60afb3bb91;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45b529b5504fe8133c3218eb9310d0ef6324e88328b6445474ed648b2ceea0c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h18b94975bffdb2062e94383973fc7c015498da91dd203315efda7bf007ed3598;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b78916bfdbce05ba673130c65ac71c03f2cd91a58497cdd6d1bd4aba436ba3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h695be3dd65e16404aae6a9d5fd3128e6207e5bd6ba31baffdcbc185df90a0fd4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7e2dd557512c10b89fb6228cea660900ecf2d3b342e173fbffccdeef23e416a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38a653421ca08433e95365e7fdc37cb281cb4b1dada3f1504370171d325f808a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8372fb1e8342d2299b8b5130162cc5df6ec992fda82feaeefc1313419c0ef6cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39d46c01a0b1a51a7536c21047d5c7b9846d71a761040c7e6f402314d1bdbe63;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd71c9641010280e1045deda5c4e5ec28f788cae230232b4961ff3a2b645ff141;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h313d1bc9575305b1fcd992327dbc5e872aa3f8c7191bb23993081a1e8e82aed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2fcc9459a1603972bcf9897eb598af22e561c77bba6497191f811a11997592fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58ffb2d6a2ff0d67bd76152a540e55a998c8345f526ee84818e8a16ff239ddca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1cb80208ddb31acb2bca1b145747c8843a9b5a4ad5dd94ed98495cdd257e35df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb8076068896c28365ffeae47abd745919454469488cd46ad0e5c732762d535;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h612f5ffd8607aded8cfcb38a9246e6bbfd2c72fe2459ec9804c4ec13abc809b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he6c89b7279010a0584e79b8d75628bfc048ee78de0529ac7f7c43980921a77ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h175b32a0c6d9f4e8c16855da52ff1dbdc829d8cfaab2816f845386557745aa8d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3c6d7befcba00b5640396871e982e22c5033de66d61f1b606b65ebd81b89697;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61edb5b18b00c0f31ac158817aefa24fd9a150f2abfbdde0747b8eda116be665;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46aaaec7cc5314a3415736340133ee89818b7cc4decc2f11fefa89b7f1cfc978;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a7d9bf2fef2b5b8b84948da7578673418e4610199678e4530dcd049aae00c29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d4eb84c64cc85feca23d8e9b324c42d0e1b8ff8ab1ae6b259e1016c20276cdc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2356edc788ce43018a430a63f134f57cc3223f88d666e61d5bee2a350e29c65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h953886ed697cb96f8ff7de9bb9b5b70ff0680a94a7ce9eff0a575ce46f78e762;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf355a2c89f7d01e8a647f892c20f6211307c52de79dbaa943c7bc3c8d562aa3d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4996eb1f128af41b7ba9b64e123b3b01b547eddcd3330386e89f76460b67a34;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb219b5e26b050ffa46b2a1361cd2e6d0e092b0260391ba23a3007b016af258ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha55291cfe866151003c4e17be45ae806a22e973d69824becdba5971ed450d1ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d69cbe92b89a20c818a99585838d660e7470e7d77b7a3c2ca43f3e98b0ed9cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha14f6233c4003619d10117ce6093a421de7bea68c431c01cf4e4bba203f0aeb4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9630f96608cfb34d9e2b0c413a2e53e4073c113db5d220c814c792951e2df68;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfd07f271696709cb2dae11f3c1d921cbaaee2d27066651eb681130c31f2ed6c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b06e0f383fc00a1fe48bac87833eb3a2495e758b4424b57c59b4041a4114d32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4613e07d77463336f7f700c97e0470d2a8f00f7be466b068d5d3918329e95562;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57d82fc281e55c29719b722be7cf36ed1b9122e6b482e6fd898020b88579b905;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab6be18d256cbc7e354296d3f2883ddf4893e75d039aca054db285119b6185dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h659e82107ff040322f3cba4fd840bc6eb0f6d0d49f90c6ad3ce3a846b1ef7e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4d5ec2b62bd2bf506ea0bea84faed92a2568d046bea005193486641ca8e0e34;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1868c0ed5ff3672932e6490b94b9ccff0a9396d169ed6b49654abb57c82c1fd3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf18cc3cd4e9b92bc574e95dbddc95e3c8989992400184a2baa9cfd35d008d99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a3a9dc52428c88d48f4dff8ec62f5bc13ce302dd3a6e819b1d5d12a8dfbe1dc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74b9447a7d62ffe3c2a2d9ea5e11aee31b784a3ede580794ca9639b2880a122c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9574658bc81cf770be0efeddbeefbe790dda57f4738b7f5808edf78eaf2f61de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hece43ffe3340dcf15092534ead8038ebf0c5cae19e9bf66722b0b248f2160d3d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h67f2cfc070e37da10d0eeec37bd0854d8ca583584cdd1cdd7661ca67d78842f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2fee5c2d3877b2b1a2312e10212ca5d6bd9b95923b08c994f3da2ee3732749d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc34dafd3f2866b2563481cb183a6428a51859b830c95c3e805b5c24215c6aa6a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d1e253e01368be046dbef6a2ac7364fb7e61c713e9b77d02a9f60035281d530;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4462cd6d5de0c54334f54acfc9e1c6f127ff908b51634551afd8f3e8dad282fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45cf3dbf0e107b90eece5cdddcf40ea2c8c77d922ab55786ae1bf41596302f21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f5322db414fa46c8df5190df9b681df126a00bf10645ec8c9f76ad9d25a37e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf14ddeb0ebda225bddd6b66895ecf6761abe8b0d532b5950ca0479e3fffadeba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7bcf784693f7d93294e89637c4251c61131882dd99fc7e98dae0c15a662ba55c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h750a4f78c60185f71323fa9f6497ab9119fc80750aec8aefa207f2efd9e164af;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66219392f219627f43b0e8ca6a36653fc4da901125b09ffe3f05bdc5fe7bcebe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2af390c54f57f326b9632b3dc6206909451a47ceb164455484d3fb720990adf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9962c80874a84ac0a635cf1383aa4e2d6bb88d1d2ae9874b2bf82d8c1fa0fa1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b4dea1aebb3022ef2c45177768d428437b40eb2258631152e0a73da7ee61f2d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4048b3424d89307920c8bd17994c29513487883f04ea28362ae4586d22a316f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha22cf38496b844603e3e3c33d1c3cbfeadb339c1289ed7f6aecd32730b140fbb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c8c74b37a9d7085d1c9e8c58c3944fd5d65e8c8e271ce1b509f6039514a2e6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d8c91ea97ccea8d8fe77078b677357ca9335e5b186ff7eb6f68c8f2281295c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h939d0696bf36c1147d4f9a6cf0337809974746e35cfd4536202af3907c48f8d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c92d128b26ac12577073c2dcd8d727013bd89c1533a1b8623c8d026ba4d6e71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5adc25c26273fe2af7b6b9d8fc5eac819d54d0af65064a7516c6a0fa5c82960;
        #1
        $finish();
    end
endmodule
