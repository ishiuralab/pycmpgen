module testbench();
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [15:0] srcsum;
    wire [15:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h126c0bd081cb211fd4c9bb72e837e3dc20ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9a3d98c057bc6b2d1264825c914cf774fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f16232cb14d5028c4c216c4c45ff37cc9f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he01f959d53f96d41c5fa04de741cca020491;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc35b46b0d185c16d23448897e71b7302597b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99043c8bb5648f945fec6d2beb2ac65e860;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd82434a2e27fc0f6f43f1192ff6ec6df6d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf863d9b84ce7d8c626ad23cd7e3d78e354f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd9c59e4eb27209c8b04e3865594be7bcfef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66f048c8087a7c1ea5c6803c4d41f0e39e57;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h531ee2ab9e64365a03be22dc1ad24431d268;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96f5b9c0c501fab832556b622b5b59736857;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d53608e6bac772b19c517e17253135e1729;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6180e197e7b5ee3bb3fe9e0bd05489c24c55;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9171ead76bca68221199e2efe1836cee1372;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ef9bc5304d2df7a1b705bd1b9a630551fb6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68a6bb141b85aaca7066d787982fab42ab12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2db64b80dfa2e6ce2bce21cb5f29536a452d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16f1ce969b61281aeb727fb3aa6e775748c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h823cd15fbfa3c36fa81d9cc523162e3787bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd322748b0552d9e8ee4bfc09f720f52357ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9210f655bb5ac70bd0085274bf27f24950da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h663aad827e05a3c1b0de86e845ca0efa1dff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he22cbd5bdabc5e28e8d63f814bded0cc3eca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd0bdba0c05cbbdb3e4a4e8e4f878e51c970;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33996abb6de7863fc8841b5018614dc6389d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9653193d66cf118b6107b1c8aab436d6f613;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h725650118151332ae694bed6a4a07ebe720;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he42bbd1796fc85aca9f7af7da6b8ac62af65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99fdef3104f432c0f02e8ac51aa8485d5aa2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cd1d7abab68e4e8baeab29fbcbed89aa51e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28fdbc5c10a1576bbf8e7f232842ba298390;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4494b2f3a51332c88968f044b9f93718259;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63107ad13b75c47b0af38ca885da7dc1ee29;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bb4cee07a4b195bcfb683662e2237263f34;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c5ba2ed02948de2651473280f75ae1a2ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74995320d88f14ff8b4b90f35d680a1d8f2c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe776c7af3932faf839e7a3b1624bedfc1e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6075ff584ee24ab4851f9ce0110e1a36a8e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha18adfe15b077f81d2e85d22d24239192ff2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd01d09c234367f91f3cd01243789353ccb69;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff1afdbcc9c27e10c7df856c0cf661b99a76;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27467aaf4fa673e9165f22e350c991386234;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b3c841bc26d853222c32db4eafb8d2755ca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ae291ba59d15a822507da14fa7439e29560;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdefc07d404a1522306e0e21f4b61b703d5a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc4b7cc9dd5993ed047abee3c731199c4fa7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1afae32c71ae5a6203b67360c6e4854bb91d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a572da2a4782866df949dcf2bec677ad077;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haed5783132454027e4d8f994c6db8ee871f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h634baba82e5f9e7fb5f3a660e31f1f8161a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47e2ec981ad058aa13476202560669253a23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15765445d783a29db147c1bb85e6c81447b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8437487f6290d172e1566399162e0d0929a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a31ed1fd0ee0e8e6dcd8495c8deaa4ecf87;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c8de861aa23fb79942cfe8e36f876003fb4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40e94a32848660fe19f099f491eb3fd56bd7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd0d15076a6fa3d1624f1c1de859536f7cea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6feff8af265f635be729ecb01d5706bfdd8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h114822a965db04a489506fb55cb4e70b5371;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbcb50bafa677cadf3db6259695e589a745f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82d09d0fcd4f59f00172edd70cf6e199f13;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha3be91e6ce9b9288940ce1bba3af3bcfde9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6104f0687fa6163a3a377cc3f614f9615d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3088af90cc243ec2689c211d3ff0b849c789;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19c00d7e449f0019bb26a2cd55641939401e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1c490abc0f95ade87ffdf5a3af7057c8301;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe0b3d53a3271a99f39b53d6040726a68112;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88a156f5aeca699f5d5cde489a5583ee6f08;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde9a752b7aae56dac8192a807a2dbeafb7c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a658b3c438cb9365266db78192fad220fb4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed575b68b2dd652ca7cd02f3d1024ff72e9d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h342d9a0816268ea09dccb8036b530ed6e2da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8014340ed73952bb36833b2b5d803e7d253;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4384daa44dfb6db57ad28c4e7d9dc3c6a17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d6a36c0e6adfb7bca9d3e02da3d222195ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23d87ccc15e7949b56673f76634c752e76f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h107b0311cd76eff43da54b7873eb5de9c0f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h402e2f543b42df308b5bb3390ed73d9490c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e89e2d4f9a2c65330e23099fcc2e1b5b692;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb3817cd3d363711e5e95b82f80d0c26261a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf595dd04c43588f3c09fed9abd1538543394;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb325106a688c52525414b23866cc0f18d0a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8795236d9b6bacc8f74625c3f91871428ad6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha3476aadba32835bd2b3068a7f8b29f1837f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb964f0f91396f5d45f884f8ad26e9c738e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2189f444c5d12916bdf7b39a9a40ed88140;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0fe382af8a762ebbffc85052d675bfa75a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f33124324978ee46fc5a1657563ad4bd229;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd72f2a111b106355690ed7c1146bd31e3051;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h171914de77689ff855d8cbe34d31d5c00413;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40cfd83b61b86a9ecc60568fad867ef69084;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36bfc59d64e1a34c1cb8453d84e8564cbd5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h813362340b25ac4fefe642c96afc3f9a35a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ac6124e2f5cbc7590740f0eb432fa4b3844;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8ae5ba470f2ea7055b7e17ed75f1659776b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcabb518e10ffa953b1f402b8b2b26dfd151a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2e5a29051904fd45f11cdc74be21e97c7e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bc3088cc3fc47f66f0c4a3bd27e93b022d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8328f705d458171fd1dac53ae88c87a5b939;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc631c43ee6fa9731cae89df829161a8086b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h206edd1005ed5efb7bc3c397301cf28325c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61f43d6eb55603095c05dd59daf2d74401c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf8022ecd4479b203fe6d76de5f909a70388;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79b1098846a43eac895a2adcd3919aa1ed5a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h380f1bcab42b0ecc7309219b50ad3478303e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1e4df6ed69cd226debe25f0bf940a55d94e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h101322f97fdd48f84f31c2fd4802f04d52e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ed7ea951cc604788eff1119d440d7767780;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0959936dbf1fca07659857ce7451307dc3b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7f863067f886d3a7fcbf274c32e203cc4d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbb0a22392ae4293f6a4a306a03c63939fc1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb867a8f988974ae88a907389499da6a53dac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdee149c4667f489b32fba90cb1d30ae62da7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd382e4ce1bf4186040f41a214eee64b0a53f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2da334df78577ed67b133a7c347c8db3f1da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea55d5d9a7aea8b26221750e6dceac45864c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea6ea2ab1b1f815bb82eaf9aea0ac5d1864c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61709b985551e51d0c49e725c0c59595e328;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90d76d728480f5a5fba6da37f382cc57ff10;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h587768485e4c75bf4945429334a86173794d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb66ac967fd95b6076150ba8a8b9e650eb67b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h586d06cd10ee5b2bf50f8493532d4ffb6024;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ef8f90880b3f289bfa49e8cbc418d927cfa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha67a9ca6f174bfa3c174884e0b3fb1f29f7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1bbe33650bd5279a7bcd1de7df797c660294;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd929afa0194636e70bf1d6ff6c5c733f6b27;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha40ab257ec04c29f64fa4fd79b3f0b6fb14f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22fb47fae963dc955e161b4bfcf093b42d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b2f94715f7c880227fcce63e2c598eac83e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25b6d4d2e1b789fe0ed28d36fe5dd4fb3669;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef63d2a8591f86478ef65596b65be342e05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc93def9fa6fe003abb56e5f51f0ed59fc63;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f18b5656c6cdcd78105f768431063f2e3af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0262b28c06ffb1e454f47acac69ecf0eee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4244c706d904f68c681535f4e028da8dacde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20b2fa30d5027deb928b4ecfc8e07433be6b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c8430d8640e24666ab2cc4b9bcbf901ef07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b6e247e21cd1f8dfb89d9093a94c98a8de3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h22d77fcb7d27c1df094e22b71cfdbae3557d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf6044279f5e1c4442374aed742d89d53325;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf00dd6a235045523cd1cd55f7ac52f90cf2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1530c8af89ed7939b3b76b0882f0b805990;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44d9575b4df2ddb2d315dfd6e767a653e45f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91bc039f866209cbb684eb50b6b5e5d25844;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ea53d6b8f0881577fca9a1bb9328b59293a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b4c5c4f83cb508dd3fc53a35e4a2e318bc3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he57a3cfce0a9fbb36b555f2db453e32a74f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3d75003a31c6bf800ac6b098db6e37f47e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac9bd6fa485c846a9b13de5b8b98642746dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha52a3083dab010b735c98e37a4d7d5852ef0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a66cab50702115f94ebf83640c401db3059;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b9f755f504b0878dbb3c4ced27d54c8ef43;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had738bc44a820d250447047ed97bc24ff3c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14a783c11c6969926d5b00e4aec76916fe76;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1123630f05b674bafcc35913b3f95226ea2e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91d9d9a7ae8ae2f9791dfc4a40034b7dda69;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0c4e752aa3d9b6be8da1efd1b058932950c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h676fb8f00a28f86d773665906b0fb2f83c24;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac31a44e04054ae87802213fbd364d7e2ccd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a471b3694afb81058ac3f669426b952379f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82b217b49ed2a689c2f346ef7bd437c1a765;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27646bb2538f301db5e95c1bc83c20ff2ddd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h440199ab9ee0cff6f4ab01e960a64e7dc178;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h690a9aa6680defcd8505eda90b26b3b84d91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c31a796c2b5e4c0569d97b044bf98b2f15;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98876e85acfd3dce29fe5443c9313ae3e74d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8859d39fea22799954d37c6e27e787c33bac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91a596aaae7b37a6c3eb02a0c69ec65edcb1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14e601ea10cc87b546ec09b9684b5e88f727;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27c3f43dd1ca99b5f038c77887e7b961c3d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ad015b5c01658e7aa113e32a8db274db49b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h131f023e0b258d2cb228e5cf093d65e32b4a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5a468d290317e2f8665025ccce6a0772f29;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h983a6b3e71e08d6d2762c02538eddfff3b03;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6c323bc00811b0a734cd1f50cf45409d841;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9946e79d987c8a04573460c3b1668e6f1372;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f19171b69c4acd3c5cdc43f615fa954b775;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h969fd566f9e3cafa6a9ccf02c1ad86c5b834;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb931501faecac897615d471c6b13ac74955;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd0ee3fde4e046dd87884e95928e2ad24df1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haaafadf589a5f1fdbbe55c5b096d0c1c87bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f74ee894e0c75dbe9bedc28acd1b9c57974;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfa5e002e9154c78f1a3573417202aca5c99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbdd6e1b2f613765d55caf8f43d79437ddb1e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6049bc0812ef12c122830803e4d5f6047c26;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36db4497b2e1301ae722609beaba0a62e210;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd828226069ac981d78e6e62e6f4cd92a5d31;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c56b23a9fbda8caeec1035408f1b192080f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f4beb8427481d9d0e2f6b69f6a697eaa377;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1d4b5ece85d1ac8ba71ec118c52878c7205;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f7a218f9c9cf3b2d7f59f0e2374d0ea4d96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9568aa38c7fce1607a29ec793f8da953f82d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2949c59114cf3405c53340a20e82882940e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8646d5a4943cf1a7f15c24f3ba6d725406a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ba1bc9e4db8e150e76af35785ebdf661813;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83a226cfc451a03028b5ec5db40bd27c62aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc890fab5348671010320a6349fda2bd73daf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14afaa7100b60e100bd21a297783b762c521;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b7c76663f1d435eda3222cfc363d52c12dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b5539e521a205ca921e1c08c89469f3c2ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he778f9d3b75117af96e5c2cebeef5d08673d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafdaccf58cbc7717d385ffe967c5ba6c429e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74e662526d4acdee3587275df08808661a0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hddf3322dfecbac2b5e9c99992a2f26e8332e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e8747b043c2823f8c240b3f5ed585971af7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa9d761bc47e8983c16a7a5e34fc7881349d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60bd7abb01a107b9bbd00a1812da31d40903;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca298aad41ffe1ae0013600e99e936e7d780;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1fc2762359337bb69ad703276612aab0da54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfcd6fc005eba4bd6d37df812cb5967728698;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ac1577db3c32a30497b14246a3474319668;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfcd82b42b25be71fef0063bd42ddfda4a9d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1031c6cccea5d061ec4185a70974a2d32ceb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcec3a195cec8cb7700a63a52bd9ae258be59;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a0ff869fbd94ef4f3cdd0f4269c0f11c3f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9673d3e52550703a2f8d0b6bcf9d5ed0e012;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h32219937c6b0d8c6d7186a0fb4caee2360d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71e2af3760ecabe09037408cd67726a7c9da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60d70261121d459c5d5bdc7c6b9812247fbf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha15bee91a39f2c13f453e6a8769a52f3798c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a9d6a0db4f631cc2650828ed15ec0413702;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe3d323655f1606688715a911c865f36fa11;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a93c88d409c1421c1f8094970f146641482;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5eac7a1966f1b8e63c006461bb6020b24893;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf808cf80e749fbb1120f467fc03e98288382;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h750790286f19e3233b3f9a0460367413f900;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e20fd81b88110eb5061df2cd2f2cc069404;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8cdd2f3b8c32c1fefa23fc8d8f30eefb50d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf441829578be06a2787454e9fc2e85dbf37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2938a0562eb387c1947d00d2738e28e15b5a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ba49645f85e0040228cdab6a6b97f76ccc7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee1e98a5e58bf640b02c61679e92e51a9c0f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h745c6d4eee7d49843abaa574ffcb1cfb5126;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e0ee53ac05a3fb386049d71abec8f4e2166;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8da1f5841d466b2b84aafb8056bf36618c49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha994f3bbfeeaadae0bf886fd7cf3575574b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafb69419bf777e4f3cbddb2064970454a4a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cbf394cfeb4c1dc7ad6db7f4da9ac15135c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h582b1fa37bbc63401210f75c19bbdfa9209b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h253d21388b6b05850ddd4f2b1bfd6895958;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b1dd3c31725c3c841d5e09e975386087f22;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab59b2fac8cfab04231341ec669f6e90f17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb510f354ada6c73b7dd9cfbe780652c54850;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbdc7fea16de759a8dd849c1efbba7ef02e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7cbdf90f3e6656f33002ccf6297e153a80a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14df3aad8f59df690a5fce9f5c4b7629cb0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9362200407095947beb6da99d352c730b54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4473e49bc8e00e922cbe04b172a5d27db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9b23ff8885e546f2c4a67869c776cf25e75;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb53328ef59a6c6652a99af475c0549168c9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h644a74a64d9bc3f5094ecf276b4af6498822;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f4a21731a336abb35a471aa66d192ec693e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82ba58a90c83b857d33c19673c7e4a83ce37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h754c04e5d85037ca11ec2440b53067e74e7e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb450ecead148a850127bc4599336b21dd844;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a9c29b0e709d523da16565d521c715b0288;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hded8328b29206ef370b277eb0cdcd1ab6f61;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6d4ab96ce3b01ccebd148041db79d3563cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1771ecec05338f55d86c1b65c74f3878f2e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haea8a4c23a70df5f306d8a5b244360cb60e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd39c9d6a4f36799f25735b9eb58fc5df9a08;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1f5db2876d12969fb44a11cd013308758ad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd470198392dd1f553aa1611a71a0e0feb7e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bd21938d09a3ff061c41cddfd29ceb96e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49029972d7b4a99f288f44ae4924af7c4dd2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d8bdd2096019ae37940075d40c9b44e6d86;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha33f91df31a39702ba133da57a8660f28eaf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4532fecabfef91598ce5d672486745cdacac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69fcf6ba3cba45032c1ada1132df0af8817c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h859450a1290c85ba186650a1607f79ab4baf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h335c1a0635c1210ff67b57d504def5a41256;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68cebef1dbcd577635e41aa1768e181e6853;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76953fda7177409133c45f655b7ba844ec82;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha63c907bb0df121b366aab2ec704f1edc91d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42164bb2c021ce5648c07ad0e03f338b0f87;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf51d2af40172a6550e0179c06fc907ef450c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62bcd69a32dcb37948cdb7b70fd9de6ce3d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f2eab8c2da701b71ab0bb325474f386e06b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71225778a5ad5a40531ac2fc94320b4efa7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebb77ebee2e6fa0aceb28a98a713b596066a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1f55e9a59ec2b6d17d7460258b0d98d8668;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde48a3b6dd5e3c55fc0e3e48bd7a930a5f3a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h779fc5fdb8d06c086804910bce3abed53695;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d32c98b7e82a9e996318440c502660155a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87822f2070266eed606ab4c81b5e84285bd3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb00df820ceefa529da67b538bb0b802ad7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c777d5d84ab90e387e7fa866f1e0b0ab6a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4152091eb0b5d93d4d255246148bd878796d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3049b464f58d56550b71cdcfd198923f96aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha80cce62fe47e2ff5f1c99175a4952d120f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3f9a900d1fa2c42ec7a1f49a3f4a43882d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55a7ee96761ebc740bbb64e97db98d24e62f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3d0a21683887ff1737f49c3536d9e04e601;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1baece36a12e4320bfd63a7292b33c534dac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda1cf94707dcc1ad6dd938858ce275aa2d8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd91fbf1a7f5139f7fcc7ec409f7026282504;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha76b79d09422e068756f7ca938a12082db26;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ab28987a7469853aa24b31461a99f6a5910;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6074a08cf52be74affaebe44f5adaaf51641;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hceb3fe99e5f6ee6167896ab35bdbf9b10680;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h606375b50e37e43abbd8942e7c41f0e15630;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h942589cae322fb48bf97e6d458052a1461b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb50589a6cc3d13ffaf4bbcd2c5d789bf6694;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf433a4aba372f6e05c5452f0e5b61d787708;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha91f06655990efeddeef003ea574e64e13f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h32e757f1033e6682e68baf9e6da15162b455;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h641555ea51141ab6e1fcdfe7448d26897c8b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc40baacdc071a5ecf1d21629316b917f868;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb206c4711d08c50daa41b657bbe2ed856bd9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34330cc29a6a260955c0ca5c465d708d15c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h829c75db9dd72d545363c64d7c75bb4c68b4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c27ceaf022b919e4e36685f7f2df22ace30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b28c53fcae2a0bf0b48c01ab4703495d332;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1ed6ec1c6e435e7292500bf965baf36bb22;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfcc65df25151cee1b9db8652b63a09fcd02f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac68a81c128b0ec394ad2a1db0eadf98975e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7a3a21a181b3a638ad61e22e6318e1ddbb2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18bf8d40b7a6d2fa61107a73afd1213b2619;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8810f1bebd9256694a47982a8e010c8acb70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5425b81ea8eeb32a94e115d571801a6704f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a45dc753916fd50e2d9a3830efd4bf11bb4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3bb4a63988cf0e3de4d3fbf3e55abad9c723;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9147eb87ae28a786ff55840b822843ed7d43;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44fd3d628588aa74e2089421831ecdf41a9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4da3057a32b9f6856617b17f356e4cee525;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5395f8ddb73f3ea1b3c7c0879876cdbe2ac7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3264e58919b88447098e87117e0f884cbc82;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1c76fdd38df3a39416195caf89ecb66bc6b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9716e0b3863f42b0f57840c70406b933d665;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b0594a5c4f1134e7e6c63fcf83a4df0e30b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8469c4183254f2172796fbc27da894640184;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcccf413aee13ae030bd906f9dcc6a9f95431;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe0b939fdacea62095ea770ea46a731c61d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h41cd22b869b9fad334f8231f0aad7691c05c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf05df0a28e7335c9cec06038cf64eb2f0121;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50b001711de7075abc5dbbdf20d038e7e972;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3f99414d1addc080a732fc07cf2ee6a6dca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf06fa985e02ce4968d9acfb15030bff7714;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc27ebad66de71d5637d32ed0a0cd7f17f657;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15441936dc357b593cd4c65244fa2da107fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93661e73fffa47853354f4817b827b268b8a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43fe22be423f84b4e35682ec6d4396a4930a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8f1df8055b0966dc12244f0e37a3db3abf7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b9ad01249da2c18e55b06029db3b0c74010;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb158016fc8f0d579547f917ad4d59e5f181e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85249f6ac2c8f3c20e246dffb44984db99b4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h138610665a36af5176888b328cfc4912cba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf90ab284826080abbac9bbac2db52dbad218;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0b35d154402acfa06dbc9883b273136deed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc83e89df11a0f67326f63e03b62eee110592;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2edb350e59335039f7fb033e244a36805087;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7926145a6778122a40c3626fa058eef9a33d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9cd1fed7468f166e88ddb1dc6e2a030ae86;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf79a8da1d5ad0ac010f593af717c2c6184b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88f9492d68fc924eb8d70c3c69a90d285707;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e4bcd897ecbd758ca79ac87e872ab2ecf3e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2153e80afef35d80b47183dd73c54581160e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b0ca63171b0d2126fb7994d2a13aa5b01e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd30b56f7fc5a6060a3eba9f2730e89a3d84f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb82b06495d71aea280fb04fdb97929d20dcb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86b77ef80809b679fa826f046e7b142d8463;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ad7552c931be2048e19748eb9f530349aa0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc87ff1c44c91caa617d90ae3fa9523c95e13;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84797be1b810b1b5b73edeee0b1b4243ca16;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1021962f58192114d1dd2d1e6635b2d4f037;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4085a46572d7db62c0a366c32bd45ef2bb7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha15a8962efeb3115bd4e7ef78313d55658df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24478d1c4167a23d72041a58b62ff48a1e15;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b182dd597581d44a6630e9128e7aea2e390;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1e7af413095d6a1ca120e7b9e306793379e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab5b42ef343a164ee65f9302b2331dc3e72b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h870f207b69614871fdb6ac17f421c6a6f685;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3fe13fa2506d600a57680b6da1c48116d8c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2ada8293100efe8b4fcd4c57f3ea3044b5b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h461e118fd829065f3ec25778faaeb0414292;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hadb21f0f7c6422bb623fbd48c39f8a32c7d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb629989e2dba73f3b91b000b2a9a5b98083e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13451d6a35a3a99c10395468118587fe9c0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4229ad2c15f98f61f1d613596dbedd628c4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h782fe76c1697b9d21353d5c805e6ea8e51ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7231cad01ecdd9aaa6dabacdf55411253423;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40451f301ad0498cbcfb59906251cc069142;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2ae2066f6feb6b5701240b8ff8b85003461;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb964cd2175ed80c10a34874db7e223c472e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h304ec79bbefe3701e3c91a3641b51895111b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9a98d032418a386f9d4da23dee037c7d3f1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27889acb334801c0cd0a3d96ae5c5ab32ced;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50a46bb914bc5fa0d77b55eac442f5034c74;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb9da9d9cb9238a11e7a3caf77ff1b72c713;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4960bd25d69bb2522ebb4101a015a19e840;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68175df7bc6d9fc3109f20426b32fc07d31b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10a5fdcacfdbda55d12439a6b5463efc514;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h280fffc1bbcdd0654ce41548cff34d5bd015;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6bad0d357424bf1771078170da31b9c66ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h637c8fbb9dc56ce7d72a89930d674f9f9db3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70f53067ba74f812fb0e7844fb4f556273bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef6eb7e07646b800cd84e98267cf640b035d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfdda4af654e1fccc232fa53e96fadbe4db2a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91a1f961b24804e1e50c487ae9adb736478d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd37ba6672dffff364f88eecf804256aba9c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb5ff6ddd69d96053abe0a98c35de038551a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2da4116ec50666f7964d68d927318e4f866;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7833643f748401cf48571dc6af1093ea2528;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3886635f3d4ed367a7cfb4713cf9ab98cc84;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c056fbe380b9d1032508a7ca6a611ed8829;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h349dedbc4b3c993b1370a0f67205091418ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91f8cb6ce09cd33671f21ea6ac060b850caa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15853b75de8cebe66c697c90210c691d400f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc52e96a41a2edcbe38b77623a2ce164b0915;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h440a1b1011f1a8b181e43ed5ec0d27d844a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habf71148cf596e216ed79e1f3c131455d81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b6c85488c5f26078971328aad8450ab73d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0bd5364be90bf56dcfa667df6e9487be62c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88b7bfea75e2aa7e1ea59712ec8c2e2ebcd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f617fb86305d75b51adac6cb5314020688b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c3dcb20abe716a60f7d7e7889077c25e8f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2aad22f725d88ea2e45cff9cf6bc5c996eae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha3b8719ed5f6e2af4eee06a986be303e4573;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e6b657628d0dee5e912ca265df0d174cb2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd42ae211fe7db5553d45a5da52406719ae92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36c2542c2dfb8db7e1f287a811520228c812;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5843a3fbe27d4efd7871d1130c994422c1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f1ca19df94618bd042fb5661907a954fd7c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he17d35b5dcd42c746d0244310bcefbbaa291;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4be3e360022f8df92bec0ba9ab632620e1a5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdef149e5a0fe693e1a2de63280bfa4c73d8e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a31f3b7bf18969ac5582a3bbca5c7094920;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca20219ce922045c23b2e9ed120b9fa719da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbcaf885e1481beb8dd538409d9edc18aa22a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6df0230e6753677aa5c8136a69c2e19f92ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc338c5aec0877b0dd195335986519343d8a0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fc7072a26cc25a3fda92789e362c2e57163;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48170a1768a1caafa1afb9ce965f296c5361;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68a27f6e94c493ea32588c200e88bc1a4bec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c8e5a76a02a1086afc59d8f6a577fb11e7f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6501089b1024dece5c7b9aa1ceba3510152b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h555847ef4965db0763502a2af0cf461d1a1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43a9cb8ca54acad00f754d83255b75c53e88;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3215ee168cd577cd01e69b5180d7a87493d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9646691f77071f487c9b393cc1bbce9e8a64;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa03f16bbabcde81372436b368ea4868fe71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67403cffc31902e27333e19f5c899ba9a09c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52d17316ed57e8986f707cc13684e7609abc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1f8ad5c314a05f1de3d273e537f7d9d788b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he555b2179f5ffe8156edd901ab210f93f16d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8ceb47f9d0b7590bb55438b8320339ba340;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f7a98e93928c6a1fa6a89b7ebf6dce436e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33550425ee51f38f2cd402db9a8ebf9b195b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61a899f517cb64cb438bb2b3e46b9c39923e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda520b5cf66e0fe5c5c3524459e63c750d59;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ac2fafda6f611df858e4abd26afeefed68d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83ba7036e31a44e4010a1f6710d2398d81cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c988471aeba2e352d2ed4646aeb8caf5e6a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4adef8e8d81a00dab28ca58824ec460dc60a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7091317489bd99120d1e79ba9b8c8065cca3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc22201e9d725dea48a0d5c0e69f5c2b705b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4c996d1b324a8499c8eda73b209b51f06b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha50a061b12cb5569cd5c4b5f0ff0e087b2c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heef1de68a7761a0f86c5707132f9c4324ecf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6c082037827652d72a917c1cbb7db751546c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4217b4d121338462aabafb5e6e6d85f34720;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c76d05294de25805b781ee262990de6a8a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdac87a764300d94e4b83daa501f4b0c919de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf73e4f1b37e164de47f7eda7287713476014;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45c45b6387776c5676979f3a053d8e1e3f05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1cc0e59cd65514175d5cd3478efe47ad90e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80b71c545c8b810a8c7d78dea21dab6bdcc0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf620ef3c2ccb6e068132e28303f7c3be6c90;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34cdc2589a882b7f2c7e7da06c158d7fb4db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ba552e5843951295f77f0d656fe0c6e8ed0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a5fec1c08a8f0311bcf7b59a2a4f218eb43;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he81dff7d7c1690641e86c1255b76269fce95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc413a0f5be377fd2985f24e8009db23b733;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h107f9e241f810e4fb1bdde4cc9e08f7f8a77;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c7b4c28c2eed1f6ea66eeed1584a381c7af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafb48928786fa9d032265478302880dc1bee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf10ba5af18af449d180864381994f9d7a2b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc81d6c61bd22c271d7cfcff239b1dd10582d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef1dbe7e0010c6bebc7730fae90a129d729;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b4bf351a4b536383961a6be5f35203731ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc67d25221a49de06e736b6eacecb6dfd05d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b716b4d7350de5218725e2f25164fb93856;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d26fd98a8cb1786cb5895210e9a5986c2e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h568292f980c8816a7e63e59e31ecc163906;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95215d321033ff53091be7c43f41cb278957;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h731535348c43de02b9ebf1a2241aaa04a1d4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfe8442e4b4da048374cb45c0fc8f7bbc948;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe472b03afe5f9e8bcf849a0a6fec012d4ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0a0abd25807c9813460a3474ac4162630dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fea224a639c0dc03ebd724a3160d284cb59;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc346e124a15062b8a5d43aa790d6b2ca25db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d33b285d59f26443b3579cd33930f86e6df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h184fbf469ff948b36edb36e5c5bf580f21ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb57994f4b171ea2a5262fb0dde3082b423de;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94b4706e877e3b467dd776057e8fb8e32c25;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba0e1ef887c3b0375cdce8df7c44c14bc066;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10a57281c8a7dd9ca247c7b72ffd6bb5be48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4a0f5d081bbf780d19d1ae62dd9d1cbef7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5164738d663e85b7269e1528e2c94e2cd7a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6bccf3469bee5e5e04739a56c83c9cb5f5c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ace758bd43608d069eb1c1c98e1cd8af731;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11c1bb618a25e2c59087c64ed5dffc97b14a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h562d5ba957fa944447976d71b6f59149934e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6fbfc8aeec12beb154bf24e23a180a190fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf09d130cbd9967f31dfd531a363ca6058d7f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc173be7c5e3d12634427cc4b616004e85f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50a72b16759f18c62e30741433076232a2b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h156dc5fbf4ad3c54d527c26f23fbc8be815b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54d2c3bae1be4158800b99482b23615d1181;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc21cf8b2466b14daeb5215ab2a2817f224f9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54be02984aacf58937ff9a55174c67fd34f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90d709437781c36647d7ecae64bccd26c95d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbda597b708a623cd5fed85095e2b0c52e540;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b4c49e00aa278aaf7d9ec563f4d14fecb1d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65e43efe6934e38054ac61d9c676b7c6417d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h124038131c18e005b043b5f3fd831e205c98;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6c5b358847f0cb024bcfe762351d6de3970;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f52a194cee239794031e580a4afb5929b38;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17db4ae222870e419a656366dfa1ca2928f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20a44c063571ba2bb8c69e8c2fe17f1c926f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf76e3bbc5d77ac5216eaf10d4cf8f804fb4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0a141d869b27bbf3f14941cb125f693abfe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf5fd949f953a6a619d376e2c7398369175c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdaa1948030457ec8d88e999f888484cc9a5a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee8c555d93ec8d471d12df992d06a4347841;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc18e5e94e79b406830177abddcb886df76b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87ef5cdf464bb4097e0d7d492e4939627a52;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78af2b6a97aa15739eb6d83eabdd5fe1a1f5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90dcd69800500f4805e2c2fd4bee9dbb4837;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5a0ecd194193f14bb301aa757ae36f8a782;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e67274dea7671e419b9e8ed91dced33f4e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d93ef794069a19df65c69f535d101cf0e0b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98e570d544a34f992459f11d5ae9438190e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h213c577a3c1cdd9adf685026009ba54dbf8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3581fd9d88f19a5bf91700214b1b51d41c8d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf47d55cd60368ae0eef83129f89208a0d14;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6cbff56b8ac7c5595f851976476485a64abf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a4e3a65891582dc9eb1aa1fb37915d7a8ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20f9156faaf6ea78b284cd7c3a957baf83b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56c565fa0e5397132a73c4bf39720b51ce20;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1683f4e55080f6e1a86128f6f645c07564e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33ce2be78d281a9d5b5c6e306220c7bb011b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53d979b1b66543ef426deb27656b137a9c34;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3bc88bf98d457c4f1e24c0da36dd791da001;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca15adeec0a384ea2ef42f7a3df199d8dc9d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ecf0e0ffe6527e49bb1bd775195039ecb64;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73ac415deeb109eb716cbb2d505a4a998caa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd62bdc4a20849ec75d65f86841bb1a44d883;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b2c5ab9d5b0363eb46a6104c81d449c252e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83ccded14a22034e92514f00c5a1ae7c4c9d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91ac508fbb16a5a801a98dd597094a792bc9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69db7154106e679420df4f4e683da2a342e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f3a4f3d4e8dc981863fa536b2be9d5edf67;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he54a1568c441e5aff1be4c902f6d7611d3c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7eee4bacd88ca8b8f05b4628aa69bf0f1d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d2060885f33db04b9dca3f4e193e26ea62c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13fb8b3eda27983507d162caea2295327d8b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbf376b16b3af654304f2b8c2f65ca254ba0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hff8838cf75d9b6b67630c7ff24f0f6667c63;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ee6a37db006b2cbb6e6b968b082c2b0f26b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc141f816bb35bab4564c89c4d43470983d29;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha65c6d2dd400651b2cfdb86a3a0ecdfe20f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd90aa8ed0af9bf03c4dda4166f2bd32b851;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69aa6e702480917cf109be3c9332afb8ffec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc79d0a9da621c9fe37a48d711ed53fa263cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15a4f8c3260841749192848d833f53eb22d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63c7cf70d6f7968b9e051a65a9a8348001d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h521bd1a1a4f137958bed136fb352ce62f510;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5666f85ec58852743a6de1ba83aa904910a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7dcebd92547fcf03022c368d4023ff04a68d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h585298631f865bb86d188ba3df58c01e4608;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e26074af5ac00013469d7633e9977c5162d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38cd249b3cd82705c1baee857e0c6da81652;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h264160d2726a384cfa9cacfc1a3d600d1d65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9750179ec495c8b17c25abe7c6bfd3f5722d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0fd35027b3328a587077e6b14b107a9c170;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64472cec2c6590b393a377ce8dac4fc34eaa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5706d725eb8e8eebd544f5cf6d65d838d21e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37d0bc3aa5a8d706d42795315c236312d43c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19fe2cf3324f67f75167741f91155bcb996a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h562f88999a8b8022c384e2648c1c898bf47b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5583877cc1b820bdac4fe3360d3ac8f688;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe9b1397d0ea20cec95db18985d8050a1881;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8752767067113ded57c56a728c445583fc1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcbf735fb6d7355a4cf4fd50ada8fc612d238;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b49e320d86dfaad034a4814237528ed06fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e236cd511feafab6bec3f97c7884f085544;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90e76a36a9630a65a91288101c0848ea4ace;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb339fdb4c79854266a9881d39800edcf5709;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec5f8184f8f95193ccef15e385491adccf00;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3dd18c60da1a8e2b425c6cc9526267282b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97c31379bea49654f67b75a51d1bd5e92554;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44762a6d3d8933be510eaf21b1e43a96eec0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb864edc65ea2cd85270896a0ec2b4a28924e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0b8e3a4626fefb061f35b291bd7f8cffdce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52d5a8f8e7e1c1c06e97247051257b9301d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbea2f5f18c9025f4103b9b98ded4222b7ee0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h906f122786a8b8c525d3ab7cb6b146dbc17d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c48084a19fce84d318b3bdaaa5fcd54d3d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'head8726fad7863a1795719d37d52552c3f7d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85a589880e01a898f3f4de93e2d86d2bb80c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fcc1a9a5423aaed7b1815157396bfda7752;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haab61b9c13de746be627bbec0055c105fab0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf13abf80bd665c62f63c30578b2f37ce3756;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ccf64d56b4fe5146c2da80498945c98a03d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c4ec25f01fb443bc64743ce0d993aa48855;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5ac29bd87e977f68686656c2b994d5e6c80;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7d70dbdbb7cc46710f36038b2dbc3661f3f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d4117bd44ffbc6ea776dca85373dd7479b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81097f91391521dd8b252c8fb6be283ad4c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ed970a4e7930e50c8671dcb42c7fec68405;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbef27a8e9b23205bfc4eba25e7aaa3c0f49c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4bed8692bc6f73568f4c6dc98ea7fccb90e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f6d36bc0958b72c7840774b2579238002a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3349a0080404ed193fc47d1520390cbe5d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c31ddcf27140bd50c141dffea6e015bfcad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42f6ec0f88426f8d12c0a0f2fdba3fd4b70d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebb907882d0401d8e63b5bc8c35bc689d531;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ed233f3590b693a82be12f321a71f321104;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8dd5faa7166261c258ffa3996009b8075c1d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5485e09a253b1efe66cc1510bcfbb657907c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb68bce02e83a98ea93037b8373256bb5f07a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h71a77fa9b32923ecd0c8972853fc5c690e62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfabeadf0fef94860b31f7b1e926c2bf349f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9b6ce7abcece28559eba4873c622506c4bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55ad581c748ca78e25ed32415e97632d2a2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he2b68cf37d77a8e65427d97529ec519fe6f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3da058718cd0c822e3e2f4a10f2ced43171;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74157f7bbdd090b788ca36877e267c1aea10;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c6105638fa903589b87ce1d90c2dd48d3cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca0e1d1a46748321047b17050d63ee276499;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha00f95eb5011d909bdd40f60e2db279b57b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde530d0cccc08456b487895b45e05b7b4da4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4847a436fb4bbe4b839401a342df3b00780e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8d950e024ef709e230e13f55bfc7ffbe696;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc09fa1a4cdd12ea16d5b1ab5e0a50073a4fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15c7c94e1a59ea2711453e4ebd83ff0cb0ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e1a93ee7d822ca74a57976b1d9d03b0a7a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd658852c3b51ecb97884cfcf9d3467a2271f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2dae73b866fd73ef41f29ede45b189acf12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a7f0c75c8da4391f7e62daf21a17f9f02fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h653526baf8fca66ca5af2e62cd8229b72186;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb13e4bd7d488072d9f90602e537058041e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb69bb4e8968fe1e2851e090d8060be7600b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heef27a655d6162ba495a40f7d6c36db34785;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc3852692ff56ef2bc9e0f51b84995aa1882c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48b1caaa958fa7b1f0d9e35297a5008b348;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf629686055e68e76b1e12119af3cf6a2dce4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2dabe6308ed0756ec0cd4f3dd3b59e404244;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d5b7181b58137e29e7f7d81bdbe66f49f83;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52ff3c02fdb3c93656b5c13b915862c09575;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hada3e0582d1923826ef867b23dcb4ee52dcc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha09bdfad68736854954ce24f5bb690d7ee98;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80f78b7d5398d9faa92fa0913702261850dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ec5e27d68d6a9f3e0ebc6c1be6a501a354;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7c757e280fbfe9acbf8fc3a3d8a0c9f7910;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h23cc5fd0a2c8917c2d359e4e13239ce2681b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1be6adec20a9ee54885d6c8dee526aba2532;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc88ebe7e3144d94ca20b9b25badb9f23876;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e5041e1486c5e428fefaa0e31ec478b83b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfea6bf1cdc6fc7deb70b8d83b208ca0b283d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8aad06ccceeac215dbfa7a89ba463026f3c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c92658d15d30d6516e3dcf7f5c749762a07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8410d08acc61f5f83dec337170a8e91daf0f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc70fd641dc46c9263f5c1a66bed1e7f543bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2b462c044a77f8096d9d0fefc907eb25939;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h457a8a46cedbe52aa9fed1853de229718499;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3bb3a2ffe8f3b0095ba933736efa1762349a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9148f8eb586f7eecb2ab1bf5882783c179d1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a34de07b395c77678175ac84127001295c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb64be5d2aefa78f235bf77b1fea0071e7e66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50904a3ad32cabe935b0a7f32dcae1ec1e98;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52bbee2b6c1583b4a5fb1ada0adf0aaed616;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61ac521d1d3c7ece5009cf4af1a049537723;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9702853682c15054c2d7773ea16ea1aa6b74;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd316954b1722ce39eda65c20bb915bf686d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h857a8c7cc7137f1cf4b1603baacc4554ab27;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h456d9ba24c2d34dba62a88c096e0de4c18db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2eec0301d0f20045e97854c8582fb27f0b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8fea29ea1d69f7b11062755415b14bc54a22;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha997af6748b42befa71270b9b9264089610;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4148ea14bcee75d9d5944ca3edee0628aa42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h719b490c48a12ed2f1172c13507e41294755;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf4fe9f84c84a87811b867331660ed77d5952;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda84f6a4cf3162a820843c91ccaa9a5bfc24;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e0a17da50047f393c243939f4b1739c9611;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62cd927670dfd3b11980fbc1666dbfdd53ba;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h900d3cfc89dbcbe9e2900972bf1dd1d688cb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0266248480336ff4ac5472ac73318b8f3d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h180e418e669d09b32469c5e1706444e8cbf7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5299a64436fbe1ef509b1f6db84a8783213b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59121bf3677628d5fd1a21a2567f4afc049e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h371ceaecf06deb0959c8ca066b772bef7ebc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h800ca776bbafef0871eb71e862ab924033aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6457db60ef8e8eb52c048ca0623ad21958d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d5831d1d8bacf6c01d244481a6bc6733c9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he318805aa14dc37cfdf8aab4df12ee349e2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7f51fb6bef343c905f9303d712730f02991;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd12d16e98f738c662901fc1e09d2606574d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb9331c448176f5b06a63e28fcb7cad8a335d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67a8694f65734a0766198cab3a1642722af0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3300d08308a96d9e9c709dc4e0bd3ea6b89d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbede4fd7709710c7e073aa6a302d015c910;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbffdda2386bf4ad03fc117d71ec76161b32f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde5892d8899735f87329b82f9fcd5a54686;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2af6de8565e2d98fd63be62769601a900e70;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3b0ff14fd555b96ddc2b163687940806e8b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a3f20aeb6fcd048ec35e5b39eff0cd68c42;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bd3f39cd56f77962abc217bd4ac098e00f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdaa09f50af22cb03eae3beaa0b4d34f2862e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ea0b134fd2e4b3a8fd3171b25ee21203df9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7a037b2bd3c4881db6362f6b75e8ff85056;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef7a906d450d2baf82f184f2c672d6f6ee43;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3fa8fb372136e7c437e93b9fcfcaa95f9237;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b34192ac5a4a62e5bebf180006f334b02f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb64995dd39ae9c7455c475dcac39df10a127;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7e65094593e542a249b7db78b178f651e8b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68c2a089b49dc08f96598c6ef1ea7f979075;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab66b281843363c0e1c8d7c42c75942158e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3fd0b4cdf3edf9aff91e960877b7d47e0d62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd82aa1c9881bf5757142ade62f86b4b7eb71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha806f423bac9fb286c65ef84e62494877ca4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42813b92f83f78337a68b325199a4bd32395;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8de708384baada63b9851e821e35d30e7b4b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hecdd57676d6b302d86293ea37a6cb6b3b011;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h819e3adad2f022b2a28030391d26792ceaf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe2c2e8edb1cb2088bac40cc2499db1dbfb5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h418a9c5ee668c3cc2be87ac569a651466eca;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf054bec71e5583cba854db2797b446bc118b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bc1d80300bb584bbeb22db83a17b529ddea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6a01289bbcc1312754fc5a8265ec6befdb0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f2de54a86a2ab410575cf2165a085156971;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h417f467b532a7b25e6c3ba7475bf5256a6eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56311dde0c578ff7266df71f0b3ec4d423d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4fa4c4adcf4a0f66855057c25c38538799;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e32c26eb283e6142a832cbbe1c3acd4a919;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc1d3636373e30f9e1ce827b13ec126fcbe6c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa9bcac6c042f10664c6f748721243e547a3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e488f9387eae4bdb03c9db142640551e1d2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebde64c46a1ecf7873b77ee72178ba98dcf6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4932ee079512b205e737d6d814ae5b6979dd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b77dcd75661002304bbd8fc78ccf0242457;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0ee2092e1cd2a74280a7faf21f0d6ef8dd7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60ab976466debdf3f5daf70dc0c0d3d69d0d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7b96793035ae4871c7fc4d947486396065;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf04557de5e8b4d111178cfdf4d1b16512bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb13e06fe3b5cc42325288c27c10a65a33959;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1f52dc75d47319aca318e994ee5e86d99b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ca00bc1a73bfa70a4891357f67861c674ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h51983698bfd956b044fcf1c127e2c377e609;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfadd291c8c691492746cc0821355c756c301;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h495adf17ea4e9a10f417b4dea51a17dbad0f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28f378addbcfdcf2917f21fc283d19d74b19;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h487a73e4b854f626d097c5008fffad5df8fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea3722c31defb85546519dd84fbcba5028e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37409f8358daaae84b69830d0e5aa26323ff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93e0574422bc537c0011f2f3c9e42d0a4e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5d1597422ae63a3126ff42cf7214dc9ab5f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2db19d474e7314e3aee0e3bb217c4eabc88b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cf7316eb4cfc837f0840cb49d00970ea275;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ac912c47973db7eceb916c69d7823a25bb8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ff7a9b26373a7240cb0cbedc71d674af41c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd361a0113c0da005d88260c1161a229f5bc0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d29a152464b42d68aca6f9b2c941317d0cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ece4e8498cc7481d678405822b71e675d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b487be0cbbdae2453b8035e749ab4d1a0e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf060b59f330d7d32ee752c5cefe585f5f2e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9385be7111cbdbd4d577cb91478043ba1e3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d1819a037e427657d7c21939721ce55cf71;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h731ece9ab1d76e61888a5d8d4c666a0b59c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6391477d6f12165b172408fd4e7d381fc8ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4aa2754f148d3d8d6aba8890f2bacc0b193;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7af8941871793764f47645e35e629f29bda6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h930beea1ddeb73b6ee6d4d7040abfd57ffa1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40a64835da84f0a1d68e2292c2c687b2b206;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f61826179678bda399da86c6ea9be7979e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6aaff8005e4387203dbf669c399b98da5d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h450179918413f72e4fae54a4348de2236a40;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93dc22d260d6a2eeaded04bbd8cf2e351de5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16fd023ada20562aa6edc2529e906408c85e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68d4275de66bb87165617752720ca9df2dd8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h483fcbb9b1e80caeeda76ff52b926c29465f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ec5b780751df0b86197f6c4a25d0cab3db2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7665925ef178c5a7cd9e672bd8246fa1d6f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4ab4107b0056556d25d17a1ce43bb8b85a9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87f9a398cb245df24299207925736969497b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61d08163f7e3995cca2fb01d337e9a01bd17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29c2318f2b35e5fece0b9188930459feaa98;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he93b7c5b316cd72f70a52d2e57d06cf8f40c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a5d514085d7239bff02d150a5192c8e0b6f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2bde3d41c5cc8a721d115d308df05022fcda;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fd1c3d5b962f8d5659d4924fa032e0c4613;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a0272296473af33ea3aea6db0a9c8bdba2b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7e6b5715fab284ad55d156700dce3f797c2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb5fd33c87f204dff846862a4ba8bb388005;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9279d9e06a9fa61f17114ad179f2cc122967;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9df40f01f1a260a3f393dd0c1ddf5b72c07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9ecb6a4bd3049951968ea65238b12e6ea1b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h904a89e5f2b9df7e2d2077be985e5aeb2786;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8560fd0e6c493b4d597cf40f82793c8d355a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0a75ea65681500b6b0c9403fbcbe375eeb9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b579c54bf5a0978854b4a6ad6b64e48f751;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hced08b63ed7f90b4b2b64b56b8c916ec9e06;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbf97c5f8baeafe2a4f4ab7b3831f73cbac4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5ed740d9dd549176da54adea5ae14f64891;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4bca4f9cd0fb49a9431a607f1c9beee6adaf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d8b34d501e60d17990b6bc69dd740679ad9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce4c37760f8163529398b41271a37b4d990;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f0c671cf12c85bab268f65f0625665f3dd6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e3e0633529fe193e3185333afb06a4a255a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha96a9ceb58605e5ae6f6b545c915fe9714d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb90e17cc4d6f6528cf46262f52e1f8db74e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c0dce5690b814b5c0033c1003f0edf5c42b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ee8741eaaeb33f11c02304a1b43ab335d0d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habbbfd79b87a8e69b47388b05dcfe059ecc1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7590ac25812410f4b0a6269075c9d3f714cc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cd2059081311bfbc0240040a67a68843312;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h877d04ef900b6da46990df829f07a7012f92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b74b95de8d9cf685925e4d3b56282fcdd67;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35c671e1e87a9fe6b7b5e83686f1889ece21;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce58b73085c2dce27cde55492db0d382c9e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a2cae55d1b7f87c2347d736efa689ec3d05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fcdce4558a3b5282d7eff7067c82578cb99;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90f88ea0420f06036ab57415affbaa5932e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ffff0847ee0ee0e3a98c339cdfaa4711c17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha582a7935fa8237610dc79ed68c4323c5e57;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8a4c7ee941daf867c9cab757d80c49b0f95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a5ea4eeca740ac1478e88c522d24fae13af;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f5f4e4cba06ff3da280be9a1413459cdd9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91b859fce4f7f8d6d1371db4c8220603f836;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1099ece91ae9ed740e847843e9ca5cccd38b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5ed2feb9b321d29852c3f4983e8cf6ded1a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2435746119adfbb59fdcfe170eec83055243;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc37be63e9353d2d56e28efacffcfe59e5c55;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe07d92acaf4c3b60cd144e43f002841f252;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d0c69a74dd43ca6b25f91d7730a2135727d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e48cdb883c0a07694aa5b1687bd40459656;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90c3a5a8c2f7b4f2b10316567b548a47c7e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd0c64ad1ab8085cae0917ebe971a8c5c2e74;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7cb28a7541c6e7ab1923c5f77864f309e2e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba9d931ecf38540e39f6eaa7ca881494049d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4bafec9e4b1d5445d5f9feba5205300587fe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2345c8107118ec98654ca93b4c1ab3d55e3e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69bf0c6c716c36487623420eec7c64299480;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1b67997f2a78ae5e705cd70793e0955a436;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6402bed1143a668ee6cc84edadbfc4e55c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha913017f679cd22ed4f0472868898ca6aa79;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcafc06aed9adf917f562251cbc6ba2a97ea6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0c862f15fec1c48da01528d26850bc2a441;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81c2937b7c932b3a8aed8c25a6ecc93322f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39873e225e4ed96e3cfc6372e195a128b968;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8515a141e493a7331e46ad7997d402701f0d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67551c065f0c1b84e59864f4aabe9f4cbf8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha2ed49bf5c9c1226e3105afa005bf5cb25cf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0a4985e6653dbb1ae290a17b2eec06e3d78;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7240b8198e81fbdf48621b692decdfffee8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7811c04d9ee7116a4ebcbf5b0e91b142df79;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4cf57463c838822c58255f5a87472b41f6d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65e4370127ca0506c83344170e948ef76d37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h907d5f155005cf04a0c441c1014f1ea41d52;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5692ad0bee51282dccefd32aed64814614d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd31f6ffabf998f7f1c89da01ff09f6b8eb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha493fcc6d2f5a6e86be169d9fa33ed783b1a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb541d6241ea11e592d378127a2f306659f3e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebae2906481ebacd97e1335d8b98baaf6d68;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h651726d8d80ae3a7461c0b3aa39ec33114c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fe35ddf672ec352b4cb3e641bc6f8915bf2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc575997725b36520c2d8b1f7a479f274940b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb67828665c33cc74647a258ad233dc91b1a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc8fe96f600cfa5a84a39f9ddb89497f1b83;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h436dcfa40eb2353dc0bbcce46ce47041198f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6769b91383976e895ef5dcc15cb4924a9e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6315283366ae7187cb3e9bbc8693b5ea07b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70aee308e8d98149f60cb4bb772a9252f80d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74aca42315703961f0d5872a73acb33f90c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc986d1bebb0c19d6aa5c3e112a6ea1c1b006;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2e93fd66217ff5dc5d8fe0bffb50f0de0e7c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf62a99a1d800829e86048a38804a7c4aa4f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf22738c8a746fccd31f1293cfbfb1fe29f52;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48a6bde4d353033e1fbc7a1b368ca7dd3e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1d0b75e1201761df500fcd3091f72554631;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4faea94e76ffbc4974beb0a1138917105e05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5979fdbdc88259963e499f43f9c9a80a5d51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec6e86f04e72ff746ede772d644411a6c038;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h197cfe8f95277e46cc3e2ab5baf7a995429e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h619e70093575befc1827a758398960e1287;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h399259f5dd331cd2b851fdb98f0eb30cdd72;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf25246ca88c5de9ee9fbd2a7aeaf753b258;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h279d72ba660e317bcf282d5556d8caa947f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf5bab2e3f67b434f77a794ca81ab651db50;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8736e07fd3b33dfbf0e584ec28e0f242e140;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9511b4c941d65b6744645b975f0e2d13cd9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdbda0bc0ef5a8b1a52404d2dc5c59c24583d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9b0308e1da221b3cdcc16b9f519bdfe4229;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e546660e4005210da2989399340e3ad9e55;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he29938f0b346d5a51f4926644ad89eb4e645;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc75dbda00b75c35e129b7e7c57d21639976b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hccb29e94a9428a7e066e7d0da7d97e6d466d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ba05f9d57661b1a330c6fd79136d3546118;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36ffde74aec1429613ee0cfe06ce429661a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee29fef24fdf9e421782cffdf57606f112cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a56218be319d11ef623b1791eba8612d04f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef57c0ce9d6d15d94cdfcb75932fd67ae25e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1673f465b973d82c065e694bf6d70964df08;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2cc4860e36c77fffb807787319fcfb8a177c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6bd4a66bd48ce085fafe16dec111fa3f3097;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84184385241311fbec7af25238d629df194d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68072ef8b5ef8b8e0acf73263569c4f98208;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b3bfcc25ffefeadd0773dc307a38c7775f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he982aa3403fdec9da488c8fcf9ac2b0eacf9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb2914bdfd3e85413e3d0dcc0d4f4906e796;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h448c514c73df80ec1246dd503bc2a0c7aa13;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64cfbd1106b00e88ffd30ada458f7a65ffd0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h192ef8b5259c78c5bfdfa968d0648abc4a32;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ecdcb2d1f6ed34130eba8e92834cb872afb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfec183839f99e2dd0c030ebbbdac22cdd6a6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8edbd08b08924b6ac892564c37f1a032783e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h838576a7a6967f2587bb828c00db5b077767;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73a41e6162e4124fe263f52a897266782613;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96de85f8b9bf3608a26d887fb6d34a0ac10f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf980ae06b3c581805f78fb0d849f85446d8b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ee1531d161fdb7445db8fc1b62c39f3a0ac;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc0cba8b07cd9402f9dbcefc71932c5b06c5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h540abebe61e5de122af63ec221b23628323;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he03c054dbf5a7cfae06c97730fc278a7a6fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5c5acec899d0a11bb948cea670f4348fca51;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7b629d1c36c78054dba838b4979f28e0030;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b460792d9900b4c531fb1e2b34fbe2c019;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he18524056acf7df1d809c53be4d149636767;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8dd78f9ec55c2e63d90e606d670cca7e711e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he6219700ad5160630e1862e4f15b27fd4bc9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37f7ad71f72d1db4ad633dbdb3832ffd2755;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8db0ffdab6a0d6fd74c008ba1636517ba4f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1170b0b9c019754489b2abcfa15105de9bf5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9c224142c754c70cf7286524786263e69c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7ad92381290d74cbd488a0cfa3e66460474;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11e9041695f61f63824d85efcfa62d00d0a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28bb82e5998091c9c1c4ebddad9451308476;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha26829d87ea70af3526d04f339bcd7824d83;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc27fd6265480016657e3cb600595ad42d735;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he60c62210e75e1eace61c71a5740af6b676a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c42c18af3bf330ae8bc5efc33fe8bef6862;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1eb97317d4b5c2f819664b319db1b055278;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ab240905d453815c78da01cbbf50e3eb291;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2c64532d4fc2ecca7a1eb3c59135d34eda1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16c4c5cad3cc5f7cb78912fcfa8c72da95aa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68c7d11706c736fe8bd999064cebeee32ad7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9cde08b96fbfb2e9ba2fd552fc2ba54a0c8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ee69892fc8e84e36dd75bfc34db59ff54d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68faeb3b71eae3edcdec96ca9727447c2447;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd98398a3e76afd357d0954918385b08d59e8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d1c93242fe552c441896f5f60fda7e0759f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46ed9ffb6c1474bf06d3bd7840837189c742;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77c5887053cfcb6250ef1b66e718943a99f7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8f9189edf2b0e1e3d634d714a99feae1581;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb68c65a9cae76d7a62bc744b75cdff209a64;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h798c5c6b4eab21b73dc38b24c23b4de5de92;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfec5325461b42bc5199ce19d18091f15f64d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62eb308931fdf7539c4e5e28546853a189f6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ccd09097568cd1d6a9cfa4f7e9cadf8ed07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e8c0f2c75a92bdb789cd9ecf6120478a665;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he52306fd25bae67115a0a7f1509c78c0d386;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he840c711216f64134c479f65da260bc4c681;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75fef9de66b518f7973446ec989296215da2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he0d70cabed5f927f954f0e98f076d37975c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34c250ef8467951d697d5980178aff4a86d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3dec3b63cc1b0a3bb7cef322ddc79c5374c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e79809af286e71d13d8cc7b64ab59517613;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84e6a6bd7497b75c64e193e341e504b66dd6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48b083b829ce2befb063f6e8be29e4a28909;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce3f5c585297377b5323c5886db00f0cdc61;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58dc80492c5df1ad94e024131f7711331571;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8295d6093735f0fe97d09862884295c9eb6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha194fd82187ec7988c375ae245b5a20786f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcbfca6675b7fe16ebd75dfca9bdbf9513708;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6ccb1c50a9f0631b01fdc22f58b42987893;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8b1c05acb93e48e6c4625ac2632ebd89f07;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9040279be43daf9a6507ac6dc88b0708f733;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78a68520d24f4fb2ebb6ef4e5014c31b44e5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4bcf7118c2b9dd7336b9a273370cf9f2de49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb497bad697dfe83a58a23e26757eb0ea47d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f5726a244f53b229be2920841c3dbc5320;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5db45282ce4c1ebeab37e56c76fe47e45d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha563597870b7fab9bba2c7df2d9e7e9c8df5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f039c328c45eb3a8dffcf3e8226cf9e6986;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83dff06dc640f53bbabc8b0f36dabeb5a44c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b13cb34984b96d3df5a73d843c19e799c1a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6137196caf133c97fa21bfc3e46e45d4afc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4af09de7f43e6af03c4b8bbc780d9381c1ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdda69e63f8d2e3786455e1c8321ae0f0a026;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebde5b48666dd878a05941df18c436986cb2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8b68ec7a348da5c6e03dfbf6503d7ee41b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ed20d244bac7c57a53c3238b7c7b0401f63;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4799e672881cc5a974ac59f8370836a04499;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha83a9e32f9721e7b277aaf78a37421f6eca3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc1ff0e0c16e85329c8f82ad8536abe0205;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc19d8622369e6b733b0fdbad5c7decf6908f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5d172d4b993585a5818bd7d319666b830ce3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfbea777c57295ed1a0331b483d8782288e9b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h79c06807dc5c5c3e469e134547c2a0d5e33d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25a29ed980aeef08691dc29bbcd594be5cdb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ec44f7a81b59dc952411a1fa29676362926;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc75a7a8e75e404ad62636878100950952054;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had167b12274498a110e24f2d76bfce3e5590;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb658f323e456053d3c916b2ab3f1d68b5acf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bd63405e20d61f7ab8a752fd25d1ca76ac1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf8876b5cae8c4bc86f48d7d48d129e0b27e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h200e5fda80f72d245dc3794112ee873f8ee;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb690eeb900033d4cc86b1d90d6ad4dc3685;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca718b9c7c2933c2a08a50955b4327303864;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3126c345508d3a2f8cf147c39791cdace219;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac30c24e45facbe5181d2aeb66c4599642d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab8ba36e46d3e9b0edc247322a6252d0f045;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e4ecd953150a0513a02811d32bf7d2c6b66;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a1bdf529b644a5a7186ca65a490040f4510;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha385178518a4c964857475202bcc5cff7db8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha39dc69453130146eba1644f4eaeb870a670;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ba564bdf2cb3f6cc54f6f497ddcfed1ab0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d708396154e0a5126c31124b155fc08f285;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h150a61d23b5740980fe630d252caab88d5c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h616034cca2db9606b8080c45c91d8e9aab01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hedaee7ecf9b773a3da3e914dd49accd0575b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h12485cf2b9f6432588aaa5e74aea9a1908a1;
        #1
        $finish();
    end
endmodule
