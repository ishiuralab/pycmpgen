module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [21:0] src23;
    reg [20:0] src24;
    reg [19:0] src25;
    reg [18:0] src26;
    reg [17:0] src27;
    reg [16:0] src28;
    reg [15:0] src29;
    reg [14:0] src30;
    reg [13:0] src31;
    reg [12:0] src32;
    reg [11:0] src33;
    reg [10:0] src34;
    reg [9:0] src35;
    reg [8:0] src36;
    reg [7:0] src37;
    reg [6:0] src38;
    reg [5:0] src39;
    reg [4:0] src40;
    reg [3:0] src41;
    reg [2:0] src42;
    reg [1:0] src43;
    reg [0:0] src44;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [45:0] srcsum;
    wire [45:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3])<<41) + ((src42[0] + src42[1] + src42[2])<<42) + ((src43[0] + src43[1])<<43) + ((src44[0])<<44);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa9ae58e8421d8e7a79fec3a11aa5bdb02b73c24b45ce98a2986b1de6b35c63e0b7b156cde095a02be9045ca62c0c9b77bc6d6ee16109c94cc28e95857fb86b8b1ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h69d9c3961ebea08222df6a863666d3b07db3cd6f9201a22113acccdd049daa1f9df7c1342d142dee263a1fd5caf67f227e9b13abf493895460740c99a6dfb2bda763;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e2f7901cc0c9498d7dd2b3304befe101dae8d5bacd1abfb8d723c1da072e0ed8383ea3457244052b0721d10a37d4bc71211fa5ef4ed7067822ec5b3e2a89a19ffcf6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19241235d7f80dcd646344e66e0524dd7b27d81bfd14bcc621f0c46272c340b03b2fe0c0e87ab895d130add390da2f06091ac82e575e337768e03fb0896d435dc4e5e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4dc717c3d7770ccb2fb60b380637225a763d702d2c3129aed3680fb4c737c7bf4b5601befbc4043e6e19492de03046a91d3f518847cb14b0df416f399b48716fb07a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e4a58b157b9351454bf93ebe4e8ef23014a44ec6b7d76a650a79f6349039df3d3dfb6383f061f77bc627fcd8cce77a9b63a371f1e56e45ad873a5cc7a1c48bf9dbc6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8cb12252114e2412bd3e9ad89664f9698187415ae4e9e539c22af471257b15332c3ca47c2454a9c507d64d011b20372e471f33aaf4e97bcda4b5c1c06123e9ef9a0e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h50ee2905b56633bdd705114bde493cce778b577c657f11f4c1ec6bb25396b6fcaee515ba744c201473bbd78ad03cca142d9e8a2cc1a090a47ab824319a6c714548e9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161b1daeab4d225e8da5059a050514d51dec3e9c0f18bdda40822ef00a50b9d17225fff36ffcc41d7fcdb8be493b6a7b787dd8a95d77295b8c997084c560568b2b8ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1df0ac2e5e8c42f2b1254cb13198abeac455d27046a9d93a50859b1b4e0958063d3ae347d52e4f9cfd8a727af92e7a94001adaedd753e62c777e7a3359a6d5669b1ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a13b758b9599d430808c6ee1f1e4ce1e1a7926fd9be7e9420e1ab1981845c6d224e3dd5977451bf873918198f72b6a1ab5b234cf4b1cdba507eb384e2969715c03e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e1dab51f5c0ba783c1aeb7f0af27d1f49f6c21a58c595910a6dbed50a62b394e20a4d9a08453cace310e3bae4a518ecf3dde2368ae9f0b24349267449f48231a66ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e45f8b802a419b6021c100642a57f97df22cd39bb3daec31ff938bdf7ff6ecc1b689097c5ae6af6e5c51fb8189a271d92752dd70a28de7facdd94dfaca9576838841;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e24510ea2fafb18e678cfa6ecb69abde1033992246463368d2985bdadc11754ec76f983421eedf14a7ba4349441f6fa96bd14d7adc04c1d8952b2621f35c54b6ac05;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c3aac81771cec576aff655853fd146794faeec45936cd40bbcd72667e112309ce4bb604c081812b20c709cc32449197fae79179764c25ca1557c7f27bfac6c6680dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h47f371797f3db1472c14c5aaa7dfc8fe404f2fe198a4f142754ce60f47b0f56aa5259776ab3dafe253032c07d7ca83d70e6a01ec83a62992540ebc932bccc3d37f86;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf79e660dbc3ac824f7310e6978cb2af480dc204a7cf2fcfc9cbc5e18000390d16f1566b05ca047c19955b71f669e1bbe9ec6ca859cb61dc131bc6949fdf8f303097;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193cc813e77f9aac49b68a4fca085fc64b0c1f2448aea22879da42497fa3e5f0c2ab0d61f1f3b8a8b61d0b348ea531651da5013413e0a911b5db3d77f658b6b3c28e1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d8c2f26958c755c91497fe1d73f8a3f120e0f6fcdbcf2ee4ea394861ac0872bcf2a64e41d5a2f2eaefb1d1764fd17b68b60735fc797e390cc673ee2ecf049bdef088;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha4ebcd4595532c3e9641543c91286afed805ac335fa071d21d9be4996169d79fef5d59c03a3898a793748332d7167b6bb3c056c8b4c3b7c427c59db5d2374ba31095;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6cdd20f615a837eca4fdb0d5dd9a082620605ea3fefee6c2447a77af2a04fd1aac5368b7cedf4e65f55014e4d96da613bcc52141eaebb21d48b533ad17f95db52e8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e015235a736717fa7219fdd66ac09022d143c07119ff10959263ef6fd76c33e96451b916067b4321f88fa054ed80092333cb50dbb3b4c7301947790e958ed173ced4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12365fc3edd546d54870f55d1daa0b068969c56292597426203d8421680f399ccb6873ee863286a851c45785f413dda5c7038ae1eae1899d907f58f9da653904f0c58;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e97d3fa38455f3c55669c9131b47829bc1b3b543c164766526e8d1df8047bd9a28b2503d285c4fae4d645858e198fb46337e6daedaae6974e475e837ee12d8103f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f873d42b3084756827b728131aa4b29023f894f609fbe4f26dc9abc69d7f0404587eeee16fa67073f34a940164b19421fe0418b99c8ed46b0b228d63f922da3bcb6e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3d711aa15283929781b07b8f257bbc9c53818992b55b271377da876f806be28670d05257f3c2db1f09586ebcf8752bd14f1a9e946e955a386303e2b8f62282fd4126;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10d8ced3b9bfe6913900cf02077ac3942e1d78d6c6fce2499592f4315eeb14ed3bd50084999352a1912ccfaaf3ecf9f9ffe4345be736ed3992930d684cd5df5e0b74f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd07c043d69cca8d831d63f42e7b65e89092aea86280120dbeefe1a2ccd914f8240b780bb23a0be87519908c5909ffb0429690e3d9d705ffbeb91ff05b2dec91dffb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fccb26e8476186cb0ecb019e0c6de2f9447a722bb00da28d42a6dca213ba551999d024eaee7339c8a484d9c875e944e74a0e2645be13bf17d9a7bef2206e648f0c93;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cfd8583fb6a85b85a6b626cbcc9c3b3f11e4770d98ba3baf5af0918aa971d4d32d9d09fd6abc062ecaabfc2530350e63d7b596c41f8e29131b68653d301abdd768b9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e5e5344ac6064feef60b5b06ab2db84a10172204a83e7994da90eb5be98f78fd8b561ecb363e9d7f533a348721be5dbbe75832d1e015f24131a0b3163ee1c2d50ed1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7a423f496da79d321ab08b5d1ca9769d9fcdc8e2929a48cebb792ef17776b4dae25ff41a6e0ad11c61a8c937d97622b90fae062e28ba05bbdc724278c537f146679;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13e34799a8d9b398d1d1a76bf2441f6efcc4a04038c1b8577ab2f2c9053452d8488df5dc8a426387ea58c006f7d4031b68153ba0938347d9616bc64cc36bc13963e66;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d6a576b416c956fed3f3105d47a120a24735ac1653798b3bd542734aedab3ab51bd4544a19d8f38c5df1858e544463e0f401766d44a1bae95f05c845cd1c1feb2f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac285be6e2dd905558f76d7376625e53b71aa440f843bd3666e9baf53af47852913c31dbd04304ca016c9695dc281cf6fa029b534aaa2e604a87e071770ff039e94c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbc475b913fdd03ee0b181e6808a43d2ad2a7802453cd351c93449251ee54c6d9ae884bb738ecd957d5a93e3fbf0079bf20355a5f9f2830b028805fb74000099c095a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbedbf86d50df1129898c76a4d82f31aa7fc09cc8d1a5d617bcd43b5ad9b3ffbf6e170906f3bcde07556d4df28300fccd35f6056854a2471049fd8236e64885ead323;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3aec2cfe58f4640ba43211bf7a1ddbfaa174ded9f5cf9f2178aa3eece5f133bb799ce2ae3cadecbc3fd070e736377ab4a6fad0eb7eba64709e987b6bf39cf13fa3d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5f4055fa3b15242c433c09958ca83a4d2bd77fec424f1a5c71966f4e02a7ec1391f8b60e999b8777855d6104a7f60b70e9143e067323b784d3141661daac04622a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1536133acbbb4c425542c59915ff68036bf2d62aa1548de8267726b805d5e5e33e92694cc2b0a25bfff73d8f18f97ba7687fa39f2c6b90f6cfe85375ebc879817a982;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5a2ff0d6a95e81729f0135d527119858e262ac217242508660aaff1764eea1bf1318212021d266baad242c4b3a1758bae5b46e8eebdbdbe6855296f13487f4d78b12;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfaf7c0c20aa4d0f116e5379231e8ac58cb5c63ac8159e246becd0b347e796c752b53a31fc6faadbc8b6cba871d508d86dbe5547ddcf0ff03da87e19c4ad4e14dfd01;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5aa9dcd7dbb042b38d42011328b4f667cdf12b7c46b5756de442fa489b1edcf414c4bbe519c96037e3051d7a2ec03275c8de380dd3c89172a6615183864dc4fe0b60;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd61bf72f4a572b8a004ee3e785a476b98dc4dde8476e833af4636f8f6d60400c2eb8ecc412fc6d7e419b53c38584e122520dc70043fbf4aa4f5f671cc2c52d270dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f67e856f3e5ce22a8254c614d0b81c6142c258f3743cd9784cd5948776a460570526044ddd20163d0d8232fb1be1f611dca72b137b7422b0e665af3b46f84150a9a2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27e52798792e01006fbb26380f3f480285269db2aedf52a00098cb00bf9fde8bff7ccad4c46f89e5062b65b0da5d3b54fbc55b4f0c425fb18a22ff4c8cb96d907fff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb33799fb197b242e206fa2f2c26d398a9abe7b0c5f269dd99b87113dd91e3146c9a36d388c8a5539a1ed8e0f84a1135e014e1435e19ff5d67927d86ab6659a7380b5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c6f25941569df4a7006d8c616aa83fccd4272a8865f39f2b88e760d9c8659ba3f9ca887b3136e3bdab82c046b145efd9c7ae1307ec93ade454479f2f324265564be3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17b98a0935b8be985b1cb68f88d770780e81a7850aae4f7f66864c069752a229488124074211f5465830e7553fb1f253900dc50644e58f393f630d4c37ed1ecc6969a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2a960f8ab6bc9a977660c45026cd2da30b7ccb5a07ae791cc79de2d84326b3a5fd6ccfed5ac9620ed31b8a3db44c6cc70733ecf39538981282faabd8f28293247120;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13806e9c6875a6fc0929065f5b88373e7c9a5ce7ebe37b49598a7fc3e3b9fb6e9574670528ef23feba4ca4500b8d97e8ef91173545cd948f271f27c53180d6bd32710;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd850a5935457053bfb29400ebb14a7ddc563b87c436eff129016a682461d3e3c5ddd73535f88845b87474e2183cc4d2f28b86c641837527b99d61646ca427ba4bc3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b32878a0bd6ccd33a70b5229aadcefe8f2ae19575652277c0d66ec4aa1976d8a657592e6424a9cb0326fa4d7f7ab3a628daf68506922b30dbf30062fed7751889e60;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b919443f03ce2ed352a9276192307b5b86a1a260342d4c1412198b8348b2e6512235fccf3e02e3f92ba71958b00ad321f70bf822bafc2ff36d169c1010d82b42191;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f64c3fd3bbceee44853f6c163eb4716098d96fb9b68614ca49809bb76977662284888c278b0ac601b71d81df9a16d07fde32cb9e74418b7c5d921f83f5badfd0be7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4212d9d6be074028e25554e3dc8eb6fbe5fb6355c41a6b9a83f97366f21b7013be93868e5ac90749d09ebf930b8833f4afddeac994e5080f22874e04b508f10e0dfb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f21e39f12ae515fb094fd9b024fdb2554f04b8a3cbc54d7d0cccc2be4e7f1b1735adb4570daa1da3befc279d1917810a09e3a79bb613944e1ac2be61a9bf0d82824;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf63f20a599705f6aab817758bfd9ab66b2fb745ac9ab8743c7d24a34a25062047c776d8f5ee160eea8013fb84a08c246e1fb9bb5e7b64cf162dbceda0f04e4bcdc88;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14e775997e3db780d76e80f051ec8af03262d9f74bacceb6fb3340d7af013df7586c4fcf68c3843a824ab702e3be7d7afdb2a5b0eb142a6e80f193789c6676c6123d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c79a49cc308bad29cdde8baa13b3568a6696ad2b7ecd51bdaa11f995187f9c55ff31a88876d0884409428a2b09ae9b7ded85d59b42e2869f0920bf4ba5c56009a335;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ee56fa54433ea58246a5648103d9f0d502952a39cf31cb8e0ae9bcd18e8eb223614c992e7b4f5979794dc8a3cbcdbfcabc4b347b747caac1c64f3cd865cd2ba789d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101cb2b35a024d62636623058bfd2902c8f47de9bacd603d2313a5dfc6989f1b85976f002d8061864ae6437dc96129d4e814fc656c970426702e1fd174f9ec7753ea0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h176d9ad4e4160a5a83f77e4028173ba81fb0738074be5a7d0efc19291c2f34212b162c11cceb274a705268deb2344462eabde785fdbcc68d8becb5d41497bc3681ce3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1813c9f0ec09e2967379cd5adcfd1788db0ece00dfb5b7c874db17b2eb66560128785421251e47c3da2cf911f170defd06bfd529c8d5df1219f67c6ffe9fa7b613c2c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14258167088857f31c6d8fdfe9608073378e731bd2551c84cbf63793df42605783c71a5173367c5abfa739b39fa6607bbab029179db0086474c9bb106ce1ba300cd7c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h382077f196363162b2b1351f0be497e25a891db85f88e976ed308972673c9b60312e90ed8a2254f5fdba970f9aadd7ea829d4f5c7d8689bd3175b1b9a95d0841657f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10916c59b9633ebba5d0b61f8b69a0245cdbfef67ad238b3f43b6bea9fa081bf61818c308263e671c0a04fb237bcfeb12d1381e122f4471f5081e28294fa3c9955a76;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d429a7a98d1f33a00c597d085549574826fe69d96cd3430984af9ce3f6e277f136eb9c32363e88e9a0708a5ae7f854078d93e58bf744230652141f5ed09efef55ec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe7dbee7d0cb91ad78474562a260ce19bf6d6a73699684d6ed253e6cd85c71917e05d9c03e3000dc2cb23c4810f134b0c8cd071af12cc59cd794a0dcf388fac83c5a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd32bb8fa880858abb25799532e8712d8cba4cbd5b5f394f800fb0846ff5c127acab8ff85ea5c6e3d687419b778002ea7af12a613ed5c1c8d8138d2d40c729592d2bc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ca2360ebb028e9cb909a400dcbf5600c7b414f4eb0a5de772336b9b2b06de6c1d81048810c1b4094974d1386a0ba9dc801bc85f2d3ca271679b3834b32309c52a24;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e10de2ec08f43931958144a86dadb8608a737312737a45046d9ceb665f7621b64f48fc2751cccc1fb1a7cff095f3dac6c37821a96e6f003211ab43a303fae08884;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3606efdc13358514f32468cba983cdf8dc5919574a716de6906d2e6444522a9967d7ec5ee9c43378359a23b4954a51fa0456c59ebdea48c72b665c8f996ea094e01e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13710b66270ff798d94d084c8a0751eb20a5db013c72c6327ba8c40889981afafc2e6826c6ade836ff81fecf1605e2a6cdcb50d67576e1fe3c37f7c05b814327d3aba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15393c002a38750c996be5e4282ccf171bae6d801b94202d26c4d898a900623705c193fc72cb0092db8e08c847247324b86c2eaee9860e3415674d9f34a049b81d567;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea7897a7b543498adcb8720963c01528366f7f7be2b4f62db5bdef81f99cf0f095c83a437c5e5c6f7e30273d2d2b652654f14b3cae335395f3961610d205777a7f6a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193494a443f8a756190252f16d8a88cbb6d6da468235810a90b7f17e648d5dc9c9c50d1bb3cd2cc0bd22d58745e8b14237def8861558f152577902e71a37fe8ab7216;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10d548d84e5959d8770790c22c105c6ac814a6fa34f746a7663139bea97779b6986892a7d3efad87c6d1679f1bb62f3681470697175ec7900c658b9a673b5ed15c224;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1851e835daf030e02e902bdfafc306f7edc7eb5afe0c4793ea903685c03030204b240926d0016c6ec3a1429c0c6a67d46f459bb8c173c812a026f5fb1c7c1dc2d19dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10fc6e08e3094e57e3986964bbed301a3842397ac118738c5d5e59971591bfe2870ae5b06075640fce5fa2dd717ef14ef76fff449eed23d04f5cab139c3e7b454b9f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h170ac2da25ec449c6726ada3c7e91ac13ae6864e3752ab32157ca729dcae915ff48c23182e764086d6475aede0262913db22b1e38272ed5a6d7cbb8622e16e3052c9f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb33dd9c5fda625b45a54689856490275f8cf4eb2b4cdb25251d66da075a868846b967dc9c69599fc67359454c082f189a0c2d089f5768a27e8a24338fc7b662d5fec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb0108fc7e7b06aed53a7e622109ecff280f9e92a497fedbfb741cd58544346511f99e498fefd56cd1dd4425a1efcb53d3c8247102a2f7b9898aab515961cdea1053;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1673cb06eb9b0c021d550b2ece2330a734550baec93d3ea6380f42b5e73c1aea37b17003228e695f9204d173fd6429247f9552e26090f687d33dea302312a9850e0d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10cc39f9dcee5363368fa63a634697bb7d8dd8530f8abc386d17d0dc47388d85ebec3d6bb1ad27585827c3a544a6f0791b339d153ab1d95bce710c66cb666a75c5c02;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he6048e3337eb3d51c5cb487354bd74969466c3a3222ce7d9bb1792780f2c88de078aa62535df8f06e6bc6349e4f9113a7404cf7bc5531b24ba5fec2806b5f6bad445;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eaf194a6e9496c42cd312273ccfb6cf9a73f2816fadb2f6f24cc96f202ad60f01c3f453924e43a674f2570fd0d98112d10be65635b8bbaa456641a891ba38913d1ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h993a67f98b10f09fd0033af456489a6ddd225379f87d86cd9494cc8247a9f621482a2daf65c83e1f0d2cc089c2b4eba01623ee77858a1a772651c5b12472626300b9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12d2f382c79dea666b4b8bd63c2bf49f1f35a1ffa602c893f581e358dfb02b2f08924ffcfd2fec87a0979b9fdba9289eeb8662bed3b1b1fd0fd895d90f01dd1d50d67;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b38c88814cecb4737c51d755aa45f9499bfedac68bf358308c26160e9fd79e3289707e65c4335b1834bb76d425b7a24383b4d628bffb9d8c27beb99e540e3112eb34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0ec0f661cf43425de42ee280d094c449ec6c07c8c7bb97e7159fd3f3d2b48d8b24bdc64ac465d85f9351ce98af3918125a91b28f687d4bd44573d1ff3c5cfabf629;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a445526599d0ec7e1f7970bec8ebbcd9c16ca52973ad4a086e7766d6a119f971d1adc3c7ff1dff9ff3d33fcfae35af69bd58800d78c727f67d771a5332c4ef7da61;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79873ab437779457a2a4526d2e1543ff41edfe79743454f12235212dfb65c9409fa8817479666d50168ff0f8ddce48a06ee668eeb98f5c20e361bb9b9536b625e318;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h630b92fbde2403f2b5a5b2317bc1a1694f1b44d0551cfcac7988471e65708b3b8288103508d1beda49ac1f1cae429528f96399aa9a44cfda8ab0ce15349ee293e968;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac7fae6e80bf85be147803e4f67f885d3d7b125ad0153a8a5765211d92759314e45a5f078e7f8cdbc1c427456fc5be428a23b3584603d6da7915ee57f1a62e00aa0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc408991731cdae306ee0319f070fc3e9ce96f45b6714129a199929c8b88b69f1584ba59cf940952ae30a2604056d2155efbfb9e6c74f3c43f0a35f2237c446f0759f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd0d43adc114ac5f19a7529e65a3139066ec8ff552fc81a06df5a8f0eb527a3c8bc38082d20cd8c4a8de16b30b58446ba71aa9cffa48df2c54c3fe00f6ae4b20a8c3f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1833d92ebd3a35093484d946e89990ad26943273a596f76f0555a6770189ea3dbc7a710b9eb4881448711c3a8ab16486bedc1b8857fcf64a310268bd660a1a859d549;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h311b2a263d69d8e60a226eff6dfbdde3cd33268826804c044305fa569e076fbd14e60a42b9acd875898d0da30fb85f8c7f8b1ef562fc7ff50d08797605b8b0729adc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h436719ff9ca8172ff48bfc2b7bb3594814f1a2aef46bbe0aec969b26b4e638bc20a6f83efc24724f2b966da05eebd758205df20ca6423c2270ab31ccc7ebc261c0eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd0080892b5d12b09c80dcad68bdec52139e82a17e3aaf6c59c41defa1788a8209428906f9ade0dc7c56067ce7dcd62e1092a7160614eaf25fad9d81a86df00813474;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb63e26c7a345be9dccf7cf376f90d90d99c3dd8cc555f559f8ed012dedaf22ef9ada93fd8ffafa8b4841ba75c7b3586bcd7067dc08dc664733d81e41df0cc55e5972;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198b35032d35d18c773274072f26f04ea05f9c1b47fbf18e6f2abf06cfd57cb0a029a72ca22dc183449800076424698fef3818aeca9fd523b5713d268c6a1766651e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7418ad5e2e0636d2ac4b3bf54e1497f8c1c96ce50b770bb945a25914f6b104062f1c9a39ec651f414628590ad465b92b47fa722a36cf0262b333a45c8f860104704;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h144315219cc0200c9db31ee2a3d015b3455bd4307f32b6bcdc5c0b6699879b8e93f918753f144bb05ce63996c07efcb83d7e1cfb0f28f066814e73a6fc8e7137f783e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f6b57c72c7d9515dd8e70ce6cc5c1143143ae6424d96a05118da3422e87a9fbc4ec5b2d0afbef00fee87a85ecd4b86570f8ac57a35e6887fb078fab0dbc1e063518;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1032ab3c5ef24b2d0fd9366049effc6fbd8feffe887fea57d1029c54ca4e71619da00ba2e1421effe338e7c3eb1323b2bc86f3da909a84592ae9bc44b0eaa9f6ea19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdaf9230304918caaba3e40784b34a4d68d623cdae33a5ca56641ff31b5d2bb3ec419989d2c6d9cad785b83d60244f738b0380b7096446f1f655bbe76a701301233ec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5aa63598ced2dc78fd709fe3c066fdf4a6281060eb45c49168e0b3fcc034222a18d8ea0df0610db68add8ea06bff25eba680fde0d618090b364b437987ac677efb33;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19273d35ae47a34ca8f6336b5f14cad021d0af9649f9e318d5913ae8dc5548230e2a3ea4c58b3c7caca1648631df6e173170d80f5c92d81ff7d3a8b201ff0b29a86a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3b8daaebd48f43fd5eae13515baf5a45144f622a880e2e79682e106c4c0b50b1647e971f7faefbcde5271c27e408ca51e3932d76b62cd60232586007871a5e4edf7a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4826f892e5d87104d07f2177ef75f16c95bbac67578331b5f080b7e720b937a6b0787e16edbcf0dacc7f4c92fe94a812025692d2bca052b4737c153f80fc28b59e71;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194a75e219c6c432d5929c005302b31d538f8264bd975c1c3f29758d22f216a5cd82b16c3cbab514f8e4581ec894ab7ffe7e86759da1247e2247c8642b296dc22eb44;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96f7d0528e10a70b04b386f4661095566c1f3af719485d555d1813b62718f0e7b29afda786facf98ab3e5d3aa32d79f2a465c47230745eb89997f86f30315a2bcf1c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9beac1b54644d30ce30ae1e8d63ec90010739ee10f1129372a86080e36774ea863cacc1b763814f21257046b092ccc654b3aa236e7139181828fc9768ca69c271442;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbed20a38df478f899ee9c9066164324035930c2016418d59753edccf60aab64f5ba375a02a1d513a152f96da37e8acc90cde79b5cba697a74415c1c4508e52008175;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a119b8666bc3cc84f530064973fcb32b364dc0b760e533369a5730bcb78125aa34a2ebd4eaa026a193a93d1e2964afda05263ef162e9c35fadac940cc9fc1583a184;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc7b1427b4643acbbc0019571d4fafdda491468699c0fa46e194cfaf1156a2c9b91eda750a0eead09a6635b9c51149d60a6301a507507861b4586eb2569cb2715bb2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d78b0cb62088f48434fc6aa6a0c0a154ddb66b45b33cef1248794ea6585689bd5576896318afee6773d450fb72dc26feab1ded3f3a0c26294978f222d4e22d2d2f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60cad57f3930e850fae8b3dfc7a75d3b50bb2080f484de99a77732ee3221e25dacd007e020c424793113b2ed759ff6927a92ae6546807200e04cac06dd2e6ba78c89;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6dda8ac9a3f38b1632f0543d201cb542263cd4d8f51b413de61c14facc1acf54659d63785719a985b57a6f189c6d3993d67eb556d80150939332dbaeb820f306eeef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12110a15f0e0d6ecf3bbeca0aa554636749343501d4e2b7a114baf870a60208ef5dbeee3dd8475c6572d149ccfdb2da21cbf79165dfef2f24ff405a53ae2154834d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13cd2546ef7ece64e8311580bd34bf8bce915bf61e8071d94f13c563475d39ec75f30081a441e52590cdde62f0090c7503955827c4fefcc781fd3e9b50e5dae13c08e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14c572714d74416f1f5d997b2a674c5ae6d9399ec7c2c2d85c5575efd575ff26fdda404b22aa5e1d2ffbdc89b5a1115ab489d3f6ff29b3be6015b519fd5437e1fcdc6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h682414eaf2b519d5e8a827249b75466b0efc52a0afcac287bbc2b6dc24e119fbfa792fdf06f4b25c8b6f3ed6db348b5d94a097be36eb1ead280ddf595cf74f836741;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ef91177f35374ebad44f83a82902feb058d803facf17592d4a6fb191d6f04990f519229a431277598357066700c5a5d4962c43c6779710641679d123f4b220c6089;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13cd59782e3fcc5dfee52d497c2c7d28b4b334923e75797bd604bdd6998548f4fc05f7b73f708100d7629ca91f4dc289cf314b0ac3d551b9a9bbbfe11ac30a8e5e963;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h151bd7e337aef46a4903a82cea89e216fc8f9fdfaa0257e39770ada3d665bbc29c93e240fbb8e02dbba36c407f6cdfbbf3936e6445c6d52f3adcfe460e2aed8213def;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60fdc882948c30564f0fb9017f1f51e677c4119612ba6d25e0a186bdb02571de5c9afdb7ad32b8d8602d09604a30aebb928ce06ea27639a7d1aadf819c33cea2512;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h192a61dbccecc68f50cb32a908388f027508dba2e3a88b6862da181439c46fd3f4585f440cf4d2f5ed233d5aa2e42e61731c06d74cefa3e72c2e29fc57610eda404df;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h115aaf72afd4cf0cc68e3132fea06c95c478c7e73e6a55676397ef949f44ab881cecb701dbad69000fab8760e353102295469a8d9c009b9c9b611c6a27d49e4bcca24;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a01bbff33406ae0437ce3be51ba26598915ebe4b212f5db3224a43c6609aebeeef1d485e1dfe8f23ab83b8991f6aed7fda1512985d14f22938928859032e8ad159d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91a16ff679cc724d10abc9a878660400d355623a48b76e0da141c0a6e4ae19d6715976c7a3906039483027f3098ea3e3052ead8ae965f5affaa5d5f7fdf7e5cc06f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18307e295203f0d74163d22777cd9de1ef90c38b9c5742768c413c9e122707be64637b097825b7bc1742121b395ba07b3d3f0e7170d8071cf61f219e49d34f72d8391;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc8f7f56f88c6e3667886dd520029570e73f6df5c0ba16add41b54ba39122318b531d21272c569f4d41afa5f4d7f67629fa546076c56539c909d597cf7f6494de66eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc598eb57f4d73a7763f993b57e0dedcf9d505d698bf94790db188ae4866bfa07e46968c61ab0cb17bb024d50e59bfcab2d02d587bff158ed3ec1d17bc2534d1a63ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h76dfdbba2e4bcdd7012a483b7f6091a963aa5b9c7f17680b1825bd63813ff5a30a6f542881279b78fbe584e5aa2499e6fe6a79850c1f60d7ddf66c35d5f7c57f6884;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha326f606d4c25c579adabc6b17306cb3c9feca815245517b233aa07980a7188a9c92eca6520b65e4d84417c301864eb7d23a42f6a7fd0fe9914ce63331d89b5cc633;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eea46b6b0ed25cc62447d0889d7a841fddcef4dfc0adf5b7acb1e08b3d3d3fc20c417e5cf3915d902456966a548e51717940977fe482b6e0cec455318737792ed6f2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1870a958bd8fb3b85c5beb22bae3401b6457395ab54592a32d9a1dac3eca9c8ad41c6e4d2d3e31dbfc02b7ebb8fe5c6ecb30474332dc373a6d4ad8f8fca647750bf22;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac9715819651391dada2b22c5ce8f60fa53449ffb1177d4082f793d3c11e10a65c11b45c0ee60bdd099646f8a4f59eb74609558fe840a736444612eaf98a883b3830;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h109eb3eaab0778f4b93ed90422ee080d3c8a24f1f5a5fff384f81b1c6d179e5d847ba9dcd8d39b683dc5023d110994c34ce46ac970ca3eec7bfb50f10b32e8e15b335;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef512ec24e87eb3f805929ee99340c83d346cf14ccb5a47df431698558804681e5b5cbf08b2cdbf7c61f2731df66a9fced40cd0c001762918935049b6e8b9f428d2c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h773788a3cb76f8e1c9a27144e53ccdcaaa830a700b60c3698818c17515ca04467ad87fe35056cb0aa04487a1026702a7b2509c92964a324a76d398143058e3f299ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b4ffe6e48c919e7b7ce415c8491d48d3f2c5021d575f506e01db5e8ac6ec3532cc6157274ba5a730e7e9ad5d8b91ffc0007638ca5aee96a82ef4ac2ef8b295a4d8d8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eeabcb46e2d9f6f81efd65fea627ac5c5d38a6c129c5001d151352012673c2f7ef6d33c4dd780e61b9cbf74fd1400afc8d6c76dd07ee611edfb648a066f5d15c17a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e24930b76532fc0239e292a3521938d6fc501495692585e69c91a039f66b62feffca7f7235b8b8512e7c1d9388c7d5426aa08260d3cdf10d77d7f3255b3e3308cab0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd530fc5a1fc5a3a0c99f242a2264532dc62a464e979b5476ddb26eaae999bbb7b5b89d50bf199c11842f56b3349747ef53ac764d8469e37f6800717b21450784f702;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7fa304cef56a5bd7719edf3d24d8d659bdd5ed25729a84d44d9bae35f2feb5c634927031a53a290773caf511df2be943ec3a8490469a6dfd7d6b48832efa603302df;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h62e6d8bf6174703a49a00d55011c59a9f672b25955d1d8f67beae0fabe7c69be51bb856569899e635155a960a3b123341a93f4011bf051f1e9ae65c1b0bf87dab4d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ee1e30cc1441879c2e9c2b85d9943ece32450a2ebcbbbadfc6a16178fee0e0c4e0ec47003096df36dc7c02d84ddbc58b296458f538ae934a29b1f0d585c83f1c0c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1838ae02a58e7201ff67c02a290431e3c886edb438baaedde3c627ace61e478470cd4d85bc80b73019e9368bcadda5554b466f0115684b7deb64a22af99b066e482e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7283d67140f6fd823df1adf221c07264f214d8385e21a764dbb774f35da0839077d358909cbd3c1c60a1856c0a132de99d6475e514a54644b5f1d613e754ffd4e1c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2ba2e3ae36ce47d69b2b950822e93b6b90074194a3f7f0b16f98c27212d0b2afb5dd09fefbb0a0c214363a2962a3750ac579a3fe72e9aa9448c5a3a0500e1b4000f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b9bc5319dd5fcac337527fbeaec186545abc01ce3d18e05b2d97c23ed88c6066a3304aca0a62cf7276e24a8a75355bd0d99e1288b5eb685cfae8d5dc86940cd58d29;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1927034a8b957fd15975d83f43f2a75aed9736b28ab292681a6f09cfedb2e9385a846401bbdd4c3e67f84c378bb07e105e7bb3186a6b669c32bb3aef9adb9e0a690fd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7de84028d10d77c9809d23dee0e45d759ed94d84cf7ee18404f0bf2006017bd8e8c698f8ea34f3e143183b815d51d615ffda214306560aa5e4b28d6f25c0d0c61157;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb8ef86bc4a5720afcc4d14063ca7d42257ae46fdebeeb4bfa454cdb01da8107ad914298c7731f09c804632daaf7ebc98fa6e955d3c1e269106c09cddce937eebaff4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198235ca32572609edbf0aed4d0d0c2a578fd0c45b30a87f65a61c2cfa8bc09ac560d81dbcebb1604c3001c14b2bc59177aff5fe11deab7bea95a1a354fc46be71e36;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12eeb13e85c9d0d93fbcfe1a6fcebc81391c9aae31d6b2795bbf9ae3506f49283575bd5bf6f4beea6ea696bd2ba2190e30362fbb8a627cffa99a29e3e2b1ce7717d65;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b4a3816c84938a60f6ab06e0344c7292b5291ff4077536453a44158d1272e5919f6e43105b3e8cd54c1b2162b876b01b6e759f117feebb4fc8edd0d6a498efa2a07;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129cf2a391028432004ce20a62cc8fba556ba4b23141003b5ac05c135d8070cb3287335e4ffca94c516f9ef0acfef6e6906ed17c2c0316835a5ecc9860b9f0c0e696d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b7eb475c88aefd4b22b1b31688e7e1d3442ddcb55486a38c9f0b1b785367e164e48d64ece8f91777d62e46b94e5a538d8ec32f3e9e7e82daba9a7085168f7467d91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbec4c86802c861011326578e38da769c27a9f9836a3cb99ee1552deed8a3f8069b8611815912ed214dc5281a1c8e6e8f7a416e45af8c419bef071010a0b79a4e25d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h174d90569e14bb57fa095b2bbd6f4a3a091585793da640a2caf7dd3185b9cd40fe6c2765d366624fc253de9f17fea0d5b620d475ca9a4b5940839bd58c86fadc48f88;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13bbec9933fdd178f97942e7f8e70dbdbcea6526fd0fd4d62fc57a32eeca88a6e0d78d0f8df05b16c949bf6496ef5743897e720f136df3f681011829dbe1e8dbed060;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he431d6ea18cc231b22ae97d40f6f2e4dd37c5c882a5fe1499896d15aa60bbce6fbf9f84a70d0385f4152a236ea1707ce77357776e93f57b68b42b693c3d01b846a4d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9277f22b77444f13fd121a96f23fa3e28175577c1bbddcac592ee2cb3bd60f28cf57bd51be2837072ff09344b6315984202693149fa79b6c91bbeddd65717b0bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19997c1165134a61dec024dd92872a55895eb97c30aecdcc1286c8258c63d2002cf47b4ec96891c802f2093a3fae31d6fef6bc84bcaa7d8cad9eff83357b4f6abaa15;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ea0a23173c3b7d0e6ea7cd6861c8a8c6d3bfb73497c93bcb8b26cf9e99c2c0bcaa1211afd515d2c0a51fc7b3eed5d8f40c721b53bfce77441d8aa1a4f57f6048c72;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe632c167f99ff55c8b3bcc09bb8fdee1b58d4651316e25a81fba74310bbb72ab09a3bd5fbf064688cffe016b695d1dff2364c6ad3a7bf8825573bda7c94d26da9fa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h21d1494596ef1d4e003b16a2c7a3e5d784462db872da400b85bc90062d9ed7052f026a4c793d2d978e6ced614f33a83d7fe0d8ab3eaebfa946a26771342921fe99ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165cd21060a01998abd6fac889e5fbd209d73bf271e4f99401983856542d85ea6a49d991e441d10573fdab4aee2f87cf82d8118ee7892a0c2e237fa010b4ee47bbe35;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h669e440c5b2002ece12c98309cdaa7cf7e017b9e91d68f1706379c9625eb07a5b6715b1f0456371b47a2381b3caa554241e04798d0446adc7e173227d2430cd3c6ad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11084a68bf145780a455510daeef71a471c87de34a27e078274f0c699d3a18010819376c15fa3765ce5e4a578c1395d08d63edb89025d8489c583a91c52e2a571accf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h59b14b7eedff220fae59d00b46d588d004a126265bd6ae8a4a0b8f23efa4272647298c99d16dfd0d79e73daacb2e30b7d521d5f6d69a25161c44bd572c882dbf4203;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h95f8a7b597d395e69a9d6f6085ee9ba2ec470f739a7096c154b710efbbae3a162559a52b55b49b2206f56f1cb620ced1b46fc00a084ca205defbfabcd217126dd21b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hda806500e5334dbf08528604a19cbd8eae5328ba61d78e97fa400a0d66ed585117227c21675a39f913f6e67bc90ad8dc5def1cf4e86c144e2ed66ea0962cde997a77;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h141b143f459b8101d14ec3d5ef92cb733b2fa4c00a307ce90bd7eaa242b579fb224c49220fa4df8114b9ba6dab5c9c33c1554f38ea970657dd037c809908147f66eca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d0f730ae13dde8ba72f80c78967fe7572d284eac50e703197d418c5354dcbc795c773eff9be9c025da82fa4ddf12099584dd7ecb4fbb3fe633d566dd2fb487f115e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a69c96e17a0e9c9b42fa038f2b8ac2a48feb14c9831a060b403f9c92624a5ddc4ac2d4509282deb4727f8fb3391d4aa8159ee9fc7dc19f2afa9eac64a33023f35b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b0e453fc2bb80a6d9cb6ea0131aa2f8b15bce4ace0656751124d9985ff2c0156ba5043594bf185cb7bda2a1ecec676f968a740fb44dd8e029b44efbb9544b13dd84;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf6181b7f760d8c1fea0629e8966cb583b36973b2703cc3d8bf31981d13d64b6afb08fbe6754f41af072c6b7b1719cdb48375528a6ce71581bb8b05e15888c4bf4796;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd93241bbbaf2b40df7195504a2254aead655d1bfed8cc1bb585555bdceecbf1ad52fd32d5cd9d5a4052f0b97e65231479bccf924cfed138d801971e54cdae040da2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha09b936d19d752e05fb25e6314dae127bb04175d41db16506b651f5472fca57716de3fbd54982b7b8652cb8b8ccb4f8f4d7681fd7ff316e5771eb8dd87c1820b0ba4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h532da2ce99b0a655a8bf794b6b1a9f76b0e9019ba388dd7d28e7905aea01399bed2badc0e9d05dde0b0b5e6283911ac4608209b495d6b552c4d974fd5a2994fc4f34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8b0131892e65fa8510ed939bc450516648131242b0fe8c8a6c3977a8aa01a07187852207e794627ecaf2794d209db2fa021acfb51b664dd25bae201504f8c5641de6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48e807e88fb17f6c0054bcb09bd366635e60cd477f52aa525bc81b29723f74a00b1a088fa71ecd5a25f5332a2ba61026b2cd5081ed9512b77d1b91c0219da605ce48;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h21ff8024917e2c4c69c732be59a717c36313656273ec2f3449e8ee630b4567ee3a4191a9e84de75efe3083deab9e6be537cea80159681b26c382c344477fd3da875d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da50b096073cfdb6c692eb158f3a66c3ff137822087a9bda34c24e01414bc057ad8e3ff87d47a86c1b29c8ac6295038f48ee67d2dbc032dd29a2d7117ae3a4ab51f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a6e1225236c18f850911258391490c02230fd731c926659823526b968a88a5ad335d942a2087e561ea8dda309b8a9f4699694ee8320c26b37a6a84dbf43cbe6f3f43;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1633d2f87ca7653322ad3fa434f580c79c33682deeccfbf5569467398bb008eed9428a1b95d557f1ff8c283fcf98f4ab16d07318727b7a061879ab7882e09ef04d7bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cb328f1fe482d601e14f23f1ac6ba7d92794e17f3d2179f8cdccb421a6c62b05629c6dc42c6c2194addbafc637acf1c327482bf5febe8d3fc7fb20d6d9baddc9aff7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfb5cd93aa08969ea0c48be791b44cbbdc506816e5448cb79d0d5c44c0f42a6c7cf114cea96bcf5dbe1e0c48b9302554054d1da13896d7d9f0645b46e6948a8a041b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h114fd8b317f098a2b94c56c66097515861f9d4d64cc50a3144d3f402a685e674663013a850a0e2f61165c57c17806b8a3b95041ef8912b933413357772ed34bb9aa8b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2f5ccd298e2b153bf8a67a930fff2cfa4ff02af0c1bc103b50b732d5e243736d68898d45dea6743dfbac976add31c1f833562de09fa58ac6a6d09d811d71ebbcc2b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e8e8ebc4a1e66982e3fd7ddbbd6acad9cef9d630d2d185e2c758e80d8b616a96a6b5b23ac254a8b5e390159c33415f08c52868c4e4f2b8fbb238878dc8177299fea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1426c255b6bd7f3a85f0361898c9f56c57c2b3b28c9c4892e017ca6700ccb561006e90f21b87c08e20253921c98ed02e4d6ee045b33e2419c76a24ac283605fb69f7b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc62a927aa149e02aa106fd61b2a7ef3dc36fa0e2d2e92e49f6cdfc21f5ce013447bd17c51ced33670b7fe47e57507617854236d6ad227c8874151e254da26ead172;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b2d22ca27a6e643851dbff983cdf0d0748aa160ac7b24fcea8e4cc09abe3ac8cb0c77e0ba4b3573d8ec72e42fce23a2c23861686cfda0d9f0aab23993bfc61d51ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8865c2ed541ec90f75544b92323310e4a73921c875b890f8e0b9f619e7e53b49449f89f16ebd8bc177ce0f92effefb84f24bddf90a04868670e06dbef7e749428048;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h76a148f9687066adf8376a13ad6da82895bdf58661333001b05999c1aaf5d7341c4cd7dd9e352488531e1a003d853f91ec0d5c09c3fd0f9ae568b915736668314790;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17d2bf9415a25a22b6d632cdbca244a6d46457fb4e3f6e7ea4df92595c425b152d393c5658879bdb472b12a6b60e019830d06dbe1d3c3359718ff86466a2195cebeb6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1567f1b8841195d8732528e665a2a356e0735dc8d475eaf243f12ecb04ff05ea62acd20923644cd250550eb695ee5719acf1a28f182ef0d73b1e46ab7a07ee1ee2a35;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c66c042ce2c9d63cc07f057f7c99d7a05c7b97d6f993ea2b103a25fd0b618cad66fc52b09fc7018ade0ef6384b43948aa99bcd2471955953111b7caae4015f4f1aef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c26120bde3e2b9c40c446bc7aad76c46e3c4b2a8cdd68d61c7afd28ac23c6f1ecb9e282b4fadfdc7a46287722a65f06978ca69f90c7012bcde65255f8632b0fa54f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c5c2551237a66c09fbf5580ca52cf6cb7df53d8f58bed0f46e8831320ad991724c6840c097226bb9edc8cb0dfde8c0296ca4ac3477a56009dc82d594ec9b577fc04;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19bd2ace6b7ce1b3fa9e5ffe569017f1c33457d8c735a4a2543c3dd5b56054c84614ce015fdd0dc7ca78d870a801e96bade39f5e470fce8cee37e4b3d3c649ac6cb52;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f710010958191b06eb35501691159eaf9d59e713c82167173cb2557b55ca9f19f54865b483079c93cb25c2df5f81c5f6cb60f12cfcebd5717502fa5abf331d1b3dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4633346d1bb3d98bfb0a9b5dfac3abe63bb587b86d64ee4b2c9b1d75dd80d60b1940055e51aca93cb97f02771fbf1719259876534c2e5429c6fcdb89ac7e7068691;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1db65a6b9a92c79724564e0d3032052984e03830181557cef12d213ef08729526cf965f8cbc204dc0085bed34381bf63dc423f4e84241c950f2ea234925adec1fad35;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71ba9293c5302b6fe63885a4a1994c808c4fd114e556c1442392c321e9ba0cbc63c9c35e54cc2c08c0f6e397cc0db4283a4d43293854e74dec7d548f987fbaf87cc6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171ba16acb6b324d4108c7a64610315408293371d40fb1b20c85c52599928f7fb772a27c1d8822403c74c710483a95dd428b0aaacadfdeb508643bc3b00f40fe08868;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b544d575d18fce28c4c7c1783d9cce548db759f259fd64eadb3a6eb59b84cc221b66a88ceac70807c9bc1fb77b77df5167bb0bcdbceefc9dd056678d01e75823dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c2bcab9742acf56d2691c9deef89e628ebfb7dc31eb765d8ea4c2265e1ff09d64251aec8b892e253ac0c3334546e35244fbe77702d0b9ec6770cb599bbcf94073d9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11aa2e1e973987b9d00f2e16b230b0df2ce24c5d24c22aa0506c4f2abaf21fb50ccd6827809173e7b906cb4b3855abdabb70180c17c35cb7e7669ade034e3ea4878f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8760d4e3313e4a90693f4b2ef291b7d93e0c58549c6e35dc12e1d3856b20eb9db7f260d8dfccfdae24a05684b18f2d832df7cdc7d4811c7b3fa77f4bf292c4f98690;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d3f4c08c4158a53816bac948f477bf83f40535738004cbd20feee790315d1fd2f0925716587ff049ef2fb97714a88bccaadb26bfba880615b96e7985e705764e82bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1441e4c06cfd763a9b4e45b3ddbba5429689e34dddf43e7f3f0d73a90cc0a9c9a43dfccd8a2ef311a230fe7179c44613d342bec38599b7b06d2bee06f9ef695810869;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h986f36f7d7e941df1cf90138bf37a938b925e632c80320f0d50f4f17282b15f6ec39f818b04d11916630ff606026a74e074998b71ddb7bb25c39ab1102ab755b3229;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f4688632b58fb129767a0999f115b9076ce0deb91de9fde399ab6c21afa1a20eb7fec9e85b83908c61637bae3e7b1108e99be0a613190dd6e0157c3c71ef1ace584e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a5e05038bae9a65ab7825e6ef3bbc9a2947d322fb76c91fe2965a1e9b518fbc52c7a7da36ab69feef769d31dc57de657a0e4fae3635f51648de26b728f8e0ed85163;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h147f41f3eb3385c7ad7221dd1bb27a77abecc1a983d247231048c53ae89b9cd577561316ddd9b1a11a1b1b6e2e82f82436b9a7b5464987d3a7638d0cf8ec350108c5d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b1fc550ac3ee5f37990b5b4b503693fa0c7600d171fbb295175d5454b274d9a3167a8c38fd313b53b7e0914b254bd1a3063376aa84fbabe709eabcea4df14c89fe7b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14198ed28e88a07f6055dc54c1f06f70d062ccd643662855f2d7fa3b8358a9401520a8a231eeb04eb659874c96f28544c20a665f8f31aa54bfd3878ee975e1e154707;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he85843d8742f46865696d487a8bc6afa3555ce15e2f08e24e85b5d9b63ed03240e2393e55e2b9f3987453b7633ebdaa7da0497b6c5ef42a3b1abcaa1f5cd060a990a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b5c905b7bdafbe05143b4466dddcfdf18f77e78bc8d65afb5e54a1fe3b83695d9c18b1c6d912692c5a237add15fa86a3186f4264921b6156b6113ce7be27b3d2adc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h26ce396a19b4db86021cea71b8bd3404fb61c8a16f39745b74846443c0121e9e052cad9f9bc821a788b5f1686af5f5da56e50b9b5bb012b945c192c8ae0b8ce1c7a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a63574281f90f8e90ad04fb1fa0f0968e8d05c5f2a12741a4d0f64f2af39e0315289f71289a280e7b064885aaf29d4e88a4e5ddd649f8ecdee488850482affc221f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18492b1233711c1679359590ada5ab8e6843afc0aa8da22253e0fc04fb684ff055ba8e60fcd9cd1f1e236d7d0555ac8923c764f730e094560e32ef420144d893875cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5a241937ff3c220d89eab927bddd8444813f2900dfdfa1fd8d920985f200a5453f030666bbd5859e189a5e35c780105f05400b9d0ffb0a734b713a51a63711e48afd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5da1dff612be0680c63ce4c7aa171f4fd4ff4f01bef2a53a9c2e7866e4cd45a46e27f3ac5435767992ab6d4e800bfbae3cd8e69f3176327d6d1aec42e96ea8c72526;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2d5269ba5d716a205988ea475d0d4ec2686dd613b15a0bf754e48b6d598b82e8962a586bd52d56d834cf837b013b60a99b1ba9357b85178ae304ef413b491af6b448;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h36aa630d91ecf0430be1d66d3322b0fe6ebd79e13fbc5f70e28f7d7aa4b7078ba22f1d105bdb0339438c7da204f546a49b75e368a1e488b5224444f2e336f37b5e01;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d7fc824ae473c802b887a98d0c8ddac628b196865bb95ecef1c5995fa89c7c835c0e4c927801645eace31d5b73ab930fc4746d67f9946435152d9ff0c6da39776c6f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e911a5f1e1847e86ffffff01a1b66348be4ebf10b563dd5d4213cf33488587db0b2e4ef04b0fc82109610cae34729268fd372e68c290d5ccedf53ebf9da5583f79a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h26c55049ce6703a36411d51d02b4782e49760fc6a0a5c58579c00b9ed5273ea0a47fa07adc452d096d8fe759436592388b0c6b20a5c6b5e7b2e40487c83b1d8a803a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdef04a5648bf7bbb369dae09581b0923e981a275067e1626ec619aa3761e0ff1977246b2673f70c7bcc128948023213c83d1a2a889f1f2172659858232baabd44984;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h32186813476395203c9b64c0b128af22d35108da2b7d8abb6e556b85b577af422e4c5d861843356c22427cb3c4d049458f01a1b62e11ab5fe2f2a874559d5bd63d77;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb7512dbc739617bd0f60ddb8e67c3f90e0863e19e76e640e148efa2578666fbf2d5d446e3228e627f18866c3561a7b314a0e7c4d57e133e3382a3b770697e1d48a7d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ba1fb37b178f7bcd9444e9a22a0df3d46b471af0dcddcfd69983a74e752447132232ffae177709dc07743ca52e2600ea37fc993253cb832e154e1e782717533841a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d8055d9d08b6c59297050071d4b06417a2010978e16ab1e0ce9b4f7646a2b20291d1ea817ccbe222490769757c3a3dd42e7c6ebf16d94d50e69a820e3ff9d844724d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a359b4bdfd8aafb08ae6bc2f01777a9468660b4e643ed2b5e32b76f3ba8c0956e94ce400ca9013068f9e35e03c8df734bd67b261635f96ed62e3af1457010a3c289;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbd62a59a54b281c9f974bed1ee4ca3d43c609f45e6d21df5bf33b42c916a66df3d33ea8f2e449cf0bb679fca2cbf5da52eca650c05b327494e40fd82fb2d0dfe0fdf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f64a5e4969b2d373d40cd6a99ae6ceac816fb10b933d24d05a8551e5388571eb3f5f53701ebf9bb22fc986434ad1cc974e5be2d0380b3298ccaa91ccaf7ae6a6559b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a0b18ed829fcb0e72a1353055fd7071a53203a0d6c5cb7ff3bcc36a2be008b0325654a834527a4d51212f5b59a4811fc47b9e3ea37d9ea45c3ea6eef0a75e79b9a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ee4d6e0d11452bf4efc0e910b072a7058e7000a5e2a704d56248c9af48417f84e366ce47be758d104244f844b851ad5ef406d3e2d88089736ad85afed38d255021e1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a8e48763c9209489aa678435285dbbd4d1fba52824addf6d6826e0f8c62da149468ea75d686a0ddb081fc0582660126b9a4694817b0e507a1aedbc3e02d4e57bf87d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc2489a76d38b06f658c531fe50292c80eca3fa9dca21628e6a260e32f99f2c395f90a52ada413b300c1f70a8fb201e3d5e832ae941722e6a4663d6b022355b9fc7c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a352e5e528da027a6039837c556d0fb6c6703430576e01d20da6016c15e615314d31913a6c3069c39e74b383a693138d01c14b4019ed08614bb4496dea5164aae1e3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h336ff290d2f552ee3206ef22e706e82fa928992dc732272604702e397690bd20101620426649646717aa783a6b27ba571e99b2098d79328c0dc75655ae90e2fc1193;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f54d1113c0c07e80827b307f8dcdc9c09b17a696432a84d2155059c03ff5c7f816e1254e13cfcb492bce8be21cf61a380ef8b9df5669460e20dbdfbc91b172398193;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hec351d5bfea3da2eb7fdd1c1751945701f15e99ece4538dbd3a9e00d71c79c23ea43d198de434b8c63f2c9e84564b6a4ebe8768ba6eada7be5f7ab7531d3f2362d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1401697f09684aa1c22eec6de8fabdfef8ca0d3105596ae1909de271979943c6f7c488cc0bf80489e67724a12a5e7c979fdd0fbd2316d5e06d4a3bef1620094a81bf0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118c60d8fe4e9542a0071da45adb0980736472a81b8e7bec0a6f5bbc53af023bc3649091ccbc1f6d64e961c7f316529498e71844b7103573c4ca621872d8da8550b0f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf2dbcccec2ce71f596e3bd2a41a8529c5b183f2a6012dc370fdcb32afcbd2fb5931d0ebec48d77c98c9b7047e2202cc70c4fea8bf75fc664eb4c1dc036023a82477b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfb38cc0b6917cbe637340837e49a6dba0bcf63de1ec97e596b6a8682fdeec500f58c252ba14cc53264c0c6976a7ece7bd87650b58d996074f715dea3df8c2c872388;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d1b0065c6e7837cda64c9bb87d0babbdfba2003b13071528ec5b5b76425394a675834afd85b370d1cf60b7da651e9ad6a5d9f119e65697c832d0d6558d5117819bc2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hddfcdea5d33b84a2aac3493e0307988c52dffeb69593f8c58a56783b20f4f50ea7e22192940457f7fe6040e10863e4cdd12ba45efb977ff190ec4ce3065ac6a24530;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71907627ec4d977237705ad1535f6d4f566d944c517b894fe8f0e2371f3c1ec1d2c7d88d172084736dfba6e5fb3b14122f3cf8e3141a2c9cfca42e69046891aea2b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8bf294c60746ad2ecd3b4361b858379d8e494d65caf38d3ca5bd56cf30961798c2bcd0c12cf93e3fa32a6a3d318c788f41402a0750aa893a69ac30bd53cb52aad121;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d6c13d254aa1f6e738c7d0f4462babfea048548e30010268178de7e41f56be33cde8faf1fa9fbad9f27ac9a9d4522b1db0ad48025d7133a15f7b129312c0b42b75ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9733001412ea284fa4e3cea6cba4b52683951d184587965bc67cd6764ff1af7f8f6948b47a513963445613cf19cfa87277fb168c4d18303535c294789fc16ef6325e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h450e1af38c3af26f658ad37728d41b88d69c0ec86dfb12ca6af1986448ea2e1f037b992d035d3d070efb484200506a6c8c70ca74578c43395c93da9d4cbd5d4e61ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b981559474eb1b6b6c8abf1167f522d4c20430cc1ce57e87ec9536c67cf7c1379539c73dac19ade3f53eb70fda1ce4b237ead932ed8a98fa43d3241cae90820e590;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa11c80c603eec7a7a842ae2ccb658e1555d3909483f3734ef134a2ce127cf1706e04c4798ba8816d447617d78f3b30dfceffef879e1843748da488cabd20b83bd63;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11d44e53251b1fb344010f3b7008bdd684a587bcc7cc56d825f431a285e3a4084a76ef39d686b7d8749681a0abde0c719c6646e0825c33e064dd346c9599d7650a95a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1969c4667f41b4ce861fd22c2d066e43bf598e275977dd78e933146e02a2826aab90ba3a3e8deee0128815d6cbb9a2717e21ddab2ab21016d4d11ecedf6a4bcb06b76;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10d828e1405c8122f86e1cadf9c05eaa91f8a23b8da4dd56aa81a505a9dd5e1fa9297f8abc86c89c8eec57235a1ce7eced60c717acb275b88af81dfff9ce9d905f66c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h620b951cd978c378d52153870cde28c165834c976617b7636448d0cd1eb70784f920ebac0916dc5007450ef0f2262e4a0a73722a7015a0c5ce4303c20a6b5f317016;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f8d857588771713b8c17a8a52e4cbe7913b1afbb8e33039889cc71263ba4d1ea5ed11c46ca2736a8f10669aa65abe89e3ac35424a4cc5dc2fe852becb2da32e1542f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h137c124a8ab2b392fbf389cae4e9192b463b8d7618c567ab4a16e81a67dec6f0ca7a4b29a3ea2c4a69a6c1c8ca8deac6e20a61abe41bdc999753452b13032d8a4f688;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac657d425b76e02fabcf694d6095072bd2f6f4e0dd806be832e19b0c3574501e553d87a253f8612407eb316c5133768c415e77a4117a49d67833f40f107a1d63a09f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15bb2b648262cdfcbc331af6656446c47538fc628a1055b226f7c3f1efc6d9c280781f0818c151309ffdd2a16c8b8fdea0d1049c7b6ec257bd433077587549330704e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h32feecef72974017e74a85d2c98d9ba94cd675d6be944ff98ae3ca587b77cf13e6c440d9bd0b580636c7988d53cf373ae01f7eeccdcf4e4ce29ca681e3b31299fc33;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h370400a6efe2a4350f80665ca25583122ae66bd6506048740d220c22d889b83bc070cf628edebf7af22774bc609dc07dc43faa4300ee0ffcc1691e26fb532ea71cc2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165e2446b93af00b7c433838eae8f0ff35e3bfb1526e2c0e428d55f0ff5776f3b3c9bb7fc64fe72d190bc3a553dce7fccfa833438b28d0b5cd3b6e59ef41ff9d504f0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9f5bfcd0e4583007f9f708273f00cb550ddd3e27f16b07c7b97b67aaebabc81853f228223c32a37c36abc5bf9e08a3e59a369c818aa03135e0e58061830a3644a8e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12ace9d90c01fd6a1f128689fbf820bf60a87fec5dcf359dc6df103a0e43d5300745dcc04cf11ff4c58193cc194287429803ec5e6e50108693d912d5bb5088db42cbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h115c9193cfa5a2d4bdad66717d3ce797535fd7705a6c0e79afa839730ca2be80060cecbadf544ebc323f34798dbd2e6a6d55ef82ad03267abd449430920be225d1446;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f7bbd3c2abc2785cdc8ba4328d751943017891ca40ab717e11d78aa590ec1bce277aa7f3c979c41dbba7fdc296d618d71a848925bdbdd053dd063af23ec4620adbd9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0b983fda792eb4720f37774cab3b6aad14aff604547542fde5dcd9794f7e97c8ca2da1eb1619705ec7392f55aede5e29928a5d3a3a2255f8c68e8ef3c7448fb1fd1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ab6e2bcc8e1fdf90bd3c660e49bc3d1f4608c74ee6eb048f15bcb5fd2bfa0ed7ae1b081bdfd5bfaf459ee5d0ebfccbb2d1f012e10825b76af20ebde3d960ccdd9a8d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a81b2b8bbf9b85b3a51a391ce01b8dc5c3440282316cac95187b58047a423d77c0b82766d74a39aa0d720c159a569f67ac003d19a06f84011b025417a37a3de140a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc137774ef9532b470004a50b69c731102fea9e2854345cfac9bb3471f89ed53587ef8911047711bc2bb405a71b266cbbce54a4a349b0dc575d49f95854dca052328;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1778a864143b91d363118759f7219f3c337feca83bf67074d35a41d85c3aee44738abd1a3d77000b06d907ac1695dc128988969a8610368e08a330367af5e8b88cd8b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc1f3bac507af1e35c21e81afa4ffbcff88c121b0c37dd4bf93f8e1ffc35c685e18347b75a9c76e474d7b5427fd0e9a80fb90ae5ed80a42f35d02a25d5f8ee2de1dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h207fdc0af609eca79c3619ea01742068a29326e1bd942fc06102fd1a799d12aec3e501f102236a41f14e853009f060b50ee65ac7c90c83f1d109374b7c27a8933b1a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb2e6acc765ec6849f41c144a851cfa0abfe9c0dccbb8c44b5fb6662a46f26b6c721f35810a798968811e277ff21892ad5412509c342ddf39d8054428d836a3f4649b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f8a7ae6bcced502b262a98db501555113a8e6c2749c2c6151d13088e009004f1b2cda405ad5e7a2f82c6e38824058dd0430d55df1af1985ee37df5fe2af8bded773;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h684ca931c8e0224400e9cdfa4216a2dc637e0ac5dbb65f121242b65f16bf6953bc4a8c5f2b99581564a07310c019bcaa6c20c3d47fb5dd1aa0cc2d72c2201bb3c1c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15aa4991ec7fdb60204a34ceff7587aad1c3efe76b4ea33b096d264dc7ef256106004eea8ed4e21273dde46f4fe3d15553cadc533b29830b7a210aad28f987c58bd3b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9dfb1f7977bed2fde37dbad9f5fd0373ad4241356776211eda0c1dab72bc61bb94bd71811f17231be27633913637bd0b8fbadd71d221425b47a3c836968638be138b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e26cf084dd7f272154d61cc8c97b010f8b9656f07d77e16d8fd4fb271a289fc4aaa22d5e856d9f49d9534f114dd7c6b9e541ce03b82889a62e4a9583df5b3b62d6c6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'habbe86f9187b15ae0289278f66316b7d994da1a52d8319713aedac1e6037a7db441dcf94b4c9aeed626ea696f64473cea4b241c19ceec46239956a0f198fc86b9b3f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h153c7aab0b88b0257c59c4770513cd364c94a705feb236a8da29c121051807771466e656ec72e18b7cda1f5942add0330b7d8a7511166fdcf3910ff876a0e1a40432c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149ec33b374cdea82dadb633a5b1c47b5f8442663d4631bf007c6eddf03e2b7449d34925f85974ea8329bcb913849cd22cd423e8e166ff873a32003391793ecff7ed2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15ec8763d3090e90d3df0cfea03837820eea10e69048cf416a5f007b1cc802392e1ac8f4354bf0cd15ee94e1150e90c7af208dee69ed03cd259fe3e3cad7b3fe6c6e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h177d88170114a80c8f6c746fe185ea565d661ba58b27f0ac55c26b5a853e58970d60eb13dca8bafb989726c2c8b33628d7d4d532f899748e061e118beb7e2a5f32496;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3b01f5e29b81a54116f9ae8915916f23343cb967b06e9f0b0a58d8b2e6ceef82be01b3e21306d775c55ab6c641d26a8aa779c4a11d9044bad682c6fc3636bd996155;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1940ea01057d682f7bc3146e17f5b5ade29a726dac5392c11ca33de1b29e26b485004e5aa280cbd23fc049b5df60e151e57949fdd47c281186bc274f8b2a024e48ca2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc7fc075fcb1832991ec3a7b2cbd6dd82fe5e5c28d98808bcbd57d2c40782f4d2a2bc8ad2990b2d7b98f7d55c43690e61f5df3272ac3740a88607ba8a3da317205ce9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb36eeafa05289366ec31eb5c187baca20f6745ae14faa52c4aa6ad94398b3216ec5f4fd0ea9552f6697b461c1955f65e123bec7730884721ba9a7da2b218b20e5572;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73aa692dbfe3c29acca1ac8ec6352249ffe44cfd24402989e444b9a31a009c0b291d40c8087e349fcc2aaacd45c561f8dd58142cf4129e502cfb3d7ed76236c2a399;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e86177b311f7381b3ded0cfa6d9de37a33aa383e69b60af08ad122692f5799bc533005577f2e2de06dc6ccedf36c628cb3750483aed0323f06cd6b53874028fbef15;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he0f42e76aca5a508ecc6056164c0616306b2ef22599c00a153b0aaaa471b95e1ebecfb0d703d02b31cf86ff7d5d5a311df6a0dcab442f1151589d6f9b377ab337f4d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he00d78e1f15f8bae934dd235ba8c86c1152f59ca89be67e2339d7e01085e850329bc5911df4f9266ec9efc338d0c01e736b7ba37373be781ac9a3f1b788d504cec1a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he61b1634a840bff7007f8e29b70b453bcee894d033248c2ae339a4eefa838d4aa5d42d6c539921e774758da4e98df1a3249cacd8803f5991c6e68b02fa801918f25a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab1607cd2e7db95c962f5f380fe7ef9b8f881e1164521f669f69150870e56699ec8dbf21ab8709160e60963af50c40d54e0c4b6fa73263750c9733a03a13e273e2cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1090368febccd1010f45bb889a52f78429f01ddbd000e31c608be8756bf0fe170fcb082b2fb02ec0d5bde5e54c80deb6677b8f56a0aa3e97fe5882ddaf4e6099d49a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b1b049c9d8c28a1da4b64ea35940913a0bcd2a3401c9d2fd35c99f86549e407c4e9da2d7a789ca8643ff5ee9d01efeb4f77e2725681765eef10afe93d3049acc211;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f72c3b78e712e1034e8dd91cba30864ef2c37699a7d64a4e4da88ade0cddf4ca9ed16ba1e5c8d5dba908fcd758be03f0822c2470dc6c5ff1ec67f368bc7e9151514;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8c3689b5d139f7d3043804859c33db15f600857381324607e7900aa8ee95203be8716dac3c6839b60b7677e5de961ccb82c283a8bbaf78830a8236216c13c81cfce2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11cf08316094a3eea2bd0ab8ae5a88f854e09dd69c929202323caa0d92845c6f6a7338a300c07f39fdcbf128397692a05569344ee553bb868ae8b05bc59fabd00bd96;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a0426ab33f1ae539996bba0c1e7d7ae21ca1e60faf2c279c72da229d2c7ec6c50284c0f85e97bfba759ebaf47186ed524132c50624118b5195bf05af8ceee6aa56a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h54cd5ef96516d64e9f95440254baf4b03d024b9b2ab6d424cb79af997b53d5b627f13f48a4c6d11f3c54dcbd0b693578a25b21356664c33ce0008ed016ad773aff9d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12cfc181c24fbd27c542c2747c18b05594f3c4346bb0473d14051006ca194215f0254957a2239c157840893773ef8efe4546b179868e01c3a67df13040738b6f0bba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f85c3074b51ac74517be3c870b21a050f465135f4a82025957215caaed071c384e6c297ccf3efbd03037b260ebbde8b4c8a2df42732954ba1a6e37ecc85b3cb49854;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c065309ab96d02543d8db1e0e4932edcdb1d055149bec9fea7588c7c1aea642e6b55dd5dfa72ae1a2760858a16ccec1bc0d17953a276956ddb0c8e8fcbe6a4a2f428;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af3b94088cecef588e7361ccf872710ddc86d7d101da894623ab9a0085d4227de6335a83b6b1bbc45d6e5dfde3bbe15211abb6c312705a2c00bd6dac2d504873a88;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a7815040b18e72182423ec80fab5c44700ac3139ae6eb76be54dea148ecb761668459586c9353de8602307ec1c63f1a9424c7f7ed8fa1d524c3a34839ae60742259;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1773bb0da3d88a7774c665523b4b43a0e8e26258adfe757fb1759b1afba124b889179d6cc119fa1dbd9a1546c342923f28622f354283e25d8b631dc9e663b103c37c9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d8e0e07f854c2cbaa2ccc1b64361e118878c588e8150f319ef96955feecff758e395afd5d0bc6458df5cce19118ae076a4340b0eac268c20e11e07e91c346598f6de;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h106c5abd536d67668049df1e03783a13f453fee637504903c256e0e4244c3362873bd24f12bd7d92989851646b24d4120e6ff59f96f36e12867575a34e8e59540ed42;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h800248ee3a20514e4e5194faaac8a3fb2e67140d9934b8b0e55e7ec60072542bfe501ec425510c26deb6f2ce7ce4699b008f313b61c0e601ef903b1e15fbe82e4a42;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a05644502b7d47e6f1ff04decd8b3151ba5764ed75a759c1db87c534256c789566f504954fb63d43ee2af6301c35be702b1130bc914297a33ce3a6a6915141127481;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1777be45349347b8787f6a0c551dc150041c463d7f3987e226d9abfeae2e9083ce164c5c60c12c5d18c8eed74ea764345936bff06eea1448cd8665f32a24e91285701;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3dee7a7afac534cfee5fb2648ab4bf49d3e0d0d82165c1070c39ff3728fbd061cf278b1d863b1484babb9146de924ef20033ae00e3c980a7a5354b6ee079eb6d1ecb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1960331d38aaf8a574d67c7556302bca9296000eb4d40e2b0c7a4ddc9c58c322648cd8aab5a29c852db94dbfd459f3ae10a630990f5b56d499dbf85bb2985c3d50b54;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h112e1ee841fe2cc035f3704a18be57b9db89823c89de1bb5d0276734a4879c1b46184d0e5131db71a0ced5eac8c03da41d05e90f74c3cefe2d89b0ca5f2f5cb67797f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10bc9567a15267031f73de1a5052e523f446dd47edb77a5b1080997f43c7c01d2719182f7a85eb90352119378d1c197a35ff49cd692e3e499c300629400c4cdedaeb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd38651ee256aaf57a90edc08b683d9538ed49c5000ef164dbd26678478e3926e1263cece1bca4b6ce3e34697dd7a0d11dc9749bee33abf2af7a73593bcc55052329;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12cd320afc75073c83f775417bfee7f6e212988d3bdd813db758322e8d129c5414f086ca24b5adb48bea52e449b971d8360af2ad1dcf6d4afa64ebbb4b5e79d471af1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ce573c30fe22d27f55a9e1ab0a753b33a64ed0f7ae2f38dc0f454c89d4d0f271d71691dcbb0503c2da2f23343abe32df4c7a401638532fb40fe4e080be62f469a015;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3149a5c583a85072502ed6bb0ca58d2f363c60ba92ecabe0f04f10a4009d483106be019eac91b2cd8deddaf2a287c337e42e395827108f3060bcb43d6d54f84f2b59;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1338f4429a3d9974c31f12369a4f8bbaf6f52d13e4cc6c08d234aba5555eccffc4eb132fb246503a30db750143499c6e769780d37cf511c8b149d8d1d68020f3c3930;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd61d5daa5e7c99f32d481b592a58f486b32ce1a65f6b5c9e6f4ec5daacd0e4be2cbf35b173a3cb8f0ea9387d6f72a99d3789618de09655ae89ad5d3a985feef0932;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc8ca42d901c3bdb6f47de36439fdb626bac54e1bf046724675f65c134938de1fbda2640807ae950de9fb96b81ee6ed8d483877775de0a3d673eacb1a3d6adee21bcf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9588e3a1cd5731d8b3f3deaaa992f6d64e6b32cc47ba04e5ceadb88ceccb04d629ad560f328c3a0bd40f95cb82673682c709da6ed8143acbb3b9e2a314aacbac69d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12db18e5b8528bddc062313f199d42c388b772f4a4902967f1d644131cb5069cf44b16b1ebca52066a4a2fb906cdbdea980f353f5461857cbdb5e1cbdd0d1a9cde734;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdef4e7e588d7a2208c00833daab699e57870740879c08885bf7db7b121d593d6fbff75fb46d1d42b43b770116202238b3b7e36dcbad85d97e94cb92dd0e192e11cb3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h58757e738fa8bc67632497727796ce47ea3f624a2a3c214540e008de7abd354bce05f5305a04ef8f107958a06dfa0fd4fc7e59857586a3bf6381f73a2ea0f58b65b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2fd2ba41908eb4abaf848887e6df6e8b87e194a9a6479eec0ba16aad45221924cc14380b2f593cfe71733b612ff9bb3dde2e782d942e0b72ef365768535195ba27e9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105bedaaec7a546865a7058348650385c1baf65ebacf8645bf602d3b391acb64f74a3dee6e6c3ab0f75e7c9d2f93b2e1f954ad16dea513bb01e2269f1d5c14f840cba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha53d48a6d08f22c072441c2360f4691acc74590bd2878d7c45f19e106fe7ee8fa70f9fc36e3bbee3d523ddebce520329e2f40d22e26f2a7e19994602772fe2b65793;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6946174e3b9a39fbc1cf704e89e39c169dbb39c78ddb797d43d5865ed45ab13fa2efe9612f30ff22accd16278ceea5c626603004819aabc1a4310a424fca6894f0e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2ae79337febba0b3c0d01cf8b0d494ee33fad429682e640a1136e68526b64401e77cf1da6821ed7c1c973e1d192c48e24586eb3316fcad87fe28b571e211833ae906;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a3c4358f405b2d0490172e6f20b8e4fc60b2d2c39fee473b9ec7950356db737706fc8df1e43b24b2972e67b7667b25a2683bf357c5cfb513cc5e346101831c211c6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1de5d8d28f69d7778ee39695d68fdc051f486dfebd004cb954f27cc0cc1f29af9a81a66d7c9839bb795f51ccf5d08d0f3771a8850719c493f945b39b5b2a5163d1c28;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1027550a2d6ef920ebaba9ef5816846813e3de94c583398902c877c03f07c924e6032b6398eb32584dded3ac221921db6aad0bce3b4051993881266e9732c5c635282;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa4b2028b49e71959d37c25750e3ebfa1eb0a22796ced69f9e1259f28811f0ca7b79edb914350c7c6c3df726ad3e11ed3d5acc7fb482fa8760f4b0845a8d6e3bd503;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1ad17e959cd4ee488286551f4636ea13c94183ddb070d3afca59b4188a1a056c59d2bf6f697c5c4994713b4937d2ef9530115056603f8dad07e21b7ed9548586aea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16b5573f643db432e8525346fc6c3ab5e8fb48c71fa38e7b3145c5761163acd1bafd9f33dc9c3da4b2be26cd404c1e928c212fb6e6d5286108c21111e709e277bddf0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca7dd4f3cb789a57f29b037fc62e4e373ea8bbd03f8882db6063aad1b809692be38be0c1ecbc201f3783a1369c6cd5988f8b0343123f5003d07a42fe6d8547bd1cad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1428d2c740bc8c6f74b22fed988d7f841ecf1338e5421b89fce88ccbb65bafbe267562a37be8a6308b1c46825bba07de9ee1033cbeba0ebf0277199c2624ff0e528a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a8952b7152562319cf3a9d69678383131f6948cb763223967a44c8baa1f3046b30b3c93301c39466a8e937f6e7e6d0cc01b7c2dd1b8ee9d0802a71b3fbcae8985b0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ab7804de10ef61efdb8a562a4265cf1d7931ac6133dea274eedf0c6341e47df9d0ae51d03c74e7664f604bd79a51530859247b845a0ea424c126de23fb6af4a03d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1de87e1964122034ff93732cce2a042cf4ef5ecc666ef613cd375c118ddc9d3b95fbeb8d54956d2558771fc9fb5f5e4feafdc98fcaba575917ae4665edaba245dafc8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27a54a1f15b5a1f2cf871cf11adbdd170e70f8174ae13e1e78c17a456f2354244dc79f36d83cc4dc9ac3e88822355c4df918695319152f7ec6670870e839c276a1ec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d13a1aca9f6080ef367f18ff3e1d60f08d26ebaaf5a63dd428e38204e8e1e518c0a274ef6ab7b90adde1837d238918fef914411599d7dde34ef952ff43f71b893103;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h134a2bb2492eedb37f5ec93389c98fca76d56d089bdd952229544d767b6944c7408b370a0e2799dfe48716cbac0060f614f16172e536578c63858b127e018625b3a31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d020d8af2ba7f1921ff14da5cf68d50004b763933e13411a7f06a08bf78ed16c0b9d7404c64c2f2d4fdf026cc9618bc2e070e673094718e4831a4421b6a0fb4d159f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1386e958568bb0e9520494c194467021d06122dd71d71291f516d9eb5ee79129aa7173cc130498b3b6d52744740696035f44737b1c552af62dadfdce5dfcb2f327f20;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he665c43d53bd126d86e32129e51bde7f8d127140e4837cd7f33fd6dce0e233e6fe3c307831a0740edef0bf2185a5310448a3567c7f1dcd9a5e57edf08ac4a3fb6da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7e3e0ace2b1e0092aeef8a815ada81e42153ac3515e95594ddd6b4b05499e3898b29554f576ae86dcd67f027f5e9acb44a61d925d704b213144173876eef63e3a19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a96fd77e7588187edefd4e07f05762b47188823eaf6ee17c445a804393f5bd01960381f5bcfa51edf0ae781ccaa1430fd0814f5e5a4acba8b1ac2beebe497c5878a2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12ca0ce727f74272418c37e04267a0b1c47576b6212950c6dc218a23c982e74bc7a44175261617ddd18ca0cc3fe59c1eb0e7e9a5a2916d994c5d6cb2ac900d4a8b58e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12bc08c0ae03da31e2cba141eb5af27d2e5b76f879bffd876d0792c3eca676fefb52bda6d084987b68b7815d9c7f809b7cb3e82e8a2796e013d7c971e2c20dd60de30;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6cae651f49fb1e80deaaf03394e92d91b0bfe992f2e5e55f1604b3c3e2cf9f8689de7c6e509c0e4696ee703dc46b6111a0f04f19a753da1c81988ed91388f7aa9cd1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19e59cee9488b1cb9445bf139fdb5d2a6f2a379127731010d5bb86e91b5090eb3149581c38c27cf656d44930b903c52c0f3e47452c7f04370d21b50af9e5ab738d981;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12815b8e771c81d7a0d3e94d5661de517720b9909b32b6c4fddf94281116dcea35ad7fea64b2e06e3515f7bc3660e71e25ab92996d6c2ab2ca073465d925d647d105d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1acba130897256c1a48c2243903fc8a3b124dd182543dbf66357501c1d83bccb53eae3c41a94dfaaa087650925f06ccd39736dad7f132c03b3599db95f3cbadc70b91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b03861b031c8bdede4ab0084e38d944a099cf17e40b5561af67cc6db09c6aaab583a92ad3cf6795d467c7a93bf56df7fab8cb68922c2020ec8b283af4f09bfe529c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f06d2b22178538d30ee28789ea7e2389f15e224975e3c84cd727e7eb142e1860240c2c8311010246a465bd53f9e98941c8dbd7970202793295283afe222cff773a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ea6abea14513ed79be3e5eddb15f76b1b2b5b80fda3c59803783595ae56b26c319e5f15ffaca736d6d48de4c7c09e4d9c9376322fe5a59dfd12353c3603d6dfc55e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c4f9b63285726cc380c0826d09e23a38e9e4b4411b51dc76e607aa58dd31fdb79c6608610143cf1842cdd706549573d41c0a522db4f232ce1df685817070e985052;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7bacbd1535844ee911f07abb3d3b863798d2fbfca575e1e60bf8502ecd930917af41ef29dcfb6cb408b7c998a6bf911d0ae4cb9aca01551834a1c9b30bc71569684f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haad4ef47eb38a7926289f702d866e3b7a599edcd82114ef4d63376528a130ec391ccbb38223f9a846c4dd2cb7267c5c1afedd2b455e854cd3044da3497c4a08c77f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h21d41a1adc41008cfc4062ef61738f2e9c0c4e1d6c5db6965497b7524324ceb382f1ab930dbb058a25fa321f14a67f5a6ffc43e94079686ace4eaeb43365ee55783c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e16eae6df4cafe2319c21368050f03408add0f71d74fc20a008e289d1e90e09d625ce5cdb993e7e015a82813e38a7ddee6b3ee54bc088140374599a1e05aaf6cb635;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb30f52dcb7bb9b383c2d8565db969f1d8ad9f5720ffada45dfd168a83ebf06f6d4e9d76803281501af27b731153ff38c6832aa797f5a21876fa91b9a4ae83942e88f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha7ae4b9cbd31c316e4484c867dd5f5d6541b6f6e3b810e0fc2f7645f8b5dba21abf9b4e851b1087b146670191c421a61934812bc1e8734f8f6f259f66c134ff03db2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67c38e8c6b8e566b6de702300b785c1cbe63731e3715d88bba2c577f5557c9d83d58a70ba163bbc87a5a68be32747c13238b971566363fdb9268500be2c5a2588ba3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h174822bccd8c997910230db8414855b66f35497d5b346cf14e996e257b73f499d341867ed6abbf0aa4b9ac2545722fc5e464e083278919668d1bfaa919cae436b887d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdf9cb05b74c1d6a855f8eeb2338eae31c06cf9319709a5d48378265338a6a76857ee083f678e3f1ae107683f5c18e04bd4c9633d2d6a5d95e6e7f2d6f48639b81b31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1103c4935e489ef0a54fd19062f3f2f0030bc62beed78528f4320ae9bc09fe632c1c818281bdb7626fcdd2fd108a57e17f8b575a4bc71957464c4f24fff2f71086cc8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab280a24f27bdebb347aac0d394500d529c836c5a98bb6a5e286a59b6c0e000855eed0e57dd3a104363ae4e3205b81471e41b8aaa92cd93e7bf72df3e22855d6e7b6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17ebfd2a8b074d136eadefd6fc48cae1b8fac2099cd1c16a14c4ced5077f4349a5236ab5279923551033b1bc0d5b83f4c5555ce9a9fd5526ef36f62a54d3de8415e1d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17924f2b04436e1dceb866914ef578acdf292822a355215a66b79ae8d2429b3879c3e54eddd6e9fe3ac088d7d5c26bf704ff650840adf5e9e2053d29fc00a6cba4afe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb7d50263a0e48edf103cb0cf4dd876265a148c9a0ce7b2d4b7a1269641cf6735a757958052d22fdab7a59a486841d7dfe53e56928a1c18631b33a2b1945fe0a3b55d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103681aef110b23926d538accc761d009be731b23c579ea36f8a6b2bc87a4dc4185e1fb005a733bc350f6a8fd34a8caa88ca718f7b330f66d2b202d8caf22ff6f19a0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd891808204d98f15fbd222ba3b381d4d0a0b761ab51eacbe467b5dc27b7a2d885c3a9ea34c8da9eefa39c23f5e098b541e08f185fbe46702402410c0d8a0e912c17b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7e9f4dd28a73938f2f0a33e41b13334b0569dea1f8629b4e66774bb1dcdeaa87ac7bc6713099e0dbea7a665e9c679f61637884f8c6b3d03fe89039491675241f765;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cb0cc850c62cae9ed44fd0abee372fbf48723b9f31d6c58017a71c7921924cd1a7958258353ddfc1587f9101c67d5711d04fc00a97bdd864b996772a64f6ee08c1f2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d49934b268c44dd78ab6f1edc75dfa8a4b86d10926b5f83f2b79664cc95216a8b49e8dc7e4a1c443a1f2a31e92e3cd1225ab1a4e2a54cd94fc737c60011d39927ae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc605fbf50423c56473b92146a89694a45ffd9b8c39f95cfba125d833f7f8233b282b85ddb8708a1b7173947f1dbacc77cf56a34cb675635be3677f52f7aedbc39f64;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h20ff7f4c8782ea634d22c3e8b7f406ef99c390b9166d685c7ccc7e093600e741fc4659480daf8e94230b15f772aefea870903f65b66e77de2bf8e86a84826af3da6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2a92ffd19679622e3f710b040ec5619d7f69a62b027b072a16b031fcd0d9395592adb28166c7d1d38d4ce4eebc8d041d1336f0a4cca348bf44e5e4dd9a1c767d5fa6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4dd877b13b3e7109fbe000462207cb42e3ce5b1b7ec3d9b20cb9c8bf0bb7ffa20beb95bdac3c4d870f51afceb4b82bb1707e529694a7d891701eba15953938ede65a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dc6a4a064ec2fbb6e2be6a13d76d89fc9fe9517289c99b94546b37868000ebe2a21ed762861860edbf635017be25a1468061008cd0f8300d7d5eee6a7c538aab3236;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h932d783f5b3e66162dae00a35be739c0a37656a7da6ebfdb854359e39d7d9441882fac437488b3aa89ecb1d766cc6eabf2b3a98c83b1dba45c24d164a79a043cc911;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdf79e2a0f407efa9c105c1f330a3a7a1a0c3f13c465e947cd5264785f8ff26bd0585ec24c2d605044a3e0eecd966bdd095519d6a899b58d1be966ddca833950cff36;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd9a2b5311f35ff14b3af55731759ef4f10559b644175048bff7d075e68a78f0d7637646e870a7eb182c0ced5a52f02f78760e27bde6c9eed37b7e0ed1ba53d93d508;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd8d7d53e157c6c9abb60021fa72ef78f3f770a37691c2e2c20167480abd992ee142946bf1e1acf2c6e22219080f386b996ecd65d7018302e7989c05902619dd49f4a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e716a36dd1363206d66b57917af574ef26ac11c5059716d6606870cf8247dc8f2020f29cac9d243a34085de56908b52db55618cf8e197e893fcc9bdbb6e6eced90c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f7a2e9a623f7f0820b4207d41b2c8e65b012f9997418a6c1ae9d491c54b8cdc3c8feb365c28ab9cfeaaf5215b5fb6723b45eaaec4175b596f557e9983b0f2a08e81c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11316c71c37f904333fe1f2588fbdb3f1e50c625c0447852aa85e0deb3b6c55ad4d3d3e98223d6a764f3837e0e1564c7a39f0cb9d2f4d0cf5ce4dff6fb2d369c40cd1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h94134e0e50a8c890a7c3793e8ed1bbe9402f1baaa5fcab98752dfc4ebdbbd991e57c698cb1ddad0c1961c48be8cf6a24d1f1a3854eea2e8f860004982606c3b07b6a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4783e581b6a492e3cc60bce0b41b2b9d590393532abb544da94e18f44bd084cb7bcb67d23ced9cd339ffaa535e8c1990aae435c2ce86926f2d5c2d2975078e37808;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4fdcd8a2ea0eecdab8385d52906b8b0bbb1cd8c3b9265a3d110098f626f7167c85950920dc6a3b93624194c7e9b587bed11eb8b4c84c97df1016ed8dbd5c132978a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h313d08fd0d8b6910b3356de4d0863f6c606be58901e73aeb0e267c3d274a466696a7d0349f0b7a95a30e236d445d369f000839be04631c59e812d8dbcc0ec8ff6cf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he8c901cbf2cb551c4bd3bba4cbfbe712b2b37db94bdf75c70979d9f9bebeda0ad85c992b5d529d5459d0ab3ebb0a30e76c437a964c26c3596c60df940194ca34ebfe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f78e412640a62c80d72f3e18fa957e61fac6b7e49836382ec844870cebcc041dce52607f216a4ef2bfb8d4264feb83a092ba91b3c511d136e0545991afa98ef2b91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c969b20358bedc575d12dbc6fa456d77c41bfa17e9c3d2116630945b76a2702f299f36a86454a72d9dc10acb01f75ed17526a3e1362cba3fdd2ac38cbe380c5e8f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd1ed2d56eb0f71834f34e12fae46151b0f399ba15f7dc2ae2db661e1f8078b8b285d4c607f4913e736a6f91baa3b81e3a5a05e065b232ecedbe657e864859c783a23;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha81ab4d9fe41e7b8d9f8cd642785a7eb6282a9710a6b1eb8667b6403b1de99f0b772badffb99280e3bc0638e2321784a5eb2af04610aa74d7bbd9f6b228282f84427;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf1ceebf76de871fc62b2e2c060e453417f42b3b27f092e132dc6d7530fa9b985ee488222c68e025e300b4dd8fd930110d0b7305c577b53140fda8af55adf26b9d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1846a2765ff68e050786549428459891994670b616ebd17c49c7e33025cd63410cab3144eb38fd16061bdaff5264381545dde5ce90adafe5d0db8886c19540d6445cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af1bc26f409f7bdf02a563f7173e5992782849af35848013adf0fb4241ab280787f805c8d2d124b227c1b121d425eb700cea3d08659c1179be7b81dd392a65bd598d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had6faf842b4d535c1e24d93778122f9d04a9b17a19c6e26b1a0e5121abcd0f7a9fd97c474425101aeab1a94493e69d26263dc2c4bbcc99d0597dd583e03859f05f26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ce5e474d036c7127a9e4c4f1464773a6d15b00a35277371979aa4df9e66aef9d0f17fd50205acc8aad1f910f01df813607658e71277047a82844f96d0a00dff72ef7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef7b44fbc89ece14718dcd1480be9516af5ebba4e0ab721e91b2d01b1bec938d4ce7382ab7a8f51646620a7e51d1aaff7ce219de35cbc4e00f58ba3985373082788;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1785f9c2cd1d784fb159e5682f370d6710a93a849bf592ec615ba46accdd53c3977bc5c9f746ec804875cc5a75e5403d0bc77af696a851b678dca7ebfec7bb85acbc1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108555bcb13115cfd8554461fc5828fcdafd6707f915686ed3871e85bb33eb40643db56505be549eb17ffa8bef4da4b8acb4ec8f414253988681a88c1f5c5d645261a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e8f9b43c5600f58e5c33897aca9a6dfaf37b3980ea956f056c2aedc47ef63cc5ed2969f7dbab5b2b69292c7f288b8d0f69cf5f707a374392cfe7f45821c95bcbb809;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8673f8526f748b4c5588549b7ab0e41b8e41d25c2c05a76ebb3df70545eb22358580155cbc3939b8dbca84f9da6ba0087c870e491ba7e6158dfd3d10a334a7c0cabb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9bee5b4501b25b3ac65b8df61246f75c95d2beb2f080782cf39412fb7bba53764d7918d6f498c147f3fcef894b40697c1debfe8a463fc77a49e07e5ed3ab576c8337;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16adaff70d200b8439f0dc7f7312d30b3a3d016448a3fd98ceaf8ea3c2ef89426ba0d676ade809dabd3cfd952ed6e01771c253e65f5ed4c98f160db6c3f75a0fb8c0d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha617cd8c3a306f8fb337f858b29e669b77bd5eabd44d35bb72eb6d6e6e58b03fbce82aeb38cfb0bc51ac485a4e8358c9d46400f17ee4ed04e9b03e6fcee065633d5d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e9798ad0267b268a4d66d44046e0a132df366c4ad15add79ee8d2301ef31ecffa075ba2376b3a909db3bed578e2f2310f0265b739c3546efb927cba7dcc4539aceb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f1020227852107567d29824dc4a14f27fae624c7c354f11c5435f2b59f32acb8a64e15fd4aaf8c0f28426ebc4bc17523513450fcbeddb0d13e56244112b446944422;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101f54d44227505212ef62308d0cac6bcbcfaee2637f67be9cd3657f856eef2bd262b858790e3c81cd022693e749d83230b50e468da4f3be6745017e3ed99d61e04da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h836f89298e4a042f03aa834a121c67ed5ee9aaa862644b668705390907327c172eca2026b07e8cd166bb5f6d48b3974dc67d1e7ca78d2496a60e77b83f5effd7480a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b312a42f92e7f8e1dabe9c6124a20b5816bd4a48f2b45a5044f0bd537e735f84080ea1284a1990e439770e67baa8cea83837252f2ff1e559baeff9469c10f51cc8a0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d764187c41cba0cc09b253203757f30490f6ccb2a2e143e5b90a1812c51a2fd2e5abd48ffdaa4ab61f937f0308c1de00b96eb3e60efdb6c0c65a35f8cfc08b8b1c2c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc73c430fb02eefb43eb2e36cbcdbf3b59cb661e07e976bca1ae6028d85e5711a9e44068350767a3a945e4003bf302006d7bdbbfa5f4e94b5f2caa47bd35bcad97d4a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf8714203d36f1dd69943b6294295be05177dc8eed8391681154d54f2e7d5cc8019d7cc3927d795e5c10b6fd566c576a133dd713909a8ad2123a2994161fb763c8481;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190c54fadb4e140dcc279aafe10429c3efe28dfcffc3f823e9a7d25e6da9584574070c9dea584394478df4fd578172d79dfc578d1ff156d8b489081083dd78c68bba7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h64777d60429317bfad7d20650b542d514a0f3834c90932ad9fa08728d00ea484159cb684c86c62c2651649f7db7dc0dbe9bf82ffc6bc9df7f1d122ff7f87fc05a262;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3a997923381d654564a672ecb51b2923f2602ee954b39ba2409d9d4bc821e33322503fea5a86f1b9b78a9300d30dce56d9080f8c260934990151d6faa4d9d6ca0cc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h574bd4a10ca31bc66df442af3dc546a847cf1ef150b6fc26db8ce07ffa4fdf8bd565c8571097dfe28e1efcef75887d0cd109b22b3a26899d5fcdc27f89cae0b3f67b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad3bb1767c1eb415e62be5a42c3c436fd7feeea68585f3c568d97cdde86673f9b82bdeda4037ca2dbe40dbcf8417f057618d2b84c843cfa81434f649ecc92869de91;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f393e3478a7e47ce5cccf3c1cab56a6193f88aef31be20343d03288d573866d210a58321242e1ced20b975437f8d3acd1697bb97884942fd5c1499ad7cc2109ad47;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28e63e66f93f1a37be792ae4b811d5381f7a8c23ab5895547525fdd52b6cb122204ae32c1423b2ccaa41a8f617b2d5b376a99d6f1cf6dbf218d6971bb22eaf5108c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a866dad98a70bfd1c6619e55fda73151d2061f9d96ce2e8d63626eb105290c8e1d66175b6c0b14e16c138e4f8cb1d1b80bf5a7a690073b7682abbf40566070dd86b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hecb73a6590d3fb1a5078055d8efe212248f4c8caef8cd16cb3fe81ae7679535a752e638928e3d1f70bd5515765538167840e446df1825dbccf4d444867f1804bdf46;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf61ca018010149f2fead100d6623f7f71c055ba42061ab58e98d70e78f8d74962611ea70ec721ecb19263394826bc3e543a603164ef73b0c52b53f612c5970f28340;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h39d5bd338e2592219c4aeedbb178754fadb7341603d707350b7f634fd6bccff4d1a60ab188cf182db4b4421e426ebf80d0f3df88cf3e60a5a0eb45ec2ca076a552cf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h199b00a511453947b7dc4c02faed01bc59928c92200704863c684a27a780da42f988cc96050ae925dd5927e6b91dbeabfe5ee9781c74922b2b164133061781ab44d34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h30224fe605a0af50f6e4ebe15909b775102efb72d70f2429fd07808cf9658a8f0d020e48213a2fe2e4ad79120f00193592751cdf6dea5e32eae09c2fa224b8640405;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0f9e81293f04975fd090eae5954b648c7f035b68950f005274844b1e0642e41ecf1011502ff544d2b0301158bea436eafaf7768dce996fffd3873fdb66742421eb4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa4dd815699570b5733af41a8d03122d17143f9738ad3d0ed58d4588a67fa87f7066decd31a4e7c835a6c65cd5779bd937f7fa08cfa549443ad92f00716b51160f5d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbc45a4101634be01c775740209b819b73a2ca5ec1184821ce2f47b8af52b56cec5b8d0bf3cf1d80386b54e1b3064fd39c453cec583cfceed1aefd8128b4cee741c90;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d6ac4c0f5f32534d56de2ee6fb2c74a2ee9935ece42d44ecf9f9c0c0199592daa58e240db4f0dfa365f54575abd043d854755d4fbd9cead7b92208f389e28fe7d83;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d1d6c176ba0bf8e2896be86bb223e3e1a77389987dfed31e8e8379e1f75515b2de29d042e62ccae35a2f9c841d5dc5abd0bf8f6bcca9aba2ffc34862416981ef70c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a5ad0547cf5f76451c64dec8f323327094c3a9fe5f384409eb2e01be1d4c119919fd6ad3590025c84611853c12c7d9ea4c38efe2d8382fe2167f82cf03a6b3308a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e68f8b50ccde062533fce0192c06a2a10d5dea7f9391cc7260b7dec75cb2cfa2a431e4ad39c0743e766c7a6764f2b5de650907912e89a07444c7cfc5f5ab952f0e1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h107aede7579e6a19ead9c9a1a38096f0659ee74a6eb954cb10af917fde613ae561d2637e215b94109d55256da836ea6f1e6756a5df3b424b70522c92fe96ff5220ae9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h95c61e75910b5beb8bf36252124abf1ee944d3c82aa2c1824a53ad87e80a628d4b5ea5100ff7d7d0313212af75847d1a66edea9739ce601c07614def3baed874faad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1604c6506d47df662da0ef8792824730e9237fd18ea17d7f3bcfb6e59b135b914401cd78cb1bd3d9eadd8808f340779baf320c9bb4e2d093f270c9e5c0031e248e188;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h174a9c592bb69f00fdf99968179a4b9911d619350ba74195c908158b7b01e4998da4849c9383f4b16e486d984c45125721ffa359b1a4ee65c16fd16e9e88b521579cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d0c2bd1612bcd90fc6a8ad40e7db5ba6c27b38e51b0d68473d7b78a066ca477f9eb64a2cc2b0daa3ac557aa3886dafe6ccbe1aa064ab4dea2689e7738a6e54c8817d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37076a824caa15f6350abee038ccfab7283decc59dad1dce71ef7591f2a128e6133850885e44708550af99cd196cf25bdb1fa3231fae06fe76a00bdfddc78c5ae959;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dfe70acfae68bd7d99b5093fe8599ec867f3af57c1b6f68cd1118eaec4f3d86ab444080ecf25dabd3e164c90593772d6acc88872cec1d936b7a86f9a21a1157d17aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b5514e0ad44b3ef1e9d1af9a595b8c6518c2fe37c6ad47d9f8ac5dee4a3676e88c4f5d95face13fdc0415de6fff26f720ad39a98e0cd37705e7ad25f0bdd4c6ca57;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6b6735522ec05a481f55096a5c60897702bffc152624e09cf11dd93eb95cd295debb89459ca07fea2baa3a27eeeaf92927e59610d7b58238ab318dc507c28f4eb8c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16660219b751fe2d14ae4b6fe5a5345a8ef8cde4e8cc5751d6109b3b08135ee3bd8d28ed982a484cc998b28ab612123749fe6e4677a8f53edc44e706474958541e899;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd08529567307bf5063b45c7aa7fd684aa509de95671109dd9e742b2e497ead602bbd29e2f30de6150bcc448b0fd773f29e8160698aa5b4419d7e791978557e373602;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194ef4d03ea4434877e94d0e0f255d663c75b6678ca8e2fa89ebdf6c64756d1268fe299777099a8b36a7d0389cfa43bf96c607a1bcc00c711e10cca788cac20f07f0b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e91db21e927918af296caf1909028adac655bd9ea9ac0e854d1ea18f76adbb8a96bc6ef760efbf009713418aa96784487c9e4191aa9a6707e5706776eb7a0e865d6c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h98d0744da4b05d9e77bc84ccca6c495ad2ea351b946755b9c0ccda3c23e4731d78fea7cd58b55dea22b166a6d95e5e4b04145a6b5e11486b21e6b6a4ae41a46b9aa8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h185e7220ab218f556b09041c7146df550d1363eb719ef2f9091b3d355a6d3a75afdb6c5e89d6ccc789295a5399cd66b0dd425764abb15120529d01c7ab7d8f57963ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12685580e37cf82fcd3062edebab6f29833038e35bd4b9a88b010cf7a8cd2c7ce23078d11b712fbffcbdd211117f425aa045ccce84e84a80b18a7bc87bacd09c02903;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h176bed72969730cc3d22149ec04f50c0e25e514983053030e659367f00d9250c9982fea3baf8870769bf2ca09117e056ef4924319927b9971197534004209e8ca547e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c3fa8532bf5986f576e0fa1db9fed3ff628bb2495db83151ab84ea56ae19bf4da2a877944fb4dd5f276eb20adc62bf5a494a9c5d8ef9aefce784fa6f4380af78364b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14fe58448ccd70331ebf00dab65df04658ea6f57ef3cba32fc3d039635537d71351041e12b80940aa98dd429979f2e44be83df3c222e6edac3029a5164ac255d4531a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf6a67db1046e31e3c4b2dca5fc1a3a36c72b3f0090ed3143c3987a231564adca7c70affd93d913baf996465bf6f514547c8faec88e7e1bb74cae0f020d595f820301;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12daede55868791a2e1c0c2c03e6af48b686420a8d8d1f3d78c1281bcf606bf12bfe17651937ced857cab37c7e752ce14589a63eb50f431cd69e463ef11633df42de7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9e7e41031aca01d73eb5a912535574c912a272845ea6bf461095f151e424966a9e63fa71aa5b00a379e136205838ed801c14908c03ffada1d3615b858373a8c694d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd0c452de8458c3954ee0efb95ecbcf5b6f45081e6871f84d8581ec9c183f42446ca18a13e2156c28895f07e0eeee79e63356b903550f4c8660f00c6ce5975e852fef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a259c4cb1fcd0ca7dc1cf12f2e5c03a956ec11fbb407e6120dcba2fe323c4a8bd159cab207ae73e09d14515cbe9cb5c7aef1438564520c972cb3c00f7b27469c035;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hec92a1bd7ffdcaa30cf189790ca7cb2eed88895c98f4c458575eb41142e6cfa7e3c76858c31e47d4a2f0a116af0c3d468f38bfcf7c5fda87db65d812f1e4bb005a9d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h365819e2835a9a71933228369da207fe65b248ac0c21c9be0e50f2b64f143e173f323b469b16ea56ebab468bf6204dcc8a67286af315bd129de71e7b8f7ae86f3f53;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf501b849ba90e35a5b82db0130d88586a13695f4d5736054e1afd7d850bae68362a47d2d9558ec8aa58d99bff06f45eb78d6788b0d0e4c6fb9079429fa52b25a61f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f4bad3ef7103df45e9d6d26d7cc206c0d32fe44a72ef76212a011aae152f7d7098172f35b7379df323da15ee1464a726cb430f857cbe315fff9ac45e2f8c136a09db;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h51c6c4b53025a068cd99728217a4007d8e72f37608b3afa29b4c3ab8bd06e0bb172ae0cf64eeb45c8ca2756d666092d17bcb86320b463688f694f6009671436a1f1f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc5c76bf4a887637714d9b2906cbf3c3a934b37a1d1d18c83ec18d18930467ec1ca46fb7e0375224c8c294e2efe420f6e651411acf00186c746346781d708c681fd7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ed7bfadf13baec4a2d6c1bd9ece88ce9655f951dd962950d010b31f1d94700317a76738ab05d422fead528e3af4a4e6c00009eed56feaa7676e939768acf54e2bb4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4b2714773ee461064454a90232c68123d8feace70bc974db1515b90cb60ebcf653b656fbee52617af22584392008e03951cad091d50d09808151005e2a63719c9500;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h59a2b743822889d07a842cccc06cf2ee27d11c665bde680999f826f7f4bf51f8a849680d0f34b46bf8fdcb845925a49840130fd3626717dce55fa5e32f159d1c669;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h159935117b7cbd8168e26f384f8e525e19883e8509835028a63b3edab94891f2a19c28e93114672c2f654ae40338baae500135475f63c87a7ce450b44508cccc6f9f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had9e83d8eb9bbc0d34c012e8a67d5a885fd8789bfda42e51c4dbc48877bdc4e6bbfd5dff9a7b3085e868fe63d07aee95a1c8223d09c7006e48143d60c422f6a37fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16264b1f4cbc3d4a5ab38f753e05882a0ec7dae40b23510b4f7f7727a1e0e1409a2085e7846045709c723aad82a57a9358407c4707d43a27e2006f4711e0c865569ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd0329921bd34967fa707081c5635f0159018cc32a62eb64408e1dd96632f91dae28dcadb4bc84da977b15ba7ad6d3b4cd29aac3d0e341e227904682ee9a5261fba3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5839f380cbc1d786175426b5a66fb99da8f1c05638fc1d7781ce7fedf86ccbb17d2e088dd531bc37657aeca2546a0662e29567644115f8eae2a5f20d46f5784835a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h785145458ce4b7ea57fc0962eccb4607f1076d579a1591d15d2eb83aad14f7c4bd07de13240c59835abc5305d630972e1275a6b45ed240a799ec84a5d1980bc61add;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha415b92632a4fe73ae60cebb43271dbbbdd94c23ee1d05aabb4f953770dbd9af079b3c610e6d33d4b7bd624dda9b341081cea877af9902f76c63a250febc0543deca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb27a97b6a3f1a68c44c688d90e4372c8c5deee6888f225375b815c0790b3d6ce1639ebb32d8cffeda7cea91e68c0554344eb17513042c9b30fd1a5dbf5f1d620428c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1180d40697668eef68e37040167c5f44357ac5ba43ff3b7d469aba80b3519078f1ad470c721ddaf8fc546e98337e876ce50522cce856eb0be91a34acb66d89de6d30f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a384134dfbf9c26c940c1018e94b8e8550d4de96f6acc2708e7e66067f3a1a20c859ea5783964b57ee2d4d5944b1b780f5b3e319b2e23ab60eb68e06f6ba2653fdf2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194749d9f5d0c65751d1c66575a563dcaa6bfc749f76090264049c31e609a19da1e33f05bc49f68e9181dc42d1b6f8fb339adeeec526ef5e5ae7c5dd32058b4caabb3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he552a0102335dc6e20e171ed99130cba684e6d9f5cdf655e8cfcd18a8045ca31e87252385f8ee53ba39c8acc2c602eed1c80b7c63fe0afa5115c86643356e9db8d07;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb27e52cb090dee8cb7050bef0fdfdd99a5603dc7b646e50647c7725f1518475e891b1146ed4963ce10d11c7ce1c2270b7fc06155a9984850611cc2afb3fcefff24b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1862a30c12fab654c70327ae30358096b7ac77e7f2c187344ca49fadadddde52f93d66b15aea63a4123ee864de516dc774afe26a2fe45890d69ba7c7d6082cd8bc964;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8559ad8b8686a34c5b0e333b8ef182f8fba2d73cbef4d8db451d0b21b40be4abbba5c7dfec850498c8d1d6a751e9ca18606c8cc5387c47ea65839cf092ea14c1fd0a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e8646d3c2b9ae7fa292717c6a703d2b53b9c56a410ab300628b03fddbfd8b65b1a98b25e07e7202e2074cf8c4554d5609035afe7720675796b4f5708cc80a419d10;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1011ee88fab3a1e4181633e866d2b972485546021e2797e560bbe38ec8a8d937dc8cca7704fc32cfcd4188c13159b4102503970cbe1e521ebde52fa40c99189a51686;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c2700f89b8a76d4f6a7fa5ebd8a149859dc8f942b5fc107f60ef8f4e37f6fef127405a8979fbbb23f7f7a41213580c3eed4aff890d50f46ee3571f8ade20de8294f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h94aad96c6fecc78f3aa94f2855add9b1df7fc2ef09c7dbc582aa36bf48a84e528c936893d4c2414135f8235f6e0bc8a507d13debbdc9cd8a5296ea55d5906bb9ac45;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h459326a923e9b2dfa62a4ca626adce742ebe1f830c519ba09455beaab6b92531b5bb73fbcea7cb3df4daa9b77a2b5c22d159ddaa215342d36b0c9cecf2c62f6eaa08;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h172fdf11de0fc8f2360e67a68cb4cec94bd994afb9dc7b04eeaed4142d0ec6ea47947cbe9e4c8bac3a3e169cbfda69ae5cf350e01f887bf86f7e099d410867b5e87fa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haf144f22a00f8b72b179325324e152c68d008f76fcfa1c27c2cdcc9f27ce06555ca6bad0d877fca9c0af1344dee52346836121e645fb04655e3ce59426bd7de2c1fb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c1c08426f81c92fc3c54ccfa7b4c00ac63ed35b967c70345f1e83a417150cd33576546c5faaa7e912647577d79727f026a009ac57024d25725af5aa881fb72a866a1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1844ce1f43a1ddaa7036a5bfe1e53a8e91e2b3dab79a25bfd4386cf2754a7eb03fc93655326d7b39fa07805dd438e1e615c83333d926fd8ce10e0e4f6cadb79350f7f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea5c23bce7d4ffdb48ea1b42c5a6aff3628762d328be104fc6b83d6e0d4f24b2efcc681da5c803ae3a680a7223c3e27b5b357e295857d38d3629726e54bc5584be4f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h191d02a899abd8358a3df50ff3ef657dbd75e997d198709937b02bba85af93917334c7dbaaf5b9c612c521420fd141e184f1ad575982cb891217640f4950d276b5320;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h480cbe6a3577f73e16e76f3b1411b70a88801045a458a3efadf791e1d75afdcdaabca6307c1095b7063a9f5fd2fabd9d7a26889d35a2013ad13bae052da05887b462;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4de2446d49ccf65cdd5afcf11137c26ac305dff9d4b8c6094bf2e46842fd5641a90c3bab08706e3c2e18966fd2a4373d2f3863057a5f10b793143763c34b99945c1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd5e638d306bfbd4f62f647ba3bb0236e42e909f6e7c0f10f7764ae6239bbad5c5156ab70ed64de6f29ec1e61ad7cdea971c0696a57cfbe60f60abf68fcc564b3c71f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h117c0bfed42a628291b6ec08de14560ad3edcea8b87fd455dfbd497b335773112528cb74cc4b161f757c0818b4acdc6ebd8bad7030bf9d2d1988f276a135c458ce8af;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e1a08f21be2da4457e5c09f3062afb5d08e7244ec9a7f0674e29b962dd517b7771187a1e0254da63456d9570cee8d13c28a64d08d731fef7d40b447cd0d4d7ae956;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e0e15d55a6971a5fcb2dea641d5b9600697dc2c2642616b8e9e466d624980a263a067057f6108d9dc55e59189f148ad4c233e87ce491fceed7cc8fae254598607b8b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dcc70d7ac992fc67c40e57f563d5e4360e114208e8aead27b3e5cf7396a52036c7a6baead6db8cbfde2546fa9ae80bf65c0eed351853b084910e9166fcf39a6ee03c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13affb2ad53ab2a033d0907e28684fb66b6decd154dbffe3fc22d6689df299829253020ba1f34fdde15e08df31a8595a69e2b7caba430726ab5d08de11c484e60f980;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19aab88a13eeafafac19db0ba5065b33d7cb586f41d0fe467eee591dd1d2d99e8ca139017b8af4e53775330511db5c2cf56190a0d07277d0369ef7efea61bd0a8077a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e95dac67ad1da442b6696ddb402cc8cfca54b978e738b662a6c7e8ad24d0ae8a42e6aa94bb1ea79770e5f3c1dbfe1fa7993b84ccf26de8bd5af5d267dee90824e926;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ba9f2639a6bff20a8e2716f91a5f7a4b38fd14f383726baf1e484d75f46a3a2d4135aae9c30a0dd673569bd68cc606f0d1e670768f820e3e9151eb37f7da6e63c54;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h199ee1311e62fa094fa89e295d47b53df18d38125b75593cf71618c3e2b029a9a2af1cd9b07b914f0466dcad38b52672f91d56a67ff13373c3e99c1ae2415f241115a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1088925b8015abc46cf6c5407ba2c20d41930ba6b1e7730b4ad414f69ab80b341f4b7ed8e0235d6debeea669f61e281d70cc09268cd68ada0a86f206b4d334fd623e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19da61fba7b96df26aa64496e6dc5066f44244045f4414a1135c7a97fbeaae15d804f425d823622850666c98c2a01a1f7da1d3e472e6cc1fc1de149c6541837851314;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8f62970e469e311879ff2da5e2670fab111de683475df052c58f384c5fa9954beb4830fd384a63226fa5d7b57cc9a58b2a1abc084a87f27fb379d4e4e00969be268;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc22b55e94959b68b5a169f92a2a6fef15caa60dcdcd565f5d4e76a09e9af8921c0ac5e99b2eb9172872d0558c2d38e9f70d5e11523e2674c8b490c70a14b100be2f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h46bf474f9524121783bba40b3f7a11e717f9edd544d175ad963625059e68b0efa19ffac9cf9d5038e6fe9139dd8c1650ba2e334642acd57c88b6391eb3c5b1b41067;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc15b8e3aad1077c6ebf976a9c89a78c9d9f14ed3a0210acad1a88f68c61c9c327ddee631d95995194515c38aeda562b0f5ce6e4355119d5972278094a0197b594577;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12bc6a881325cf56efd1abb3014fde8b3ea9744888f4e34037a82e19c33532b5dfccd8905afdf6452b76b2ddea3a0fc7fbb1b429ec5bae610368afd8ad5cef9a6b764;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h166480e0b614cd3fc9285747f5ccfc941ddbd132b09f00de783c1fdbe1f596044eac970dd8ea468c96a9ffe3fcfc56b35e85c890cf945151c8b01484227ce529a5b18;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17fc6023fe2082c7b508dd3002afbc35944661f05bff09b12e3972e1ba9c3c994db74b9ebadf11fbd98c0ddae5de0a5c651ba9cb95058c09bc98b6d2350b2172f70ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2cd6933b875c4a9e62009c6d131933b6ddc339112e866a0d3df0ac1bb5fb8514c224cd06d66ceff62463304bb8904be251f584988d7328272a3241ff58bc262297bc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1280261a0ac8142cc15813bb1f9520ec5619526574c721adeeec34f428d203c44bfba76d8bdbe63f9697a1c2e735af394f282c47b53cb71f0e9dde9c0cd53fbc304a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3a8b3a37e6587e4297bf83bc622015296b39ebeb6a1eace485ac681cc70158d822aa47427ad00599f520aee9218de60be5be5a6bd4e64ad0de89b692a4d90d9acae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83321c651936cebe801b6c94aa54f894b74e3cfbce2e876ce8b7217054381745f6b68ccae074b7dba4e9c16d74ce3af119d4b0652033194626311a2653c0b967fb31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd9047c18d4f293dcd7ba0b0d09869cb12ae03b72786946375aa38426abee39627788e0742f46c9b054629bb11135b0a6d567fd33f839e6a6d3dd12cbf0a98bf6a701;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he664ece052419f0cdc25b035fbadc6722e65032312333211d1fa5bd3bb72bec53a21794475d995ba1e4d2a03ea5ddbdb8ba9b716e05a91e5d37de45ac7500e10a3c4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h172d1c850122e78538d85bd96d9b19f9824234e38c2833a86b14430d3d624b0b97650dc8ffa4766936063d7118a4296920fb689dbe7677ce69d723f5b0914a30962e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h201eefcdf1cf6750c9651c1f4959a2d687dd91be96fa854bcd52e3c2e5bf7d9f37b739f88f8f0e1c7db0c7907d64dcb1053ab75ab58ee9a5eb6a6097265bc0bf1a8a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171d510ab511d274f3ce55f1105c0bcf9cff135b64fc90b7544607d44fa710430ef60d1d900b86766de7b11f6dc7eb86fb498e05bc997395007addb7a97db44781099;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c78fbdb62506c5f84b08cf1d2a61ffb3aae837a085dfaf497d8b58d4b884e0e0b72371d4dc02b344e3dfcb7f229b5b3d7fc35691c9839c883ac4fd212099fc13dc0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b91e548a1ede015d3e7f5267548c84ca80758e09dfe533cb76e9e037bba6051d56a77be00c8a5966d533ee1a53a5c02407ebc841efb2b958b3ff1d10ae37ba93e2c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aca84c8a8880d415a8fcc68dc285cc8247af3812fa64dd0116e673b9766a11e0b9b0aad76c6ec0e65cc7188599d4213660edbc3dc25efef02237cf02c92a14dcc909;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha8dfe76e6f251856b4859fe49a8955dd634aa09d2d6ab5aa6c1f9366f477d73f09b6ec9f6221f73555e4f72fab9b9ccdf7b48b3160985ff7909f0df89c9c78e74b0e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h860050042febe27e67bf2014679d402f67c120113a3a33f547563b5fc8497802c469689d04d37293fe6e08ea7f3570ee8d066af1e23977cad3bbf777c70ea37c6b84;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6bd40641e827476dc321ccd17d556165efc51195426a1a66f461892ccce6055c0f67f93d7caf97ff6188259df8b2fc7df14bc5a75d7ae9dc19f1a0239cdf4c96f241;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h924a85ca395a0a5a15b02babbdcea6b281615e5c85cbacaaeb8db51bfc5be7ffad9a2c89f919a582de643940e5c9be51547a261b7dbdd616921ef029af8e8aadf83e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0f88319e0a5a09b93eeff338455d270ea59d7e9c92af989c52c54cc9df49c2058eae00227b2f309dabc0db15004d6c48cda52553c387b3741a53944f65e64743fe6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d6c19229e98011bc3af670db0437a5b386b31da8797da187099150d79bc55835cabc9478f78308a15269ca15dee2a90fb21b2bd617c19dbcbabd2972bfc51354649;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18486f1c342d51e5d04c545e9cd000c35ec78ae68816ad511e8d7f83a8676ce002f182bef8e57c6421ee8ebac786f30f005bd8fb3ad95ff18237bd148ef25db770d5a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heaf80d89d531184fb4ffcd2bb735ba39c90a3db3fec12348b0205151fe0622e07e5291c99bcf4e10c14984940c9495ca4aadd2532385dce4a2b2e011b29a011d6a85;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h95cfac0654a8d26295002f77dc49cc784be7c60bd5b84cb0639acbeea279ab5b4283f4cd20122f806665ec9e834be7568ba6234ea358acd9a9fa62d7a6ff3c136968;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149510aa88f0a95e14fe246c20d9f0ec674085651fb12b227b40f67601fbace6cbb8f65803ca41a9165b1cedc04e15a1a47cb80c5ca98625961dd6be502e456b130a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h82dbe038c0915c032007d9d30e9d01bbe68d80d4aa8034f44482c35e008052f0433212d9085b1617d498d9017b0baf950a93e81da4db7823348d2edcdc1763ddb82c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13212b0802ef9d7408a5d5013c6e6835c57701b813c06cac8b43c9359c6397162f6c1d2a794b8883979a2215a309bc8470d3b8ec3e8747030b1a6c977215ceacced36;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1266779c961aa3e8aa76f07eaab22224321c66222ef3cea0830149f563af4bbf3b4d3b51d05d49c07a3f53d2eb63100cafe94bbbe8f0c195b411e81448621d0d5ca85;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h68af34c4a0a63eb363c2ce4e98c030b85f902ff6455b0b4eb58364a1e3e417a978c1f40d12b648d52d3dc478af61a7f1d784427aa3b90419e6462e6f2442d601c06;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he0fb531349c7dd7932c2c04b758ffc8c6364965c09b15ec01ed89d59182d046dca8f47272ee35ba9e925e52accf0848b35f7712d8fdb65a13a24ee520c1c2cae2626;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfbfff4821b58609906c6706b8ed56db81c1f72af3f99753fe71c86cad909f2a447b042648086610b09a4c69e2879c716353bb9676018c5c35d9be1e5eb674670fef7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9466556d94767a1c1d0591c1467f13cfdbb189fafd7f95562bcad1d15a72becc3b3efa68797dcb54630d4dc0086d529bb8111a6291038eeb564c6847a3bdc79e30d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16105128a42ca8651cf3e47d87c3fd805acde083b3befe4de1ddc788cd265a8cf86a515e04e95dfae5d989a093d0891faf5b641e2641bf0c4b60891535917f20f23d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2265a78862d8c2f74ce0391f5320fdde506e70ede2501d8ea30fae1c6e522533a697a32a7ef9128a7665b02189d30a6ed267f4b5f01c184b3b718bf879f07caa4dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cee3b089d7720b9c70cb2e7d44dcc43a7d872141b52e5873efd1b699692f3507203687ef4754e52693359beb6d311ad43d83202d4a6de395a832b178db201e7ce13f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ebedf2f9e29b2ae7540afc2bd1639b089f56baecd12d19b0d3d41f54e9405babfcb5d14097420774eddfc844620b5477b3beb76306fe49cc84b02f1ce91be00a93c4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h113e45b0a9fbf81f526e9fb4a948ef4e8a6da23fdad3e97380f4576b8fccfbbabb40bdd6d79f7910f3459d6dc767bd741a71d77e873f8e341c77c0a3a99a2e03cdb17;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h115bd4043f19639671b4280d7868da451ad4f89bdb63afa620cf37b0f43a7f445a2838b0b1adc2254f90442bd8269e0ef6fdaf4253e6acef40721cf8d50375e7ba214;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h29bd4c1aed91b58eb4c2cdc3e6a54b59b7b0776b864555080f1b83a5e130dca8c6c061ab7c26ee4d462ba7bec0d3e8f3099994f1a0a5b84cc7bec82afb0806c5faa0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e1f8088d2c667033940cd2e81c9d6d3b990a18f4cec4bb48bc175d7c457a4f129fe9de74710ad10b2fead0370ae20d5ed433758ad843f7cded57b9ce0e70c182e274;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13bdce24d311494a5c3267cfaaddc4c5d8a7f8a57e1bf656e9be06d00511548b8e99fda99772a3f3d70cbb7aa4db3019734f50ac65faaa80d9cec0d3b5f9d3a2c182f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h65e15ff6c028b6c120e9280acbd0b84881439de07b9e7e67061636d52d749c3131b73f04089e2e52a1a5f892f46e86aa7ebcc4b47a6e9f19f2782a4f6ebbdc56fa98;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4bd86171c448bdb0ab32e5bd617a828c4ccf375add74a34c21a34f7c543e05fb5519ecea51f188b2f2add2fb76d3f179c48ec0f982ec774d305a3c6f9c7885d3394;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa695907b19d23de15835bc4ff393aa34e182a137aeb6892a6b1b52a17440e882ac178e45d87de638a4ff5e6a75358a6551c7d413e633b3dda75a853af78205f773a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h650da146a4ebc61e3410a7ed55a5a1232485caa0e753278268fc523989ba413186ef85963104963704b1afb4b1444ce4f9a7d70069a68d95d1e11d6cc1be7d1aa73b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af19528746197b428e81acdd71be6e284f0f5f1f0f759ad5f8c46c0deff9b0a4bcc16ca07e73b693cc9d4db3fb5cd8945db00131bf56b833c390fbeb15f0d2fdb30f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1710e16e7812185ceae974418afcc7786c25e1f4cee290b025a95d1724ad29e092265fd2f96afded966bc47d3b558215db5ced1e1f21842fc596c8f70c6f9f5a1a768;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4c904482fc4f8a04e0d7b3bdee08e3f9a25c5de7af961c24d77a4b782641645a8b8010f3bdf058558a54d937a318b832ea5ea00e163b7c6ca431c3735fd406f85cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c1e6188bec81da9496b393561e800b98ea5bf4be8f46a40b0d483cdb6c9fd9a130588f29622e470c1df00801b3e490f9857d6e92e69ebe4a457702d48ce9cdc0880;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c70f119889855f44a260cfd79e1539a68b256d89657a1036f1958ebd17854544aa0dfa57f69ab22e43bea80cb56e77e71a144a22f04e2bed804f7ca3f076fd71b29;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1de7b85dba794b0fa4044d6c99fe1ef38f01a090c39a13353e68b685ac23aa6ce54632af7878a8f66b1a6f606403db12634728205280cd20181aa41b637709a0d23ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a5d194139c90229729f7a5464c02f57a1af8bd15b37ea94781f57e252b96fe9ef59bb605ac55601fc0709458e740278daafb4f8e3b806c6760d8c9856ba042b67224;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3b19168e000ce800c7565e4d5e2ac720f77b7a17bdd472d534529f6a8a37b6979336842aaa6eddc7f05d8b91b5ac3d74884a6278b6732851d24282dc25c707125b98;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h33a0b0e2673026ff4bc6d9a075c34269fc6a07cd10acd4d7908c3b91aef09a7e3f2ee90ca0fd019c188ecb2697ae8785f9cdc5a388b84cb6f8644748cc31685c8883;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h707faaf683187f00d815d418f3bc85a139e1a1cb8fee3e1491b5d1c5e0ae58b846ec93541bcb623827e9c64d4583bd6d3779f4862f3a20ae70d5cd69d303f00e587b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f61dabfb0778a34653ed8c93b44650600879fc488e2e1ad1541d322e382fd53f8c51b754d50269520b16bf046cc100de298e78dade76f6693e79c46b78fdd7811272;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4011a45251a38989572a70c28fd9d0f78ee4e099e2176b07126f60acd520516f37cd8c456cbc4bca764b8846b06939f7c75fb0b9df7639b3ea3ab902a8681865825;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e690554a1d7c231b99ef716f53e84e637ca83b38228c8ef842986425b8be3036f092e72237ac0bbfcd59fe2c89b937422d9e857d080f732459fc4b9a1a505e990b6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h25666e99f5bfb67a257fb13828be378ec63938b24f232a7f646cdc5123d072a24d8cefe3e32e14963bc2c6af04e47de7da1addeb1795a28d6163462a8c26f45c12cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b6c6ca3e5c0f5b84f78f3ba27b55ccee7bab1a7dd082d0cec4ac19b662205bf01a4c579fdd998bd6c6823c4223f0179739d32af6f751f653ba3880f09d10f4372bda;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18065dc71fc09c444b7a4ef4b63dbb6685a93bf967d99079e29f087f63e4f4b9ae8e6c9f80707106846acffa8dc97e2a05467c6ab4c9e0bc404e54498c82a20203eb6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180c01fd06c6942a0150b870a4cca0118507c5dfd44e930fdc82ea3cbffea8c025c7031c48dd9ad0adb8ed5ac41d2ba06fd5dcb7860cd6e75bce7f69bc5d95ad72c21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16263d1483f47ecd3541e01c849089c1549e73b5551a69af5f2a837ecd652da80456866dcfed080de4146fa41863a9269109bfd265f73a945d3f4504cd15245bf2e1e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bdb8a3358f9c37512191ceec2c94e47b04b1ba53e90b36668cc069fb40ec11ab444a2a6e53d6f24203c0d5e2caceda243c2163f6dec1f9c2b3bd88d70840337ecda1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf81b40c1b6c0fe4e5a90f9548a694ad517927404df7fd7773a163ab0b387dc16d595a553aa20d1ce1e88eaa770fddee1b975870f87371760a8251a780477c850688;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ebda462d55639216323fd3c31a9710ad83e6e89e953750a3a976d0195b89fc9e5edd07cf6383c194881e853dcd6389f173d75da33be1534fc17a46b58c0b2400d1d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149f233ac9250b983b87c55ac101033128282245299a7ea2c2fc1cead924f7d1132f3d7c295cb34690216e3b61d4b5b62b5a23410fa148916e20b17bee38e564691d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha475ec6987a0395b8851b868e17a312ddad0b22bdac0eacecae35004d2a2b26e8ee0f074ce5452d7cc3f25e5ac4cd9528fbccef47121447302d4cae289b9b318b34e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h62a06a3859eea5266c4be190765838ac84f4d7f4469ad246bdeecc06fb2cfe1ad457712090dce2bbe3ebfcecc2e25bd5a0a92fb16b1b558b50f30337ad514adbf4e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149b44211a94021a59846258f5fa105d254541a5dc420fa5b1f2fd1a8e7c2d21ab5d2c8aec0fc0ca92758e872f62fee35112fb499de9c40b54b61efedf9ad3f17b579;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b2bb6be57e0bb153eaa6e06d0d9c29bac7130ad28aad63f67fa01c21ae44c2e9b3e9a7be1772c62e09d114f245e78bd0f59e36f7c4f695d8259d7949ea76190f233;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17faa44c6b9822afe8696492b29c6f8ecf24dc9d239d13e177a2f064c969123bb359dd50402f2640442dfde14aab730a353dc063c8d591df2f1684a2d067a0ba89736;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe82a27629a23ee155b1d4aee7801588fd6c6f7dad3ea9515bb4f35ce3473d11b8343808eb2b852a80ac83872672db634725121f665ac02e302da02b258d584c9b3d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f11ddbe501902843b00ef443d570b5688c434713c7eae436c0a01232e39656f4f5033b0de1060cf9637ea5574f58e9809609e8c864927f426f8e8c162356d0adf369;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0b603a7169d6385b8dd9fde0c8c5fe82c732b385abaccea9716ecf98a7fa7b6646b0b44ba7c7b6a65451e60c1ea027dd64b374711fb30859e88a13c862c4ed05455;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h58ccf862c8e4612112db238dff4e4a29fc3192deedc8ee9d6ae63e2f818c5d3db6fdd94fe9736ed47593c764cda82fc74ba45c71d6d1a026727d5852d7c366feb3b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38fc4f27d80be123cd12090854f812b3f63967ff67a90828f4ed75230a74870caf14897d6ac8276d9f810ae8ac61419f2696ab649a091f1ab84d4f48379575822e1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc1c81613ae7253219cdc56a79bd71124312c6467e801df0e37866b506f513034eef58b8c4d559f8b3f50a5d8b9f4898bf7532b0665253b3b8d5a8849f2c241b30578;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53253e6984aeda5012a9e565c7f6536fcd9a0351eee7b665d901e86085e71ef88439154251c57f3d9638f18136ae343f84ce9c0c0353ae320c18a50c58f5f409ac32;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dfeeeda86403e0c544df729305d15518e85839dfce808c92472a03f99f1e407cd83f5053701e08ff277a8fc7c7eb08bf869b7e71705b1dd3bcd93e574ae5eea05bf5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1941bf817855a2dd484950edaa9ca8b20a7a243de1824f5a2f62f19ad4156eeef5f3a9a20eec24cc97aeb1899b5c6b6991d522244dd690861adbd6a3c27a33eef6abe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17573dadfa11b01f4af2706e3ec215a872a61ea29f21d63d9e70ccb4ef8b345a891c5f3f5fe26d13307c9e659923e3e7410046863b3e29e024ea9f112f426eb70d6c2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a26e246849530d0fce3afb5b018c5310879f31f928aa66eacdb2899f67ad31a5f4112bc86e2ace0d257fb6fb05437aef81e46afd05db819f99dc9867ab4581159885;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14101e24f7d72ac92c0aac36c0112d4a4b3196209a9b6972c48761de51565b8cf7b5528e1aa4baf44640f703d955581c282039f86674c9712e5ecd2b100605dc63320;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbfb9576ae2493dd9904f53f4068603316cc5f99666bc280c7713fed7aacd5c773f8d1dfb72738d454e0f977f969524d7240f49150793dec984a6f3ad99496b9e883e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h63ce7193608db968a93bf13f302c0634976472960342c2b00444f7cceb7eff954ca66e36adc46ab065a6bf364f2b8f8a9d50414066434d8fc7095547022e6f360442;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd9a2d84bfac6eb80efc4f556a3a86dd423ef0bede11591af99031d3601c34c4907b95d44f818216c64a8d76d0f8f777adae97eb3a32fe56566bddbc9beb50c8fc687;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1200a0534bb507bcb18540a7f247a90bca88ac9926660eda4c4361ad919dc6803d3858fc150ed50632591997008295da89d9ef2d45525af98107cbbd119097fe45033;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf7fa501d5e2ab2ccd6f8780e36409575d257d89e0a713c9a884bb68697fee2bb597e0cd900e99dd73d4e84a35c4e238811214a5395067c12c2beb8479bdc41aa329e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a312e45281f9ea93564cb7e99f0b0c8397c9e37ab19b3381d3198faaf8e18f37189e67a1ff62be031d2772652bd8789ec6bed2ce8aafb93dd2f2c9a4b3b86162f94;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h127c25eac7cf736023ed70be89d5caaa474417b2a8e72191fda595f9198f04f793c713ab1dc2321d21858acac06ca8a8dcba366184751a0cfd653d7077f5517372cd5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e0fe35c9ac09dabc961ea97f898fc0fbde2df9b30c399372aef6eddb33055ad173c2c231c4e5d82d323019725fb0420959225f16aff3f63faf183d413624d0ae3d17;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd951e064145ba1af24cb3dfd3e4d614a0e0bb8939116b022e3678576f85692e83eabddc36e56d7f189d4a9dffc4c4f3c1523e0168b3cd0cb0cd643773fcd81fa6d00;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194976fa30d64e6c15b6bc150b96593fc34b97e1d1965d5450b4b96fd494f93c99dc8c958d2aca73e6d6b355696066deb2514a6374b9070e753f72e1dc523891e3a31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3b1c2b4f40503cc37517f90c05114b904a28538b32290e5903ca79208633e38ddc0fe26c03be5f084461187d61fe6502d8ba41d6417c0485245d228c44a4d8feb074;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120288478a90f27b15d503017db38b103c21ccdddbf1c33dfdd33e4da4f514e59a4ed20c23e2cb237db84f3df8327709d96fa07f3253684a28ed3cace0a24544dd57f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3bae02c1576ad29ac586ee30dcf0ff046b1ad0e9d5b7ff315f47b4c61d24f3550791d509996fe19602b8e11c8b30889bd0ed15798d7498b8c88db4d1f363aa31862d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h22289d535251c3bf11b9c5e0dd60080b10acca3a8e850f83af0ca15c8e54b5e0b4a81b27f6a17485dddf1b0d7d686f06b610d8ed8c15f846d27db8616e405d75e3c6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f4f90eef3c4c8ea2bc4f3e7224ea4e38d8d90ffac7e5a18202631fded945835224f73fe5942d5062f4a4c1dce65854c75ac4ad0594ed427b6842bc73a8f97cefde5c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1826f59283b9e867ac1a8e115dcb20315313922980a90e5dd596430c26a80a206bf4a5f1e424904cab6ffa99a02599aa376207539759c4a6dfe8e2787228464fdd3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f69b5e45ecbcaa12de25223937646df900a002f632f8978704eae89ffeb95ec9ec602f1eb7329903cdbdeb59b7994f9f5cb21418d7eb6a40a664a930ec6b00c5ec2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h563923131407f8e791ffe26346f083bce69445a059f9c8f9d5ff6ee12e51ab7937aefccb006c677aefeecff168f33ff4103835de636e19f15b5eba245f1c4b7d4e0f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd85a8d2a89082419f9ed0cd37f32535f85b5db2fef1da413f6331fb074dba209534b5c7880bfb3bb1bab79cb899c82316774f618f61642e353d80bac4a68fb4d6ba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fbe49f6bcdd25435046b3adfeb591b8f5326ca5fdccce67716271ccaa029ddcef6a0b566f2b75cda156b439da8c5b087e1c55cff7c7501a278e260fe8e1bd4792eeb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a5993b47db0b5904905823100a19a4fb1fbfe1e2d89de0e90a68f7136daae803a0f90fcf765640ef72e4410966281646fd8ae9ca88a7f422bf7518708901f11c3ee5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3f8b12ce4710fca00cea5675720bfe2893eb9a56ea3e4a1fb925290d032eeb930d97140a266bb80e5d9b3b5b83e53ac96d396dfbbaef7f5cdcd0737ad4e3fa719ae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haebee1d9d4fbe81ae02d257d60c5038e74539db5a7572954169e2388101838a7bac495fc78cb9e4029afc329a8a4c1dd13b8e82185bf58dcf16675bde868994daec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c8c45f2f5a50dd86d759e421ac4f15314f33c38eb43356f93c9c02d9b35516410f19a331364998e52e2cf33622ed2ecb3056f457efb39d06d625b190c495c5567c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a9b791027a69e01d63dfa3dd97cc77eba2185ab39f0b4ec0c000229a5ad9add70716043bf39897334021bb784204908c5cf70f5c85b5afc264a42950891f2f06b1b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17a8fd161b44aee972c44837a7f70de58cfbabc46a3f203594aab47d6e36bbd49bd98e5b22d75fba2fd6bf60e557811d0fac048e1a26ec1eae3b91462d3ee5eef072f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1267649af61da21a040a905c7bd16ef2e764fbc3099d3b46c4c15c1d1c5f2ba1cb6eecd370e5578196f432ba03a5df564cd3a011641f46a27987db40ea9d2e621b0de;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6956013358d626d5d34e13c0e894e8ba97139ec9b6b45642710cb3551467db5d22b82343b52736c53674050528dacfdefc8f03fd9e36cacd7f8653deddba8880022;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf9e5ec90a71a18b16aebd2029d866b35977b71de4163e7af03251d7c092b9108088396bebb1dfb0158b68bca6327b61e52d3ea170bb76fc0b6b9c2b354f690991e70;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h54b39ff2da22d1a3966e8b1e4b67630a0bde1dc8ab67c3f9b9071990afabfbeec737ccd1d4c548ac532bb08b78429da65eeca8efab7bb56dd49732cc26d60c5f7a9c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0f682433babe39766ba9a239849563ad9af428b7300219b50e8e57c3c08ef88ba36045b84772e4e2c60917f82bef2f6ad7283af7b82599b02711e8ec3cecc6f8cdb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67992575b41443f8006f6a0b74c53e8e94ec006cf8d0ae9030c598658fbe4821ec1f7fb4b22907ea4cdccf84ce5794bc635f041edf5696b6b31b665c39b0898cc9e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ce3b738f17bf1d551ec6a5547727ce95722ba2e327c7fa04c50ccb38a675078c69934c48271567362dcc59e14869a29ab942c8adb93027409532168412406d02e7a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcf59f059aad549ca065c739b3c2166ca1ad8e58b4f5986bca6239eeb5d6049f7cc1e7310dfaa31b4bc8fb6d4aa4608e059588ea271fac986d61fc2214074387a395f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbc6bbe765de14eff049b81b70c1bd2ca1f2e3e2c37802187a22f26f6d1acb36ab63c4a89982ad025ec4879c3f0d46b70ee9788a34ea3286fb47a85d30ecebb9ee789;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb4aea510798f08e1e5db35f245dc7b819d9004b70bccf82dac713f238a04ff7e53d72adbc62a362d6c29823f3e49acd2d1d2d22b44dc40c751a4054eedc17f227e12;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc2a157b48f4826256d78ca68ab3e730fac6b566463c27f97890e9157176ee6d8b3a61dd832fb67881b2904db852b40103840662ef1aaadd350954d0ad9bfb1b4dba0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c2dbddab25036abf9fbffa0a611543902b0e4385c4bdb9e81c3ec6ee4b44f8051df9141a85d03cbaad4726bb171a2111dab90064d13b38773404fdd1ce8717b4b92;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f6c888ce7f20e3837238f7e7edebddadc53e492c4705282e780d635d8df3a8662b739994c857f9f599c72668331701d1e4ab5802bc9820bfc7fa6e7a595086b3210;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a8f4d496e5d7067c270ad98430a3edd3139f79701363b4643a7a7d8cf56edd4dde67d75d019af625d57d59fc25857a1ed16637454a66d88e5445c385b0f43d81dfbd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae03980d1f74834d055a3a8a3373b324e1b431f9f4b92705708fc790693be1bf5bb7b21887d72313b85904836336d6963e5319f517c41994ba97f83ad215dd6847b5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d6ac2ff543d837b17148c56d86bc529dd883590aad725aeaa4402ebdd21a9ffaa86d09a53bcd82efca0f83135874971a852ee22f3b08fa52f9903778fe12ddcd6062;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd078fd3ea6b85a1832c98ebbc8331ed2f438c37c90600bd3778640ad6a6e3e67a6ba7d51869f9aa9804cd0e5599e54c3779f40a620061667bd3fd13ec4406b2ec555;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d1aaae8d586943e7f6710bc91e4c20035ce3e23bf8f1633d1a6c2af8f4e637efa5e35b7508bd4eefd5fd3760aef8f85f60d3d8e564a3467882a6297f0f2e134b3049;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he358e85757d4f1ce7bcb924ccf68262c59db44a06325e7a9adb81d659bd350faaaf6675224712047181f3bf51904194c38b8388cf1915c5cfac7c28d8fce64f673cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha013e0c3258f34ef0bdc4d4c5e254ddcd21fe3511d70606c322dd184b91411787933089541970baecfc6f772fe424cab0cfe963b5632c8e74f5198070edf444260d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he7bfce38f371ff4c8858d3c2a75d7529ffbdfc2dccb880ed2bdc3f0b050c90023f4d7f6e10493161a81e41425b6e20cfd11458d6835cc60bb64af0780e856ba11157;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1930b549ff21bfb78891f0b555a29d59e2357751f22b377b7568bafc1398422448a3d63420b61177469d23f70c74c643ce2998f96f47521ba6cc66b39bf43497680f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60dcb04a5d6c8ab2e8d61c8f662871050fce7cc69b845c499dd2e0837c234e540e59e69a2ea8e2ccf765a35e9bdd4e21d870dc1f758e548575251f6ccad824d095ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4d18e8d1b7872f59a80e7dca1e36d553bd10a2e4a5eb9e1086575ffc78a2609af0d385668540f8b6d15aeea797dad046815fcc5b1b9604eeeacea5259595f4be3ae0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2697d7d4532cc0fce7ff8e06c3a49068e816b4dffed95ef82fde8d3fb443a757d7ddab10ae7d36176b47c821e76a206da28cfea05261bea46e688ca7569625d94c3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a8b2882f81b94853f7b4c143be674e303a51efb6ccdd8d060d4f4c92f341b7668fdf41ce2708641a41291ca2a1ba3acaee31861cd523898bbc366196fd496450c1b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h145868efc092e93c6d73fe25fc082ce59ba7b32f38bab48848e1ba1b71c272332685cc7f405271e07a06717db40804b8250d90748f0209c13da7b09e70293f65d343e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd0f8c3aebf403da96e8c019966fb82889fa337a9f0dc8ce97a2a78ca3d0801d775317d29dae255c3bec3f9efbfe11c67aa5733e56cf2c6267894b69de211890332f3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37214068af2c0f27b76c623d59262e33498c906ca2cef2ea8481d5a3254d0851979992e1417d655a8321ab2832261e66a6679dbc1cf119b896b25ceb2ab35bcf23df;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f407a77477cf205d6bd78f2e615b1b44c3191cfa537c23c4e28734578e5cf5b1badc2f4f46c42d5ec363c300c744fd24df2dd2661ccdf8077ac0c01058b4e488f65;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca3a421d265cec4ca079c52529ca9f1b60557b236089af29b88af43eef9b0e1e8866e1e010a11acf72a124ff495316b3c8e02ad56becc7c7240b8ea07cd54a3d5b49;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7fac6b5ecb00d710ab3a8b2d8a56d223c4d7c44a2f1e88cac4ffd771ea7c3c971e9bc4212aa35a9aa3354f8ada55eb07d097b0773928ebaa5f7e3a61444b12cef496;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12df5bc814ca17b5b25f4a2433be084a87b5f6472c65561fc8e88d0977e8c62f38bb4370d7dde12b92ae859af5840e4960f825865c990606489bc5b83c3d0027da1a0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hedb9b524e42588682d2c4a6b94d7b80834e08a2fb423523eabdb80332b1a7b11aef96320e8de75691aaca9345901afc8db2ca05c0d5a3ccbed1fe4aa888a0327e1fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187c66c7c82db11edcd401c7ab165a62e0f6002ace33e90fd744dfc4f79a01fcc6a24f5fd63b8c4ae284f15006d2614bfd0369caf41be7e7893afd895b0baf09df827;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91f7c8674296a92b30f9ec063e738a5e22c3f067b7514056efda4ce6e44fc0b3f8653bcdcafaa6580bcbcbe4e11398211c15f36cdd4961e55527281cbe2434dac1c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c5da6e5c8e8a54a8635078c3c0e4f53f06ff5c04ffba02272bd4c262a058ff852d3114ce7f342f30e456dfd43ac6836248c20acc319c4d5d15331d68e7f98d41767;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc28ebbd767bff0eb6dcff44816d625a640f70119f2db56f6bc604ba732a40697994398e8a60a7b069656268d999e06fbe27e5ee4e212f75c9b692356d9f6d0ec437;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd30eb602283dfb550bffb105f2dade8afda0b4fb478bff7ddb134b7fbfbc90e8e1c93bb325a1b59831127d63e777d7c961b58c6abad303d1e006085144a7d6202ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f55d054d4af566fbea7120c96cf5ee02495c57d292da4f710cf441da347f6ba98e5c2626141467867e53c4ea0bd46a619f36810d5e4dd5bc1425d758b48827e281e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h178aaff17a09b64443184f882bf9edd3906168f530912c2944877594705eb579bb360cc08d50977a6f0221baca702596b6018219288023dbd94f4ff1d51d1b20d304d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h235b079fc0738a7edf8d6161075139a79d56c765dd2691eec4e257f76260c15ab400998aacfebfba76588662648916cb53966cb3a4194ce7a8e9513be9eabdd66acd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d39696efb0c447545b66774e909946a324fbb2b010d5957ef080af7294951f0178d44ad5cf9245784ec7dc5f1a3091e730b6cd35a5b019f88f7832d59bdc5834bec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h29854e6320ecd4ccc4206b5eb6c8a46bcfdd5281fdd106f9c27034c15872f3d4ed282b1de611e5dd7345c4a6951274a9f42a6bd1e7f022f2e8cf618c5211e5d41fee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e6ea20ae067acc48f2c881cbddc89c883fd072dd6eb941d13c6194f4f7fee9f04ff6ec196c6b7a5155176d6695fafc30c47dc32a158c52961128bd43bab5c4010a0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1342898c14bb2c096b8dc1620ad62a765da607bdadc72d558361569021c23264da770ea9126153b602d83f7a4c9688798c25c326b59bc84e9b57fe9e7cf5e1f36c9c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e4eb5654dec99ffaab8beb826430684b9ece98d2d3c684521ff991f1b66facae39b953a4c2258a15f53c796b1e32549c8a15e2bd5f352e810e14978c7018d0d668d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb949be68af6d20463fa79b7ae1040868611d288ae95012293a152f01b7770f19292317a3b80597ced98245af1bd72c05eff5e1e5e2bfe910b9ae46830f1fe2d5294;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f68131c1ad1be5ecbbca742e681e21104d4fb0b814267c75c198b1fd82218a93091537d991149814c0670198ed92bd1bae9a434610961566de4a8036688d30dcca5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15511b29b3766a92d56d7a45a3797f23949c916f64a9b4c211c3adb93143bbca3ee7a7ce0f7202c6bff60755e82daca445fef6029b4c8c0a1e088e521ba64ce3a90ad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h945d82de9a8b9364e08700f3ce6685e377494a460d8f45f0d4571b99fd977c60312fcb72bcc7d20ca44759889171fed6c51e0604e8c1f29be5631362197d4a92f03d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffb19b63610968fc646600b938233aa0e202ffed269f913f4fbea2c96cf8e25344c739808fd3e50279152f30ccfa7bb73ce3af6969a4ec26eddd04fc77dc69f433d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a40c67500b429569c6a9e51422840915da5bfc85abcd8abd9ec295db78eb392f2ba976322991c40fceb8bf42252df1f71dad239f574ca6de5719ab98726f88698b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18683c504ac530eccc451bdc035845e44577784b716212ecbafd475f6a47e46f5807a1f7bd99e088579f4ef6a185af511097a66c6a285292803fc00ee80ee22c63010;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1082c1e913eb7bca80235254ade811e52be779d478c2ba2313fecda16406192a1be4e37158fef17499f647f1e0892c3e440db3b3d1dcca02a0ea28652efeb23c8f6aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha056f0e886e12f7d4828fc7512ebffba5935ac028d94704536c395d00afc5ed1e65bef031ffb61a181474eeddc8b50fb156dcaaf7b6869f4f29d6c1f0586a693a9be;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h122b2caced36dc37cc5badcd3679e41691cf843ddcce0fddb81ea73b72aad0159fbfb8762e1421cff8fd7a8ae3623e09faf4f048128cab1221c8f27ccf37050c412c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h195f7ffaffcdaedbabc83446c4a1e45068d780b81bda873d864872dd8febb873d17b27c38846c91a1029b2c2fbee148e678eb9b2af0b16edc1b3d3bc4b7ccd69f7693;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e0e97b8c11f46d61ecf6c6af452ffdf2ea9c6372c1db4d4b2220bcc73bcb12c4922787e7ee3f77c7cb065a5d569e63592116a7095aa015da4740036acbd79f5ea1f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h888f21398e2bb9523bb79937bbbf15521443ae1ec13e549b8db0c2cca3b5693229cba6bf02a7dbaf03733eb099942587e71fffbfeaf66d2ed90228f35b4b6c1d26bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fa2a15e9d068ab14a085260ff13dc2011b3d99fa600936fc755fe2742719d872fc343ff7e769db0f8da514a5fda0f1b35327102999f5fc4d9e95ecce2c3029b3d8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ec7fb52cbe3b116699b9a233d3e7b8d54de81e7c4893460bd32db90331a1bfa662b95b55968aa45bf2f1dfcf2f10d4065753e3156c7b85f3f235f7cd0d30858b60c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa321a018fc1635f771eaaf3a6dbac0029eaf4140600a906c0f400cd240bc2b026200e6d15dc6e2f0d447cbdaf2a7b286c5a032a31450f4371ef1796b32fcf24359d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ddf6b7ffce545775a5d87c2daacb93cdf927e71dd0bf4669f4683019ffb0ecd39964bb0e1e03cfa3eae81dc421d19f27ec88b3db8260c14931d2620fd929779f26f2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1587be58a20211b0ea27921b71533342e7dcdf573428a41e097a3b8f981b2fab5dac09f37a7d9a3114d0a3818579c87c4b871e7c488b257d0d083bdd637522d5c0b4c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ad1e475df8e249dcb49ccfe70dcf3b54ee71065e72d3748bce39f400f29769f44a07b7c40a81bdf2565a5d0b79871976368a9862b3bc0894eeb3308744b5a12654a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15de6c5b173c6e2f39f831dfa8d07dfb73997690db07c798631b7ffd84fb5c8ace02c9f633f22345c359d76c7b823e4a1b51845b8857544cf63535c8ab0b1609e5eb5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc77353b4ad93137126a1ed8ef0bd0629cdce5ae0ac948f2ef042848446c0ef21888e63421fbcba06330e1886c967e976d1520a921abb0ee1b59d9224f8e9e6fea4c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90c8091f1df269c4d56037dd5fb1507e498decee9c277909869405412e9f001390b47d25f4b0167b7fd153ce3533e554833e47418f1689338b9ef442336e9db3d697;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c57678e84eccfa3af4135f4b2a209f3fc285188e957d370f3b1c3dbd5cc3cf7bb59caea12ff553cbe2a7b35614a7eba0abda2ce3fff1d9a53eb0bf492c0660277b1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfd7ca4423ff1bf9c87d879bf04cb2ed82e376d36cac2c467a29ebc7e24517b6c3b2c1a3ba14176aa30267bfd2dcbe2295f06ba1302635b274fb6d323b966a79829f3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17bf8dfdc9d6a51c545ba4f2097490c5f2dc1f260aba7332994b494db2abefef6445791063324a727a35153f5c29fa4ead2ea370f9f607a915e334df0969ab4947663;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b82cee5b4f7374255f1cec710989472838de45e32728e95db41dbcd48dff24dd42d2874ed6ce5eba60867b2a6e413fedbce5b2792e67fcc114118935278f0a8a2cc3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5a4df275f575d1e1736c3e0a30f52bbad33811fc2dd0e75f2ddc93bc6c1812dd530c93d2624fe4336d6ff1dbc2f6b5f83972a1b62928d2b0956a2aeca2cbcb8f847b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa1f0cf02e366e15c2e215cbef78ba40be36a4c9bb60035051bc61fb4e05428fd9716f6429c781dfb03a2904c0de83ebc388457b25c72408028e95a4f481c216f96;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he159eddae7e5d92b631f3845d78608bd78c55be5f7a615ef6a18542a5ad792ce6a8877561463073f0da266725d007ee3866f5e0bed097d3f7f5203617eca21b4c83b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c37676d09b6b8c4982d5d2558723e47fd2b6076fed734cd18bc238a464e10decf1f0342c375e5e12b9d23d815830b708ea39b3c0c9bbdc3fe64c85c8f698b29fc0d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd1a93f0919a0b6b7423c435360a99aa930230417fda1f33f89477bf2f751b409bcc7d8f28e49ee8cf4f04d0b4226973404b67317288590c6809358952e282b46da3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143567fb7c7223bba85fd4d2e3183cba55b93c595cef14b61adf3db7206680bc4fc85d3177762ee909fb9e1eed7e2009f3568ff9d92bbd06bcb3686f82490ccf199d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h953f94c52abc5b8958b5350d650074dcc6e9d8388c33af9cd8529d6a325b03ed208fe34c50cc29e99f99c80dafe4d7c1a8de9ebdb8f0e2015216c16a1983281717d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cde6ecf62c7ff3db335e60e0664846cf7eadc1328c829f10254b158b274053135aacb6e9afb5fbb39e148dd8b40d4f76ffdc9e7f4e9cbd815baccfdd1cfb885413d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a87c07615fdbec74b853def1a41f13123fe3b1d9681843c7169cfa0a5cd6c32a4bc1749a94317addc5c783ab3741ee2b1374bb5768ccd15c5c2e4e4e718e1853697;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf38a6bd773847598a411808a727c7e1f0db812eed479483d707f06fa3902d197e4313fc1e72c336feea0011eb74ed7ca79c57396baa99a1fcb1efc388597e7a19271;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h856628d8c1259bda938bfa02167c2e4f13fc422a815163b5e99bbe8128b8698f9d6b0018202fcbca315f212abf3072158291b61ada88037f5f85c8e73daaca82ada3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc8dd0833e701cd29cc4fc2c236d3f608d3207314eaba8fca7dac94c8fcc6c3e892ea07aadbf8f9d87b7eab99a2b22e7a15d9cbf3f731e62b9eb2f606e39d001431e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6aa7772cbe9bd3786401bcec019fc094a0d1b87f53a622b91af415825c9b105e6d2e101bb7990d65b03deb63e111af96b58a0256ebf7aa5eb60cb0c8ca935fb5ecf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h192a01d0d640b9db900fc2690a7318d792e14bd20ca51392e7b83dcc18aa3492601cb553cf64986d0212eceb027721f0dc00429b0f4a125b37bf50bc5b2a88a7cc7f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9528e8464ca300059a94ea8e6a9f7f9623399c6171f8c6afccfb838a4bd78b2be40a4a16bacaaa28e73839117864ceb924d2e0bc66a4891977e632fbd7fe0d7612be;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha07e289ba00987748ecacdb991c8173bcf751b026290dd537d7f336921f3ab59dbc35024bf5b01e5494c8fbc8c9953c1a1d97cd9b83a2d088bf2a37cb3e53919a519;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h950d61ec9bc742ee4f00b4b5eef720a08f0deb9996b700d3ff7be33a8171df31942e1de57cf5a91c13221dae9be7b3d38ae48bdf26cf6a31fa096a5d6cf18fc7631b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120c9d56a963566d96595c5a524060322e01739e059201e5b50bcbf00da374b7df7476d076b8c6d6f00af29098ec0ed4e48d40116d266f5cf795689f311219843da20;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b1e141ac26f887ddb5fb8a5b0f56ecc130ab74676c89292344f664fa024354f0c79aaf0fbd2863d2c3b6dbbf0c3c26c4f8ac75a97b7ee1f6d4ba020eb779422f4997;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h248a6e85da01a1b56f270b0a603635af26980b3cee79cd711ad14b17d3217cbd0b55be89731c288e30c3451a86a73b882dcbe349c94900df787938ff1c0bb1b5b8c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f079e0afe98ac86da48e8b249066c4a2137fc5ea5254c77b8eda6d119a3110f70a64c86574c93e8e14637df56bc3bf7f2336a049a55deb83e53727bb58d966458fba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba2a1ade4d0c17393f7481e202fea559a682a12e488150b06957dd1787b09ccf4b001f4cf1eac183240d61e484608def542fec3d929fa7f7801538f48e0a66596efa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a4a4316fb2d38da241d4edbf3bf18cdfaeb1168811ef2b56cb78d0b935bfcfef865059611daef530b873970c077253fe348e8731be3f46a25b08b458b2e30574d25c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1911f758c3df742719bb2c1680bd1e5fabb929601cca7090eff950f9179fdab240d07f5eb384c99c0e7d62c00ab454bc47fd57315dde8952d23aabbc0af9b183dd1dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h130dfd8586d57fc730fe7e9cc327d382616c21f51a8bc93ed1ca8642da1a1d94078d6658683379f7f5e1a6ed4d7e0b54eb4d77edbe7ea84833c6e45632a6fa5953a42;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb25cf8dc1ec941b4dce78082aa98e228df003cb268444e69c62a2b3043e174bc2d6d9749618a58cb19b50730be5e401c58711869fa9273d43abb2fe7da61280412ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1feb85f3cc78d8d9cdab5add6ff4527b97b09e88d54ecc6d7fef6addef2027cf4463a3247ea88dfae9e3ac913a8d3ff2114a22255bc1f782fe9dfa8e860a6eb99ab5c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19e87b2922ac6f4de8901f602eb9bfe9564c96bc660ace607510a535d1a060c1f4ce07e47ee77292d2cc0a3412a4d04adec36bb1bafc717aef992dc539c3eaa27ab4e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16fefc964940c627980951feabef309c0d82e991fcde880961e51ecc9f350ef7d97b920cb96a15bd5a53fd8353fc69e74c2a6b648d1c76348f20e06d4e76485c10526;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbfeba07a3bfe5a7223d9e56cdf3779cd6e9a499ff4b12397105b984d1a6bc08854365437ff184ab3a16226db2f8941676d13b18718c8c3adb901df9a5c4750d2db75;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c0b9a54d2f71f23f524fd1ab91f0a91fe8d6538b751ed323acfcb37e7282145859adf295935a7a15f84741733939c7a3df45b07eb82dbb0d10f388d41136f8ff278;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fafc46e1742eba0f6f21bdce2dff7a9bc8d814ed45382b110720e00f6ec0f6336dc540016967b69da851e4abb2d9845d303f734b5afe24b8ede70495f1cd335badb7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13b667360fba4436b6e297c0e09178f80f8faede6010d1c3c2bd4ac5b402c6c72a2595c79c490677ec4b69dafbdde4f5f7c18bdb4bb68a4f8d79cf4081e9c3d8f57ba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c85b3b5200b83319387be507a88940bfcc213b0c0fb10bd269c35d64d76259fd49d1026c0c6ba4b63b4bce44ecfe7165345b8c7322c626ac1375a1324aa3c2f42c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79c9ea49e8ca0095f7d13f813bd783a601dfc8eb0b2032d7e339ab1892f23c200165c816162e152158eb9b7a05d3cee72a69ff3f90f6b93a4c4c70b798986d24a73c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bed14e31b71d84e7b04d8420c5bedb496407b2582d0f62a6d8a8e176e8b0217069349d1186d70b42f55ec017c3a188a08ed6841af877c6932a37be7a07d77b52ac58;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2f57ed7b7845eaad44976b5acb4f39f0dcfe9c3f650d3bae31036c163bbe527c50b5ab94b21c9049c77df419a46a715a355c22a2db60c39a47fe8fb90a063a5151b0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e4a618ee21181dd60619c57858d013b83ed0746dbab02976ab7fd9f2c8ea4870d8a02c38e293072c9fbd300be6828628cb39cc21f00b07a17268450eb1e00331e9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a490ddf86d9e1dc693ebb7a344ab1dc00b3bd78020d4e4dd5d0553585dcc30ca1b78efeab78987c87aac508c2a9bdf31d8633fe3eb7ce14b32c50ab4cef2b1315c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hefc94ab8112d917b1b9c8605c7615e3d2b6bed6df0b543935fe343679488678fed23326ca59331e1e8987244762145a247cb1df032489ec9c61dfe4be73289875ca1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198802c234e2b6dfbadfede9810a678e9d797212d76195e4137df8159522a7ce7c4d58c8223520b3b441de2b916e6cd2fe4413f747b019a4f0ef8f52ca675132a58ec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h114e34d06a5224f38646369f07edc012159bd488016ff83af481c2abedc12eacec2d71d4f6f285a9d2596f30ec97ea309f4b0e2786f469cbc737e5364b689592f61a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38012e87a4de944418e64aa7280aa9d2e58f9dd29ef0c86fde73a95cb4bbf2c41f1afceba89001286af61d534ab954c0408abf45744824eeda94d2a055d9e6bbacca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h892dc1cef35144b104359bc6beb5cd93cac097814814bfddba719d137c2584d807da681c3668033796058b7d7077f83d6ca79ba92d7c97f2de7ef5e6fee286aee082;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9917c83f87582741f85b4ba10647002aecaa7a4cdd46eb4e9f5e81e3be639c1537047f516005ed90a7172dd5d6ecdde800c8bd52625917fa52eeeeeedeaad4d92114;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hefc11c9cf265b5329dc3c5297a00a9c3f729c33f6571cf60ae88c7d73389ea9fdfd1f89a43da04c8ced785a7889be0b19524094025a47c54b741caa03912b6240a20;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b830d773a3398065ea1851ff3ab09c3aa6bf62764587cfb00db085f1245085ef62f23d342b0cc36b1981cb32048bbed0977b8fbc74682fe5d73861e3dd8b7e46f3e9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h81d17b9f6e922ae794cb260a672f14507255aed8b01964cf2473b66a74b1a671cf87785889b8af99cd59cf035ea35e077fc705ec6af7056485e0b039b20964586799;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca082f3d56ebbd27930b7dde17d210a83596505fb909b0596c0ef1abf79459e65ee2a855837fbe8efade96a8cf722053ee3d79226d0d9d9977a2193e8fdeb4ddfd63;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h167e3aeab601a026112b9550908dbab0bdaf778734cede4da94f344ae10769eec1fa89c78b40391c632fe9d61ff505a0ce44bd13d9d52fc8a125c358333bfbcc03c66;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h191fffcf62801d9fcad0e7f3c47a5e40866700ed5892becd539af6259a0d94f3f612efd7d12ce1fcdfa41f6648997cbef84bb3d1a1fc045c4bc4fcadaceac99e85ca5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17519d5fd3dc49e4a29c887cfe1c19ffd0bfdb06d998474e26dae5f63bc99271c93c8473ef07ed23d24295edac2574bae7a306a11aacabe28f6bd2901a4bebbc9945f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha7b1405647e2529c688176f3a2f9760062866e7795c2cc3aa4abaaeac1acf80844e2669c8c58cec10c2076c78bd7be46f612a727c779bd532d0d0f4cbacecd0b3848;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fa9e83f75049162d0019a03bf1480f95c703a196341eabbb62974cca4730d8aae52b593607e64131bb3590a9a16a9dc726daf480a074200688f9d27060be85bf41d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h51cf6c610f98835580fff646e8fa6808d290bb08ecb1244351bbd99a463959cafd1421580e77cd4b2e991018efbc8354a155923ed20a2cf53d153f11468d83b42990;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d14d322a1a05eba8236b8df7d6a5dd5b6b73330af1d40165f53e0749666cc816f81a012e92b08171870cd2ed59bf34f396a9e524802f6c87672514083e2af962a73a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h168e64be4cb39051a042f96ebbde50fe413930989f6af18d060a9661a3099611119f7170a1b80b1c9a2a2d2747497ee1838603a1642fd0494f8da88c5e4908e2c983;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd5d4f9d425cef9b993c0693422de5e6189f88ababb0bf3756879ea266b0e9214b393744fff3024c5d49c2c9abfbdbea1a25bb866ca505dd915c60917e6f4f283a421;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2de4f1a9712cb7bcdd10ce8fbf780cfce5ebe16d23ab4baf34209f95d739d701868e55ec23747bf5e44265110a9def8c92bfa16457743aa88f27157835e5390c0c75;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d124f6290add09a580e6b1959922510f82b71465bc20133096c0fd243c9e4507daad5c16669d284192f64cf538f91801799c0a8a26d69dfe6d1b30f0d3904dc4c61;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h134e0a2dec9368e9067b70e4448a46b668b6ba9fee62af25665242c40579797f4e901b7bbc405b6509d2f7006d71cc97b06e62eab5a6c3159f0c6383518734f0731a6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b456bdf9d080846087eaf627cdb0e3c099d9d96f7329d46601eb0c6d13700317a44bd732973db3f854e63b47190e9671dbffa9112667531aef106ffae3b1b7c46a1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1263d7942ab311599904f32f2ac0eddebf5727730efb914728dc6cbf0a296d13f756688791e1672abd618f9fc80b881b2653ee42ce05f24390c10a536e179074fd503;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d61fa726187ec41f37f57f9d59443bacdd6966b7b5c7bf958a009915ea1a9b9444e78e4dbc0ffdd9530b9414d992dfe5e721c576ec41269dae4e3d349dc60c543e10;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1989782d88a1891ca55899d1a699c7901b36843659e0d99d73780ad9b0ae2c774e8289825ed77e552ce52c28c0615e8cdc8038688d5f5d41c56de02587dcca83baf2a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h197e9546a9381d7c1934b266093091dddead9e6b878210a52c3d8bc8e56515217729d1484c807123999d35dc0b8416dfcd608f44b6a8526419c21687790366d6368da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h98ec6629a288a778c26124ae5c76caed5c5a9c519bc5d863faead830f52d2512b7161be2f8df39b06bb80dc26be815b284d2374b91998d0c51a2c2cf2c363ee07e38;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h154dd93fe7489f2c86db7c46ac525d3948485d6c6e6ae463c77e078de5b388d9759b716f16048c155760474aa1e267a5b4e18db45f245469436f3c85bd8944ef9eaf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f3c98409ef75821c7c2b73a0c019df02def35aca12096f8e973c5654b7f69b3fda81363b747798361faf48a4debfb43bbbdb4cc1757d0446662c1372d602957f483;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had44dc796f88c4a9daacce81c3e1661fc3cd0503304804e84119203044f7a699cb0a2ad091a715d8b8ce496f7cf2e14b9ff91fd59e7ce50e56204b63e79455d46b9b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1774e54efd9f7df89ded817c1a68161e51abf174322b51e06980ca7fa046473a36a23d756faf2aa0d5800d5dd6906a22e175897e8541bb239edcd5ed9a024ad40ee97;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1524f3ce8e0c59ca73e4a3963f4b7107c4ddd41df8ce28eaea79cc4acb1ca69acddbb7e50527e921417d3f9179bfa35b908862b0872265584cf3f85869972aeb338c2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11dbacfec122a5ffa5c1b6b61a75a8ed77c5b817e4eeb7abd3d6623a09973bd22e49d637b7f8ad96d438bc848f413a2e7729c0614ed123ff4262d1e7429678fcbb93a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3d041114f60a85626fa7ba42ba7c1d284bec9d50cfdfd3d9485d31092d2c39ccc0fa1420361f1b4bdf8b98289c9be82522cca722c26c109040e42917b9918ba39b35;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h54eb2ec768cc5fb24b27393a6b36c7903376ed1a7ed9a548ecc6cc7e87f7a814b74c8ecca7d738d1f05fa06b816060831d3ca5b523909a2374490c71ae44a99c262e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17baefb296ffcdf8a178a75bde88e90f26b23d5bc4375b03da2cc9f11a4d6b89924b8dcf57e3f266a0267b654333999089070dd488cba2ab499e2e5c248880c67a2f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9a1f0ea47d2d1105970a6eeda714e1e05dc353423ba8d2c48ce5880c7431028d666dd861aeacca782ffb8abafc5a10f8fecc72e5698ea1c3941f5bc597b8242cd4e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h303e16caaecdff351e9867fd0fb5b44937f11829b5eba023a400f95cf1e0b23468985dd83859a6181842eadf16f3298e79d5e96a4ebcc7f4f41203b7f5d4d161c36c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1225ba9e041d7ebc33e5707bc39a13537abd3bb6481caf763a12b891973234057e7daece62e812f62ec938af0775bdabfd1721f41cfac779b49be38e08634a8f28a14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14be337d64da0ce6ff098e35dc7de73aa03bcb24d8f3b9ac8b88905bac1d4e3ad8ee4dfb5b46b5872fce1f98d5ddd0ae7635c7fdc6e7922f648f46e7ebce8c0ca4092;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6cc8f294e8017c7b54d197220c8934c5f072a250d9faad6dedc28c58c543f93acf9c07731cbedd030dc7dcfa6e859f418624ebb75db8d061dcef12b019d525d27ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14383f6bd7a08535fd52d3eb3d5cd6d3745258e239e5d6cc9669070d3840d46104991de47d3c120a64e7e1f6c4281431b06669564ded609d52195db86801d7e7b4cfb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2bc749e33f7b6ec68238cc84a742a6a2e719f21dfe53c6de51ea885c698d380c9d29d5903d8c0e962565552b66d3f1d6c4445cbc389c72339d0b4a7c382bf77f770;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d52b9c89224e53ed9203dc4b473e8224caaaf83de8b0252159e6ceed4e375004abc7e91a20b166b71b01a3fb87a1dc9a7f0a64ea721087464a60ab0bc048a4a9d5c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h132cbfcefad95c1f0ec74bfbf941e706a89d1c0d4c65951b509e5da31bee4be123eb216ab4396f156584c38934d2c6bffa825dfc4a15d0a1c8d3e8ba15bdad4e36df0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f5afb4c4a923a514eb33eb6357b2310ded6d42406efc50d3aa64e8b3b4e614ec9348e6cffc33431c172c247df3703289d9183eaabe66f2cdfde91e957879ca85fe6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ae664affdcc620ca5407e11be31cd1ef32347365a34cbbf7b5cf30bf7f8e4ddb3e6b95aa2fe57d41df1375ae2b102bf7ba9daa5f8934b99dbd8c86e85c3e271a1f54;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h189cd5e25062450c9630d7780c2771c8d8f2e3ddfea24b772a7584e8b9a1f30f4f6a7e33e412921049807ecc608e01ac751570baf9962cff74681940e1ba7cd71b09a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha5fbbc5a69b6a408828a6156738ffa7747654e17408811aada15e3ffbdfd5e6ffb46c1e45c8319ecd4edaf0d89cf6900be2269f64f77fb063079149780c801e5cd85;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a6804d38fc8fbd7cdc03da2c6a05b56d996fb3184436b9fbbc2651047bccb105939a6999b6b47e07362c231c1f9ff71df36133ecf039835dddb0a69a16c942985789;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e4e36c932c6f2c66b1eae95601a0b89b51d7d13dc8eb5c2b97068069eed91dbf03ced1f0935e4e3dc0970d55bc665199ffd987b0465409cdff7eca05a242d7bd258;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b381f23e7916cfee348cc2216aabca9450223693cbdc72b7a3fe515f4bd42f48eaef9171a83580aad7ddd954cb57f5701416ce3703f4852848a1e351da5a0ccfcb8e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h59c8601923ccf5c90cbdaf5de671a6c090503e676505837e32396b3fab4610a3b43c3b3b01139afae3d25f6309a6b60919041ea3d29a1176c4427c79ffc9be2dc8ba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1397e93a2f32f513cebfdacb424abd258bce651f6c0aaa1d73b55cb4415b92bc5fb0d59db4fa7f3c0be923963d1107d6967b6d90fa3416eefa7e5c93d9d02eef9c98e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fcf5452f71d726338ca5ad610ecce31948bd1659f7a4e798f96126b6651b86350f7c96468396c3af99d02c5bb712c1d7ba77a2aea06ba2eeaaece06a692b66f69301;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10fe3eb735ce3c43b78bfe34b0958b344a89865783eb6c1992e206667f0be1b2452449c88e66dd5023944649e2ef3dc3b7a4a25975876f4d7a6886ac1d7f6575218b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he1f19c58051e8ca2adc0e34eddfe0745d6994a765a8345354356f4a0eab299c2bf65f54aa0eb8aabd4042d80862b8e76baaa0b9ecb2af853f35da7b2d96f3ea977fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d93924420d00b83bc120e2d8ba32580c8700131fc518e3e4510959bed3d85006b46a3320804016a122f04791f2b8e3e4666c176a83c59fbc0de1295428d534962a98;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hda8b4567a9fed2565d72ef5292e3d56bf4c9ce449f3769922e1bc3679717522d98c5318ccae0b88ce2b6b4f3f28bb94f132bb966d9bef6491e72e1a2ea8001496bc7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f4067efcf669860e051c5a471db4d539f6a8643c6ab11e6cc1720c1d3416044b4f834ab3392d85f67719270b82ebc56964c405229cdab17b861954132e8995fcaed7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f2aac2ee61cade24fa727a09aea332013dd5e8df358de54504201ba8e40fe8f22c47dc82ccc78cee70a94e66c102ba9aa5f12e5417c715cc0a462b4acf6e34101e98;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc237d648a82587932fe109c6f1332cb988c9a673708e4c91b28e38896cf1b585334ba699ade7f368d41b825ef6c5a033fcd3057ccbf8debb316280509b0564f70e48;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19f09110fcc032a2f89ee3dd09db00773d0e1967cb61d6a230b32cca04d5140173772679b40110f37e4e7688e89976bad7b7c01f8aa024548d396a6ccea0f43a387a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h142983f16da3bda5b68018e5070babb7f6d47f8f15e5aae71ca1e21a1d239ffe1599cf9ef305f6363abda60ca0b7ed42e884f39cc463e0c7465873ad19ba2700c33c1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6c325cf34de55c99b22f0c154811f712d28de6cd4386323f736bc47c39797e5a55fc9249559bf4ce2c71f1ef72aa370a01e6012b8931a0d4969b37db0e99be8e90;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180e32bedac4a3e9cabb7888857b610775f207aca73cfddabecd8925faf644eb723a799f3dc71d641b5bf57b2f98b44701cf70bc540a9bd9ebc905004ff2eefefd4d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha78104f3db0fbb99c3a9ab7afc4a871467a023b0edf6b8abb4b7396b0b4d27100f8d103344fd0645a649cb33e3a5f95ca66fed861a4ac18a8779a6b1aa5eca7ae8f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e867ddeb68864803b52c9908c84acace1dc9509f1ba38310a7d156496fe9e065bd564f74ed467da20b9a31776e96e7a222021b990198bbfad5f37c21dadfc8c4364;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fbc90a3715e857350ed054202090a48cc541934cd4e3494fce894386e1bc92f1d890fc713f069c3e0695ae964b02601005dd5cad0bd0d776a393a379cca2403f8696;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hda7661e26971ffdf9db8b84f437b0a3300aec329e3e7b8ed06fab72608e52e2bda35671abec54b45bf6b32658f2bc9ca160496373e461886e88c00623fc809e30f19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89a0e04f08d5d6c654884b4ebad478e1407738100f906280326327a32290c708d53593d8b6fae14e58204759b6230d81153ffcfba9102fbdbed9c3dc331e0501e099;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h183b8e293332fb1f3f78a618e9f121b978116a774f0ccf0a977e929347e9b250de5bad88219bdfd269a24306d6de035b7af47c73df80c4d47903f72c11563e3178cec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dfd6f48ff7c51d37ae2f2ac1c49603487724b3064af46f80a4ab87b92331e65bc497a6abb64b9b3ef92b8463ddc0cde2a1b2a3e4652ce636ad3a84646642a6b301c6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28ea0764c2419769d38f406f8c5d607f87b6a2c856cfdb97782261cf6d61aea5b8776eb051ebb069a1e4970da60fb7e5afbdd94a6ec053fe9e4363e159011546ce99;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e02136440a8480c0b63b0867a6a7b71e7309bb8006f44587015cdd833bd8483939976711e571ae9892a033d59ed3fa2790e0c8903e4f98b558bb656b334996d6e36;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd158dae372c60f30ba8322956003c477542ef50763f825cc7d10934709d0639d107e54effb246978cf7186fbafac2a6f83443b80adecb95871d1d84c31d9f0c60b8d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1197cb87dff213ee03ee88d06c7ef564cc0a880b9dfffbb34d270726f645f59848966cc1148f16650489f107c5e738d9e22370b892531489d9bf8597a51d77d7c9bfc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d004a25812311c0fd5c06156f1c9e9f24b062605d9a81af35ce7fde600c389f1b03651df93c90cf450a5b0f5fca923bc1fddda4bb0e9a8a858bd03c30cea6f476827;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdae4b0310e506449cf71ec5620e16374364c7397c1dbbe39b5cd536330988ef314c4f578a8d0a4927f08d5fa325b69216104d908af1bb07baaa0a5142c9de9e8172d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h21f05f8d7eb852caae8f89e3bf1063b18dc09988e85e1a926d3c22102adcf608fe6a9d1c759367ca097cd8cb61ac8c43bc7753f8cb3ff3bbd172c9328f6a66e01af5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h234410daf591ea2cee9545eccae0aaedc5ea4d2eba1b066f32b9db3fe8c26ce856cdc21bd7991c5db98886c651659a26cc9a86d396c206204b65bb6cdfbb5509b35d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4b9fd5757024e5c1b007ecd6cee19641a7b0c2a70ae2caeef68a5e93db96aa45b6b7a93c34b7377765c8c7d3f1a85cfa6e5328a410ad5a42671f12f4480ce775c621;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7d5e661e0efc143d9d44b23f7d871b43e4d95f6c21518def2338146c82656acc1c132541bd34f9c7344e33cbd0e7d4feb7adea4a9ce6fcab049d17a5a8d135337e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h162263fc4431ebb2ec027cfdd3274e064e59bc5cf28ad4b31b90d132a86affb610ce448bd6d8714dab754b5ee8818af165ea0f85224088bc74f885bdccb6926d39420;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc56ce3eee09e8da5c7b1efbfe6153ce0d80c5a179fd32f40dd277bcd53bb632daf5687fd98d3fa8bbc46b8829dfeaa1508b6e372887722f0b75b3e350a79f1a73377;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2120ab9b496cd1da3869f5286ad9aad9e9160cef1e3f19a5c4cf9efa4c61bdddf0bb0150432486e820bc36d4af51d12cca48c5d53dcc84a70da43906b0d441521800;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108cc5a00dccb449303e585f0b89247a81e40886435af9b84587320e303285da607d415caacf48a9bc3280ced1701de226aee4a578973f33cf991528fd3f3fcdc22c1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb547e40155d68fd5abbd0cb161c06df5335e4e760347acbd5982b6c58cc1afd626235a7f14917e28cdccbe33a322688953d9a766efe011dd66cee20f6c6dc565472e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4728fa42dd8a7a329362c36982ef657e4eb6b43f6aa14d0b6be9acd325cc42b08fbe631b1739e10da4bcfcaddf0b25cdb97971c55b0cfa7a59a6aa88f67390b91e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h22801f9e7bf4b7266053c44e7f0cbab189ae7d6dc1267d1bc0cfb610472fa171853d2b3966bcf79ccc61cfe9fc0adcead29eca072bd2bfc5bfdb8ba51bea3e3239c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h43fb7b55a2b0db778dbb67b862631d4941444dfef9a45b7c1d30303c7a91fb819202ab54e73116c9efc7233655ed654ef21bf036442bd963acab8396c8d213ca8173;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h176f9bdfd9782e5f6dafb8d996b619c463de8285223708637061bc91f331c5d0133f37faf3353424d074c1bb41190a3ff1b3402c1c94328e588b68616e6499e1a4c03;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190aad0071188dd49a783502ce8a653f74830173da7b766b45a272159a17ca83d4689d0a1de6d01aa2b951ee9dd968c5d1478f38d2e7d17d0f60a2eb7999a78274be9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h106fc939e8144dae717e475d3805757b4682700114826d1c75f8a4d480ebd72dba7cccbdecc0f530eb3eee0b90027821aaaa3493ad9ca4420917b630cb0f6c204a02f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15bce14794917eb7fd59fcbe3a7f519bc656cc8abe26b3b980476a78145212a6726f13db9130a3087d4aad9921cf1a96d322dd607c881f55460cd586ff8f7c9293180;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3b22cf6c4b84faf5532746283b26290cc42723d88c57b85383dc7b20f43360b070e84db10dadd275d533b862078e520bfa7ab099e1760f78d3fc9929391fe3a65f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9cde138c8f720cd5697a9cbc1033a312933235da7fff7af46503de6092d5e98d008de54f5cf1594f08405d412fd0a53c390e721643e325bb8fd48b3a9c6a4250010;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h420a13dfc66464a0cf15aa9a542a175d102eff1961242436c642652fa2866f537dca0659e561fa9c830411f738f162617016b7e16bf645b208bb8b8249c54b17d890;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h184e6cac9f7b424a05218e7e072ec754e602b5e894cf7e3871400768bf3d124cb34134939b54b765553de1f5245aff12ad12e12f6a5a952abc485e1a84ab4f554d07;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce37861f99784250cb06361a78e98ad7f09a865aefb55e7129f908b1c583cacdceab4c4325f919ad2c795b95326d2d774b34e78306eead777fed7bf7f4ff00e8a843;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5bb57123fba53bb22f7dfbfc05dab37d94d76162d242d29e29b12f638a93eded5cf58b3489324189597da74cf8264dfcb6f4dfdc257f16800f0a24500f9d3d3d218;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1748b3c73638a82e028f3982a8bb2cf9fec6a3910bfe831ba53b4371420ec4fccae7b54ae925444c09fd8aa395bf793f0cce8da4d782e15bb0c3e5732d8e10e48be0e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149f9bb68ab3dc00cf90c8d5e04b1b5d672251952b53f1a74c978a0bb91baa47922b2b5ae49b75aa4ab20ffbf7ca09ca2371f9a744b5309902e5d0aba1831d2084f31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1096d9bb78cd87029af07f96c6ef8cefb9187e49146cc9ad6cf2bd37a2104f6ac903b63628fac5b3bf1049c0a9dc4ea688ebb732614be0bb82a7fa8722640ac244db5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5bf1db3980a58961febc53519fc7c924cdb78158e94d96361f6ff31c98dca25d5b0783aaf214c5ed6afe4197f52a5f9c7b90195bb62bbff92fda5a4d57e36976a32c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f13695d3c1788c97cf272336ae75c40f03e36ad93710eb2ddb5dd719f6757950770b19d3456978ae2e0a7ddc1e15295ac85727116d4da8c8b7e9d8c25e8759a6b0be;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1907063153ccc97c6757225be9d3a4e059f6fadce19ada42384a065954f78978f4a6786fadd9aee39ec8ce27e455c26dbd6bf9f2a91d837e838d9c5768c5530bbc686;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd895d0cdb8d052a90ff2e8837734f5f927c81e149baf6af25be8c19c433cd5763fe5b7b2accbe591e73a9388fbe354d45655189f0abba028ad74418212987d4fc5d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15765e259a23c09b5610b1faf772698cd34b93d2c75c24590682334e3927d6d3b6eb44673f05aaf6a97a3d767b1c83a02d0bec12418cbbd644dc6c970d546d8856d0b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1db4648e609d7d71e5f5174454ee28e5f29b61331e1b1e21b60be3bdc66c6ae16c241c16f25c28325640606b97b5d5b9ef1cfffa24a484a2516d5294a58b507507824;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11479fce27b16d7c011eba8ffe9a5a0e28dd8faa9fba7cebc2a16bc4ab966eee9878476b9dec77e18391331393fb2fec4a19f63fb1079f5281fb26e77a4c74d49e437;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150571af6e38985fe377bad1befffe35af6e347052d2e6c6c77d5d8e123231600e4f53e46ffa4c53bc65914a6f7dcd7904680315eb20dd9b72c02d9269f87ae42a4e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he8a5799554b70209a3a0d51ac50809b8424dae89683f19fdaf2862976e87bde86085be984904ae8bed1e0124776bfff37d5dba860979951c92961e688e516c191931;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf8ab725d4438530a341b474a701840e7ef3e3c2662f50475aeec56b103201868b26c771e1c2c958ecfeb0deb8cf0a99dad9017426cf021c67752d6bfc06203407bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13b08a830c67087cac33fb7df3f02d1a5cd04f4df5c437df474593bebc3736d4a0f65d5a0c04addc22b93068a8c7a9821d69126de35e61497f8e813e6459b1738d95;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118498ae1ae05ec1472bac64aad41f5c264ffb5adfc41481ceed5e44ca24a0132f276898fb83def8864eeeb8b528f5a37178f1d476156d8cb41b792fa5d6d67c8eab0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1531a423782792991733dac1ae44448739bc250280b8d244a8f2e75aae71851723610adb591261c897b3ed61077db8f19b030f2f3ae33ec75d885f1b3224013bb4d04;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h173e8ef8c7e0dea661df5382a9eb44e70e50d101a8aa0760090f16bc08dee8ab5663624dfc74393b1adf81b6d14f20185aabc65858b95003142a9704dd176f7a6b4b0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d04504ebd4705bb38b22e1bd8462a3b534d52ade03bb97f9e1f7f722dbd3443e06fa3637776979c7485fdba40bb44c7686aa49852c6ed22e1253d347b082045c5aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150817843b7d3a856a8b026f5dd213d33824dfd51e0205e7d95d5cb14de2508a9cd6283e0e19cd43981d763564cc8d4b76915e3e5394ca8d39c229a8a5450a6e2ef77;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186742f330b60220688e23bf3a2ff6f5fe074cbb52c33bfb3d27a8418ffce29ae0016f83a3c8a1cfdf5d5143165155ae3f02ce02815e75d0c2a217619beb5ef8e49f6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h65a82a3f99ac6fc453ccac386c079571056308f25350b40f09778119415ca715ddb144b0ce5c550c1c9e32b4cf371be49762b2f416f6cb941fdc1a54f54efd1c80f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17aa9805f215711f4036eaa4e7666d2e571574885dd94653a756f893472f63be77b47b2bb217d6415e8389eb9e820916a2f6c83112d6c517f04b81f9dd1c799802cf5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13942157a48cb8f8f58ac6622fc54ac1534433745b67db285e07a95fafcbf1f9af0d2b5e873d45abad5d1ae235fb7adfadc8510d25d0cda19d7f2b18406d4516c8238;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb2471f4f787c272ddf5dcbeb7d3249f967273dc84e3ff41df67205fb83e219e424963aa83392a3dec4a693d1d3d613df65a37c3453f48e1c4aafd4667128c713a347;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac6c2da007a8b5190cc1730dd8cde75f6c2a9e7eda4036c4d9f7d45385011149f15ccd2a825edfe5e084c1267ef7bd1756861bf6adf88eecf7f521b851a77477a92b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf155ad5378bdfea6ffc10cde0bde4b438a525a67875bd62400d5a4d6e08c72e8ef37075b790f979dd9a21d9685ee164d7bedeec96708b01b317ff7253170d6c1af8b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h250e651db330bebf656410df3d6616e43a4d67d3cf1b067e6ab654f2b5b70fbba533214b5ad04fc0ad26556365a58b42fed128ccfefe9d93f14696bf67a99b4e61e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15f69e3cb0002b18c22b82187c252414152d42bb7fce1d1d563c1493010b6721140a97372e9886203359424c2237e10a4383f904925c4c9e6357a05d8c0ca5a70dfe2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1373556c708f2b67d6b4ef93aee96b47230e43872b414be72aec32300cd733c689c1aa684982eb479c5c5c33eb9cdcfb09cb068cdd3170ff5a13a46e7f4c234024cd4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h741fcacc395655f1a94f5b4839b9dec82a422c7d7522b13cf908f1b5a02cbc13a6f260e1a7bf7383cbed2b13f2d66829fd0b875fda7b8cbb1e183ccae195a2ad62d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143448315c11c61904b984329ccdd9994fded03628726652a0f98b130f9cd7ed5d0038910bf498aa8b13f73c9625f1539f8e0b13ae81cdf5ece8327f30d19244d368a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17323a9ee6fe857a842556e33b831cbd25ef91d2ed5e3dbb88741e1525a8380edbbef2d2cb2721c89006d433b40cabb40b695d33d412bdb3ae33f83ff6ac96f1982a1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9cfccf69f4a72a1376e32fb3f04f349364d2364777aca93c90569c9384ccbdc9c3760383fe2ca9e52c743d6ddc593e2b2a7b863fcdf09edad8664d95cc5e6f2afa5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17bea72a21b97b3875c0b4d4b71b65d90924b89f7e494787674fce4df3a1ac63ee669e84f333616170c00b911aaa5145d6177a7cd5f44b0081519942a3ea728bd5c0d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h36cc61dbb732cc74e3a8191058d2fd9bbbccad60b73e21b8061714c75843434b7f5ddef8ce0e397c6c3dffd5f046942a3128fed752a3810abfc267847880f5a62d39;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2561b5b43a4ae66e7d07f5c796857953a538e01f261d9d7655100eb808aac4206053c1999fb0b2e7e1d12d89e430824c215b5b614c2b35e77254b7f7c76fc99a45e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha16026891864d94b926eb53898085385f4da2ad2bd5802b457f724ee63ec2bb035b06b3fdf1647c905b858aa24dfb5da022a9252157398b8230cc68aa9336531535b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1caca40dba338a6fcc6008c8a9d601a21c4b7ae6fa2e7a8033ca2ad33517082db51cedcb0d93632875074e8b40d1a83b84bf44b283450490373a0a7d133a8ef20bb27;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff80ee0c968700588373caf373f412a576dfeb7f68a64288f05c30131423fa3567e9a3a18050412f80598a06de8ae87e2795e8a2d82d7f7cf1b6204e4c5feb28bf08;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f1f5dad3ecf083682f32872af5ee1e25025092bb12d905879416f1ee9d88568d14aa4e19cef4637dce93ec52eb2c6cb6378eea6904a4f4e9411785cd5ea1985f84d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6024fa5c7abe91d3b474fef20edd6d27b11c32e5d3dfbcfe04ea5ddaa568bc1a34443948c7a3823ae1cbc9bf3bff4db8749097ddc7dd3e702e55cef20cb0fba6c8f3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a3662fa992dff8556f813139496688b64350843776f7901651adbc2427cc614c8a78e4d501460782202f34c7a68004c5842d436cd7891258f03251da60e0689e140a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbc8d83e1174bfbb42a9ccdef28ae29c73a8ef1aba8b1f042f234a4b95f123239180347cb60bde00a5340d36db16ff8c8573c73258e8bfc0876a8b1b04e402fe71a86;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha656cd241519388f755f7ac896197cfd450ca3f71fb6ed1f37c3b0c3472b3ec67c13b1d9340affe0f49b0a46ec008b76fe7105b101c6cc26dd496d64f07157527fbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h104c6927b43599a2473fffae3feed6fb2931db7543785ef9f8f9808bd12daa8faf8400e584019aaa32a9adf140ac10085801542ae7b1838ba885ce88e70ceae406922;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h113fea5668f606dc9c3ab900231f14182e1e294b4c96728d362c937aa562d76e3a57553bcff2ab0e3921ef8cec510876b61bdc360c18c608bfc5f722474f5b04f9402;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f650328e1a3c4af236d3113a91ba89520ebb117483dce3e8caf1abe03cfc2a646335ca4e3f6bc60819443ade42a6da60a47d990e5287eacc9a50dcfe2eb7303a15f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf2b66af65c2941e0ea0cfbba1ec465da260e4db44f4c1552df0b2d1d403c71525c1f02edaac12052af9a62d42d64fb1cafb1d8a06b45d2691bbfdc012f9c6ba74f80;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17130272e80479be990e96327c666d2658475e1978057f388095d1854ea0767c99534dbecca6770f36b0f302f81b9a8a293751c1859660d2f04d431a6ab85022b8b8f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4bb3a1a2876d6cc8433b5f82ba73267a222a6087ca36ecfb2f523137db0224c8c02d0364e522e1f673458ab3d48062a65afabf7f3993dc447af775d2b543b25c70b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf631d45164211d3993d41f2138d307180d3f5cc253bdd878a58200a26c9884540c515acee0884596ea30e99ec8f9ce00abdea077be77dbfba61f879ef8699e97587;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcbef8a811d3b63d111289b437ec2620d2bb2478850dde2af796791de3944dded6cf293359b5ebd39fe0ceaab70c4ace6f2386beb69fd29219d1fdcdd915d2595e331;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ee2edbf6ab2b0a08d36ff40350ae3e7bf55b94db4a5705b4a90b02c44c50fdd48be690939aacaee4689de0c3ffd0c51e1f71a64fc324df0b364d6d6ee30315368cb2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fe4c3e1233d548b9a7011ae5fde8325bb32518feae53c0daf704615c2ab329d7eea7085a133cb6b0568d4b7b7316aa159c2987a10a7a03c9ed515558cc4fd0c2f512;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b160cf3cd64db8036b85e9ad3ab07b97bb7960c52ec3cde1b9d6c3b0660db4ad2e09e529d5c1d42787b1b854d48a3232ca68c9868040bae818803963544c04b37608;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd73f51f323005c133c8ebd667e48c83ba1b6d2d1a8f21231f47647ff1c73e46c2655518833efa7d1495d8cc67957ad3b8b463ed8a512d52d16314db38b158ea392d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc91790e5c09facbef21f29928d92d86309ff836d61ff8aa667aea351b62ada6918f6df4adaa04aa9e7c29837c62ab7eac699d23794a343942c8bbb1753c84359cb19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e05c6317924a0e3283dc6912ec9e8fb6f4766648af0c6c02a59d5a0c9226626445ac567625fe7bc0d8062d655d6779d6ad4e8e27c08be82d1eee8052fe1525efd22f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f7dfc7220f17898984decfce9bd05e96c33355f7dfdeea43fb45236d0615b288095684396b510dbf564f0d5def6dd53dde391127623417c3d7806f8a350424b2db0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12889d86546b79c0f42ab647e41c0d7fe6e9fa1d02c195080e7e9ba870f672717f92f1ab1bf45e4ee18738a82375de526e4358597794efd5bda905dc9d50fd5f89eb4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc104d60177e06f0e0fe320cb35a2627a4fa4988c6abc76be52d91dcbdc5375f382d66c48fd51cbeb6755690afb95b8e9fadd1ddb6a0c11edd6fd6931d3b6361828c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b385cabb553a7e92289ada83424d0a21e5e06bfd3ff1615733c0c3b08701c2ae9bae4374be044ea38f5fe30045b1508675dc0a5b5c7cf7b52d0a53cf96392ed536e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a82704bb717a7565ebb0a384737f8752750d2904e54cfba906f86f3625e8bd60b9fe8388669c48ab0f9b222d7b4a98134e5ce37ef6b491db0f7ada602397053221c4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbed11084517980371e925bda621c224d59d0c69035e1b5b9c7c52f31a7e1108cc721d46f438095a90fa616b1b64a1318eecfa9fb3a0eaeb606eb96e40dce557deed7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h151f23cdd6d81478b6739ca8f308a6c7c64bc2b880b57072c4c4c63d7eaf9998ad84a2ed08c8a5244daa7b806eb0648f77f06dbb87f052063e1e4d047f8506b4befc4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf50fdb4d15eaffa99d2fa55590bcdadcc84ff3b3060dc5d411ec433cb2b18fcdfcacf7479876efc0b0c9d8b5d876eb919e3e7d38abe9500c590fc219b06ded699e0f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e88fd8e0f2474be915a50d0f151d823c8972bfb6acded5d0c0742dcef8148d315c787ee4765da081439db34c38383230d05020a84d64b99b56d0f5545700c457db7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d118ac9d4bf6b0eee477f19eef091e8db227715347efdc1492758b98059191a939806b6c8e1ee56e5f99b062d75abd3451a4cc6c023e69eefc380644edd8847e4fe1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1014f3d1efa43f49855e2201a3df1a901a12f6647947e9daf4666009621ce963a3600541bc56ece8378f2b085622043e703dedcda4687574eb53fed3c917817f56824;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h50d46d9930e340be3644e8aad63652ddc47dc26cc0ff228ffeb3e0469db3ecafb97aa6856d113b302c7db81219516b5dcd64b4bc50971b83e407c16d9064d2120d31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d16235cdaecf5ac83242c01cb4c55e1abf13ad6ccdb51c05d26b17678ca8c7b77a17d45eed10ff4dfc6b468bd2b12ec115ed246189440385ed1f21517eb79b382862;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1367ec3b3edd1e2b7aacab78b9d5410cb847924d85304c1bff4f2309d5f9ad09372b0e032ad51459b0c4b9ed234e787a889576beea8be19e168ddcef83265e107e5a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17c8516c9de6965f07f2bcd1fcc0ac9bc0fb0ff69d6a43384488d0506788164905fb34106768fc7178acf2420545e3f25e488ed2fc09da6c0f9f4adb74ca97cd08a31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1df5c86893514acd989b975244613739fcdbc88c5d49a140e6f408fe989980b3057f1ffbf7eeada279d63376929bc7134e6ca8c4588cac3864276807b8c796427dac5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c4d0229cf63196648a34db431b7795371f927a4edf3fc47295dd43b03cea1327123d1d3c2a7dfdbcc0412b4dfce7a774ed4284bd65494971ad410cabf70f01b4503;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17844f896f5e0bca7f8a836e4effc0b559c8b7f41aeb1698591f2568975f062ee3fc4d5e72febe3720781b4173cbb7e1d4e3cc7cd9b3cd86a197ea9b04debfd62a0d6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2153e97102673b4814885af5deffe3e52b8f991f98efe5e250707b0e8d3858dd5dbafcc99fb40a55faa1d89a544b77784bce2f3463a37abad89b68de12ebfeef120b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193e6b2245a5d5fa1f8039b2f1cb25d09af6185ef166fbcdf78c7b5e94892f485efcf85c074b2f75b2ff4610022f42fab146ae471ad487adaf4e93597b4b27d02db1a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf14fd3e9162327f59ed4114c8191c3edee8c91d4b31843543ce9e9c21a9c64775d965e8ba712aa427c53d1d9e4cb271245829eecee7e32505a561f8bd310237a648a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e821e2d0c24feae08f508f322141dd832f7faf86faa18d5b8f6b311b7a1c7f660ffb80d5a72a35cb499f1fe7c79ad0face545187f647de1c5b514393179d5b75b59;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6dd73266a7c38348170b33fe2237b4e905aea3a5ebc0d3ba600628dfe566f9422831edf604784a556856ac00747f9a521bad69983b1582dc3137fabf984404a3c249;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf60199cbe1d942a7b12fd0d3f54e894f7007205919c687802ca074ae9cbcd742e8ad082e1bb4f90f792cb7b4afe2ac5c8315a7e23d7be24b2ef5fbc60eea31fbce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c399b9373702c77a9e4974a2aa7af1008f1553ec1d537dfd263c69239097c5226ae510c5f71afce9bd9f45c9e3cf6d11e1fea0efcff2eafa43a03411a26351c8d90d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h537a89a342b107f1c9641836e4cc42b8ebc3ca8193924c476ed2abad424f5aeff6606a6fee4d350e555e8a7ec52a60473ad09646c89006bfa16a87c9225970584708;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4b172e1f32a79dd195a6575eb67bd8971524cb048f014c8fee9bb56a3628405800f54e26dd5e36409c33db7710c7da7690b5d56b5750b20adb0355353cdbcc9407f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3a50e86af1ac0391ce749481cf0dec5e0168cd8657f4eda21a05ec7aa4fd8e812058fcee08d891e3bd1bd9aa4bb697e68909982803999dbf5afae15b448d7dcb6ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8871afee5bad19a1f778d32e070ae4883af4c49a211ddcb9f4fc5266f9653fdcf08029be1e8a422a8e5b6b69f37373a3d93f9b8e55544537c78ca0de1ce7118274db;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e4997a098e169111d86fa66a945e7ba87b0de262fb7e3a2e5b405043fc2c075375c550c558ad15cb5411fea63371fa669e3c06161aa1d64d9c304a67d628a1156f0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18949391fb1293f0641958497d46e3237f1a2b789a4b1051a70271d1f6b800a6acd246afed67179dea506292dfe373ee42dc06753faa3449f80feebf55e06a51a68a2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf4b4a7fbe8907f837e16c659f9cb1e5f65306a73b88682226f37f5a592669cd3c67d9ab0b46c0158a09d8d7d68cd97c1379b5121ec7792051d6d606b05e509de2630;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f82830602f60e90ddbb358afb3cf848a339f6d376a4d67695f11ada95eb489c14897c96730978e8dcae367b92ee116e6163d56f30721034745b7479f2f8d4403957;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60ebb0b483bec73cde2d83e91f226204bfc9df7c603cc2f7873719d2a7166e93887b9e1b44d17741cfd38353b2b3a6401c67d0f1c64e167575c97aa1ad15cccefe35;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h349c1f3370211881d5cd3fef2aeffe508764ec3a644bf54722f6e5a203e058f77a259d0ba17a9b48a188bcc11a13d85bffbf55696023997507ae93db53c6cca1261f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd6dd32b3ec3c3ee82a13a89d3dd53f6d9ab570bbd9575cb14235bd0fab98d2eda46a4b7298708fc2325c575eeecf2228c933a32e7ae6b3c585ef17bf78f07439197;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd584789e77ac2c5edff4914803a632af22f5f77ed8f30a66bc46e7b936fb180f645c601ca493eeec0f1eaec21980539d1232a374e78022ca3363d7113a6be28ea68a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf807964a61283edf7335889e00946c272bf849acaa065ca7ad11564d49c81d82c50100225698a1e412188996e8ba1f5c37b7825f3cf44226b0b15677f4ce695dc142;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b1edb1283a43b746658615dafb5af06d2b7884443d4dac8056c64a113c612a817dc5959c90b31ca363f4d8fb087a34580ca21a6bf8fbc5740080355df57e68c27b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1353eaa907657a263c560b45771be2afb57dbf36e343f40cb5f5597cf8e54d59e7649e545018f642e6b5bbe8989ad221c6ad65f6b240ebb30328593970bfdff903bab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3a6f2aeb108fcc52732f4004018889b8b143bfc0f416c220f4b357bf7f393d45e7bcc9abe8ee805586c7ab68b70784a4213fd373ba74ccd03af43bec93253b3da7a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb94aedc1122cc6220d1ff7759965738e7b4589dc60ee15ad0e2e2dcf8d74f8d0df702345b5c1b9e0ea1a7ef4d356d7ff85c9fca6ba1df4725e7241fd4f04311eb1a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h184c932adf1012dde43091f3aca7c6137e8359cfdc2f89d8aa5c43e9a7b55461b36efc6bacefe70d03ba094c387138d142d856a68113b893266c3c63893aa3ee6c813;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28be151ff5f9f2ec88df15cfce896bc58eec4dd7b5fd032b3477886d8570ed4ca56e1f8a1bf0407025c18296179ea7df5926347f14ae03103ce0856f6cb04a15975e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9a541d82887d342b5ed8b513a83a0977e39e006707dabdee0edbf04885e7b4e75b1ee0a8e243500d8df33a54f7a7631935ba1cd6b7ab6341b8cca8e592ee545555;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b352cd7295ccb43dcf4fcdf1f0f75f5522c2a71b4173e2c7fc786ea04b852b6371fa9950f23dc65a23799f057136326831330cec160bfae05d7b788856cfe4ec3ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he16ebc1d8e3c0887fb83801ed2f18422407fc46370566d589bd82535d2d5dde4405692c1ff158ec5507caa4bf3830933f9a02d76c1986357ba8241f08ca4b0d701b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a018e8fbfbdb5b7da7be915b3f16b5ec89cb37da4ad132fbd3f3ab98a782c838268bcb51567350dca9478690a447e3e3e55ce361f53f1ff33ca099c39becd644098;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34c5ccd4b92af45c2659abbeb4859957e6268c5deec5ca6dafc5c17de4e5a9778e467df47d59af3fbf1a27ae990d7a029d0a8e7fa0564a6eb1810f32ca373bb08a2e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103493148ead3d280233936028ab3728dafa9145f8037efc46ceef083a076cb294a9178e0789bffb50bba5c9764df0f012eb6174074e4f967f57a43bfb9715f0458c3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3085991a14964a9f7eb9d85c26b40315aaab07952f08ed0a1c58938ef34e26660fea6ba77f6d8c8428dca96e2e264348f8efc9304fc8c0c691c7c16e448792794849;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3ade5c5bb7ac464b5f2b3bcc9a4ff1e34c73ee36823b95450086885a81c21e2cc052dd806eaca25496a63415255cb0e5876acce32653a08f8b2de4775d66fea25711;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1172f16e70f8d26cdef7651a6080c070e5a50c942d7859a755f09122f7e40f4a4026b63f57731496059a09f7ae96c5b6fa03ef90d9dd4087a130431491b4e96b469be;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b044b0f6ffd710b51018d5664796a1c3ffabaf647b8b8ef041c29d93bc8937d2bd1138163ddd424be015bd863383f0cc047a1890c6a8b94dd587c1760d74d009a5f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h72da00680a668f239c340e232c839cc9083baa623e36f8a7721e784fca6334eb5efde694034458006a29a3439c47f53892f0a708a0a3d08ab78ea76394374ef85f28;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17d60ac5083961a64884758d323153e816eca37da1f66095d2d8406a245066deefd20ef98c1ec73a4a2eed4ba7d875b4b1430443f443d057e2805c94df65169f46dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h30da3cddada39f3ff3520946a2641fb418b1c7729abcbc8b62c55f16625bddcc5095ec57ef473c6f41e7e426ba37fa8f0d75a510c51c86a13a31017a809bfa433c4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbfb5c39bddeb325631aac377208ff844ebf6df1ef74b3b26e607589096daaf3abd9822181708b75fa63df59206ab7c204c93129c2e5607a7dc478a8ad55d14815674;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f174387264a53627253761d1fa33fa289180234c5503824f3c5e6c858620447b1117dc20bee14be6476cf82a295eced7c44ebd15e3686849aefe717054040abdf21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h774034188641b8f37788ae756a91f612fdeb2332f0a9222932952bd0a300c2ce864bf4447838ec7b8bb8aa0dece02a2d6e6de1c11bf36c163b5d59a94c4c455e0f0b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h64a10f79fcdafd65fe1f402eb590b6517106ed0ceffa75e7b6282f9e1a3ae4d4aa9b3798ba11ecc19bb1b62e87ab661f68409d2cd560ffca82e159d48677bb00aab3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61d2ba9e398112444f4301270126a1d81d513b30d27d0ed2231bfe1e1cb7620c70ed8fefd81ef9e1e0e9b4f536a87f199c0833803733580d79a6852140fc06966d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b92cc977e8e60ba6afca29564ee625d0b7d36c9c855980b78eb79ea7c438c13fcdc42e7f9f93805cd0876c93b5b5976852aa4324e40219d944da20aad42ef626415;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4458300ae11fbafdba58c85bc5a0199f0f89d9dbe1df9958b69fbd472c37d9db5e5ab21042e9a0fea05911b01b291adc4ad0a062b36e7cc31ac7170223901ddfc1d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fdd3bb85bd7bb923fe2026a142f9826231003eb2dea8cee06b26c0b86c09fe45171602e081ad3cfc4ae507cc49380b6f2181c8090ab6e413be1fad42c77a4ea65159;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf7331ebfbd5f7fca3a3fc93b28a65bf5ea50a8ba0118ffa97dfb9f77ea6bda9ea8c2cfb27012c57e35e880965ce4d29c874d37326ff09802f1673a9294aa16ec29a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a05aa50c4ebb1892b7e56674718c691cfab30c1256ebc9604bc557d1c1c351ad9dc8e4f7722cf00c514f0c90a3fc420e038ae742a73d271d774c68374ec3d88b3f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6a514c53a8bc5e35a5e73fc491388e0b07c403dd3a096889e668157466031c061242c1054660a3908948bfcfd635b3015282b8376d0154fc1f53acaf38072d1a3f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h196bc8c488b9b94ef133f321f121a5acd7f8c659b6c74ee85312ca9d8de28763c66a1231dddeabbf228964ae584c22da21cc869ea5d77b5c513c068015d6218551b47;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105a8278ca06db82fb4d55496143427726997e604bccc931b7cad84cc4264bec44c80c6d3c23ca5a9f634f58a54661a1734498784a928eb458fa56f06045787bd0bff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19fd0d4584628bb00f44069ac7206acf503e334e5751a84fd43d6902c6de6900815a1189e7c9149e7b42c219bf25118925422da581b81128a779a9e74f79cfb909013;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4c94d1b815684ddf76311ce30135cf4bda27ed83421ca18ed5c04a9c1c8e3466c277fa69101daad22916111331c2fd6864a56fd24d24c673ba392b416dca7af4af1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19701c69512ae633a6c22505f25dd8c939be83fec6884be385aa2c692ffd1f135a7286ce21e674fd603186ca7ee6e4ccd3eeeb6184464fbe7242454624fe685f402f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e1897713eea660c427ff9d50c84e82c3d99d5a68375fc4664d0d6d5c5856b3ca751f0dcbfe3fda4d9d9f7974104521e7a4a9e38d0171c73bd08bcd3b16ff7875ecf9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h147e3f3b2c77a9927b15a902784951771c38d871cd03939c8b3d0550d98dfaed62853278235432037ccaeb15089f7a493ad479d421e0afaea451686e1d11640709d1a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd1038d2e8621c950868d8ae14b7761dd1838ff381d3c23ace23bce88ef1aa675161956691847f38c618321e6c063ca60cd8c64173a1d14ab6c53c668328478e33c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79a24a71fe771705e6fc2f316fed86de8ac440e0c790fb822723b5b0496220496e4a95012f37383893c6faf353b6892ed5db9c357b77fe3aa3bcb9f28c4327848b14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7da06823f488143fe203121b587ec4c5351490249524aeb9580a172532c9c9a73dee0c1e52059f73eb4c27b232a0570f070e4a89a668433207521419eddb440a975d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h357853250048638e0be668516fd09b355b3714707779cbcca52f1c425e8d541428959c9bfc38256203bb1df47b7960f9c758db13cd2cab8e5cc1af3b525a8ba33a4d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc923cf481732f5f7d0af7e8ee2422d778b37d7c6336c80356a1e8a08a37c6a91a3e78f4af947c18420a3af013497a7964d6f77ec0dc67a9caacbfab59b33442e3dbe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c787a546affdd7ae05c7e6367eb246bea472e93ae9f57b06195789751919292be6c651a2d2212b07b2e62ea006c504071e8c3b3c16b419d57d2d6543fe0aa3e924d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc2d7f595d80b0c68267d306fbb12608e28ba59f770bd9f929da5988daac8213c72efc4f0626648ff3b0b380852a83f110916412fdea1878f7bcb193a2dda2f2a979;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3e9b0909087e99cbaf54a0944b6b750f10da7267d68f0ef2f7bc6a0ad1e0b572ed967a1cf2b690304c904e1c0f5f56ea18b2ea78541da112446f6f8570db9728edd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea321b885a4b877c38089ec91c1b04a0f5fac3e2eacf06e6f3520ff2b7c63447ff85b01f0f478d2076f47ccd60ab5db2826980ce34b3e8794539ff52b89a5a3c4a29;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10889db8f5a592a51b4c1c17f562b4ef79c7a723ce0c8a904d8d680144160a2d1166878e4685d67a47f7906b109ff33b05280c39e70ec88d9b2bca7fc236115849e24;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c56541b45e8bddd4cf56a952764cfb5e520546c04864b45a52ded6cdd62749a72bd1856939359645a4a4f743fa43e309a1cf2a2d3a4e839bec8d8c1898234fcd3ef3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138dd794d26f83eada336aa2c6567952c49ac6b8a46a489411b778202fc59937ac53dbc57b88bc0ff06e5333880f3648fe327082c6e9859c56f03d180eb1bec5337b0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f9e188e4e67a791f12f69c0d5b19e3b7dacf202b42ead94f393edc9aaf359f5c25106c35cf637bf0790dfee2572175bd971ce3231c6e585d2edf041a10530c01219;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a4a62077fb6f87602d715cb448a9aa2116a34fa8a1a1dabb57caf26ef09465daecda51492b1b84f9634f646d411139ea5151ec91eea66851e319ba9326987141308;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7a06facdc3adf743181e9156ee450560eb7988b7ae53599bce85df452c582f29c5e544696dec960c73b8fb14f12d68d3db4c2c04f4d080f2a6164cbeab499dd6526;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he70e0cb374b88e299d6f0043bb7e436980d0d60e3addb6531ba163d8a537a8cba4702482b7dda4d8ee0fb87c2ac945fee0ae8f05fdab34341c5aaf99371683f797f8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ac36cee4d7f2969cccf534f361c7b9da6efeb8af2c3d6396225b61b4981447257a96f2bf931055e7774873fded1bb8d01dcfd9a7ccb4e689cc1cd0cb0fed63f2bc7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13885161b88abe72c89c5ad0b6229100dd398ce27370eff8dc90e2144215e1b396a8c6968fccfcf459a32e80dac364c9dbed9824d7b7e11c820198be28df2110bb707;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17c109bc568dae2a1bb6980ec59b6f3fe4df04f9fee12e4d7e07aa17f34b9c3543dd25c4f8f16d11ac118268568aa81a3818aa6bb43fbcf5f4fdb3984a59716c4a4a1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1021eec584b8d82992810ea6826cd8d0c10ac06bba17ee2eb533c623c64269bceb0b32833017bd38eff6a678061ef7481d626c07dedd6b40417f6644e7a3936991e98;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6dbadf80c43996b8c897ea05cd6db2330abe9676c420921a6d3d00061654361020c7fcc26143cebb41b9280d51927dc39dce7261e4ef013caadbe8b5646481baced0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e19c4ae9ccd74fe7283ba62f95b40f7fe6d85503f932296b125937f56c6c41f6a01b645e987bb7dfad82e97f538a44ed3cac9dd62a20f876e2a114d0face6d1c7e56;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10cec696752299e9ed345eb9b322f11994c5200fd15086047ccd0734d766ae53881d81aad974957b4ffdd4a02367304c89c73b7c08c74aab93774a678521629f0021d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11c654ddb9a9fb0d853b0a13b4672f715c47fe5ed5ecc1a788101c6ca64006bdf2674bc1a4cce669b74de735170e6300fda5fed9920b4852723a7a514227f2915b2a2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ab975960898e525e575b6d0ff8f17b9820e9c3797433746023a7751c33d3dddd54ab810896fc0e1a8b18ed5ea02625ecf713e2e833176af76fdb559206abd6deb358;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18a9e05aefaabf3b571dfb6b9a494d362cd8fad4f3f4d68b88176856a1b0148c7b9b795c855487699e659edfacf5371871071cb0da6cec5a8521a4af0d62884da43e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d579ea2805d8044228f7730ce074d03ab9f47dfcbb565f0b215ed182a9d8532162ad4fec39358aa26e31aeeec68b4d85ed167cef8b9c25dd4830f589762a37804e7f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haacf49690b41f152f769b60ea6e31fd1e337f2ea6ee7d21e367728936c41871815889703483c0dd6383c0a04000aa01cfe6ffbb1c09d950780553d2ff09e614c50a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h159e9bfb00f7a567a2a34f1921a8274b4768f2a2659d01aefa164e832dcf2387b18a192387580b32d88fff24b8012c09e6628f7d78dc2b426bf10a52968368a858915;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1222c09c14f8ba33ef775253e57ff6b7f34c4c73eba1d514af8e214ffd4d3548b0dcd4485f890de061ff86f3c3a38eeb12bf2280672c9ec29ad9b12a3b1eb73e3aea0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a3ee1916e97ec725bafa574622e4d5333317a209b38c096df503daa656969d68bb4c7665764e526da85eb7e4b8472c1d2e5bd1c125d63e246cfac8752480d2fb5c9b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9f72845c13187cff56d79687ccbf7706d524b3274083e44627729319d240472db2fd4569326b4de178d2d6904e75d62032673e25383ab2aa88346b6f866837464;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce4f2843a0e3b6b8614fad045ab155d28ead74c0bf5aea37ddf5fb3d436a68eda6a5cb0389f325581ab597748e91aa7e7baa91898de599601f329bdafa3e2d927616;
        #1
        $finish();
    end
endmodule
