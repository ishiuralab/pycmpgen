module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [9:0] src11;
    reg [8:0] src12;
    reg [7:0] src13;
    reg [6:0] src14;
    reg [5:0] src15;
    reg [4:0] src16;
    reg [3:0] src17;
    reg [2:0] src18;
    reg [1:0] src19;
    reg [0:0] src20;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3])<<17) + ((src18[0] + src18[1] + src18[2])<<18) + ((src19[0] + src19[1])<<19) + ((src20[0])<<20);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ffffffffffffffffffffffffffffff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e630d38f9cf5ee04d10e2117e4243;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15dd313c68c6b750ef725a2f60b52ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce5988feae0c62463335e1b2fb59ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2b379f2eb00084cbdcec63165a69e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h534e82a34e5b6770f41adb7f7e9e6e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6f58f8cf8dc40afc01cf658f09b209;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h737c3933f4426ffcf76a5bcc93ddba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c2bf679220a14a178ca2070dda1ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8b1d5ed7836250a89e70595da8b7f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ccead32cb34307b22016f2b91c7b28;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a2a82d62808f6cdb884f3a53d4a58;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h103eed91b7ee411d7cb3d12b4273ca1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hef1a9fafe6b2dda359f2b5ce10b979;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3baa242957fa0b05d0ca6b0e90a086;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a930d0c5f66babfdaf460c9c40002;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f79f044a95fe0f8dcdeb10f116c45;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c757850922037d7b04ac9b8f41cde;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10cc4e0c5dc22c2fce6a8b17a197b29;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d8d7171112274ce416227b6b44896;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h190ed28d4c82004482b0ca90ec7bb36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ef1635be65f5499f8bb05e0abc959;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hffa247bc5944718016bc078c36aa4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1630d0a0900fd4d16634d06c47def0e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11b57058e4a33fee231822dbe4a7251;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cdc1582248f087fdad8b2feadc7eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h181e61e1597916b3b6c918c681317ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c376ccfdf2ff71eff184edef7b331;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ffd78a53ced3882fbfccf3e02bef60;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc138718245d8736d949980f8f79191;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19c4eac2688ff3e409f2425c9f3ee9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb21d743af950db82a5747da52220e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec37093f71cdab07723eb8e3c9f007;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h840f89ffeac8371e0a8c2a2c7fbaa5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9ab18af1fbc7592f8594fa8d7777fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2a001ccc7fe4dc58fe9ee13266c0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a8a42ec2bc0e61c5d18c98899fba2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcdb139456bdabe0aecd8ed19f766b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha591687b2019f3de738cf8efa1b07d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fea9ba8b3b0c1925ac88ec8bf64a9f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h192bbde57524658ca4cd203fad24a45;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd88b51a8eaaeae3d2e3cb2786e6d4d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h85f8542c02a308ac61dc4d8b11feda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h891dad50f04e26b00e6350df2b65e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1032657a832629cdafde2eb9aaee905;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19f8f13939aef332f169f2ebf546e94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f2e8800473d3907245c6b077696d7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5100daf537f23a223d839a59f54da6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6c28eebe7b5d3571fe9742e1be69f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19be088bad54c14f6fc44f7db73d94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13cc7a7d85b8ee7dbe2f5a031746c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11bcea82a27238c61cc4279e48442de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f202a9cfe3edf86b8e7a2f44d5de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c9ab56c28bc2526f5e82ec1a7633cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82ad648553c084a8293e2935df0b31;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe5bd319e6688f5ee524a911771884;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h52e42e4a3561bd845badfbdbc726a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h51aac4fe3b9ae61ee62f6a973e0059;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hae004a97b62f555e9d6556df230e1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e9500a82587be531bc9c7bce729162;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf2804fb659395b6cc75d0827a2853c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14078500e64ed967ecdc427a8a44e8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cae119a7ef8c24a832a8eb2c9de36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145981b0b7199d4e373ff82a15d0005;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h407ec7cdab5e8c2059d1e9367c47a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c77780d981221decbe4d57061db5c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19db980970b3a241e0eedad8e78cb02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hddaf17e142082833e55b325849adaf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8c1005a461632540c02717ff18358f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aaf3c60d6d3cd748e78b52874a3db2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cbeef9f287d802629211aa7f16946d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8c8d1c18b1a7961c3c89fe1dd3548e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11f22f4f47fae7130255adeb0aa2d29;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha9ac99b4be6c04abe335787d4d36f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d5c9e15544abf9f4739addfce53451;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18696431025ef5dc5adbf9e8c105d18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8f0b9d57ae9eb368e4018e56b94805;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb108c0d203ac13933527c228edb113;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb63efaa8c8393f2285e7da9c0aa39d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1704a7a85c98d5ba3b53db4ab49bb16;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e8d6e703f4a91b47546da88c43ea3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf5af1baf0fea4519fed68bea3777de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ea4b1acf837e10e2371f67b3509aca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcc6ec6c68dfcf59f1ca38c00198c95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha7eadfa1bf57fc493efa41ee1cca8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce97df66a55d93fbed38274a582e7e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18e5352d96df2a262bdc49737a85961;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3ab93972b0b75f3344488c58ea3fd8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf977d7aaba522eba203e040c561cf6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b1fc20a87e51e3ef0935860177b45e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18da1ba1bbdc1df22fcd5cfe63d7560;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a4d3cee778cb93858e88c219dce47e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7f87b177130de2ad34c0d01a9cdd8b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6b7947b562e6e74b7fb96549bf80e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5e46be0b35b2594d6155ead3882d71;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h729be25d9050fa73306dcdd744fed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a6fc005f5c9b9589aa615332e40844;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13dbb2eb7bd9fa1f5812aa55b04d41b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h627762217ba2680974a5c0d0ca323a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2c9f1b5adeb1a94a3cad7865b70fe0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90039875f68e6f869a9bc70ff8abe1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha1adea9b4d081921e8f221b033ab7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f7bff4467d0bb52a80e6a5d3c384a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a9f3960918ab4dadd1890b70c8f80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbbd2c6eef3f9bb924785449711248b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19b817b7f64128637aaebf051b34bc8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a70e0f9866fb0682ddb7b1308e6aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145e2955e4c7cb1a235efe917a31477;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4e85c3f79260ee7b2da5ad7bdc456;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f10aee2a22a0311315516f94b62188;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfa0c58daaf2c7326f06ec0a8a204f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d9e039982c7156352e12dd874c85fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a4a433162e4a320636a9dab57873a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf8ce9d71f86e865fc1d1f8f6e73ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h135a26cdde1affd95bf933eca78ed24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13e24c52b6c269e05e0894450ed165;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197a6424c22d59ae6f684265d35519;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2c6365aba3251c672f4d19b6a21bf3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f0277bc5f63440b0822c63fa2c081d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17610b58adaa881f139577d4d0879ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb7e8207b40a2883b6803d5ffb7f23e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde6305ea4fa0978abff0916dcef515;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd55a6c26a9ca555f71108217ef5e2f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h140712c3e1a382fbdeeb2fabcb7c32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd6b4319557e17ba1383ed370311bc0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbbb759ea20ab2dcea378cb1432368d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h96b8ebfab9b8c7f2f30c72f1eb15d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h175aec1aad53c2cae41ec84d2909bbc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h60a6cc0291e55652570e29df42a8ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcf12e0943020d922ec16ab3e491d93;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2703a29ff14416b797458903cd28c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc546440e23d6650a518cb3d9f05318;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b8823fd2d1dc546d84b6817c49b1ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1292967b82d1a3afc2129546679b45f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e220b47c9444463bcef2816d99868;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14e20158624da3ced58b7a2340fac42;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2cf9ee47b068550aae413a7386cb26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15111feda7270845df8b1ea1284e978;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha8bea5d1aaf27fe3d90857960a7c61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcf6fc2cb794c2451b6fb145193d426;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18dcf4efa9f757c614dff8938c2f8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h478371ae16ec14db8236d43bb630b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a92bb2c4e6ab21990bb27303ea5f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfa51d700b5f63962c83805883dbb52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h114454c616231023ff0652fa63e4310;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17143ffa82dbc8be24d119f0c9fe0c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c13b09d73a874f4a851d3f0e8d3fd4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1092e945204257f26a4fd8066310935;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2d42da1103a42cf4e8a1c1e86d59a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f2b28d4478fb007d2acb27ff2ede7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f01fa66237103bf5262eed5291ae4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c5071853d35ab6d7e13b9ef702d291;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f701ee625c97cd8d05e139a35ea163;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce669a826b6cfa3890c825ee8e1de3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc6297385bcdbd882b9c44a2b361a84;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10fd05332b5a8abe9c17c283b7dcaf4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb3ee9d9be45cae7907da6200286d47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h154564b89985049fa7f1f88844a7bb5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f9b7fa9cdebad47414a1e931e2a4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9e2396c123c1c871537bc633fd0f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c45d06d15bf253ffb8771934c64ef8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5189a3fae0ac0fe40ce5224bd85e7e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d44155dbdd0554216ee1dd0ae8d59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e6d7a7c5228bca4581d86ba2b9404;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h225a0bbd00e9938977b220ba442bb1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd3141e4b74a0003bd2a36449dca95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dd83a0ece13fde1d2b6948af48e44d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1412aa2ea2b137437f7a0d2b2f99719;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14b82f2c2d15bfeacef2545192a6907;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19e0725f74b10100db9e7d030c86d96;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h41dbc0252ea2929e3b565984859a58;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17734a750628ccd9fd2b6c4d24cac32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd454b103cd315e3f0a72b80abf9490;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5238fe388c1b39618e7e5708c5293f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he7ab49e28a77fa390903d0d0f33894;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h80e00689442d4c342368b3e55103f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2268d3fd6693c0ee38bd7266d2df20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc47c36509ba19505080e519cf4cee7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h743eea57762fe07e76cea2779427bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hadf94c861360a2afdf687c64def9a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19af1ff72910569ced8ed5e3889e6d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h39a47e4a1394bdc3ff8950d6c2fcf9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb301e28f92e0e16d2a409ea60074cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfcc97fc05093bef8e86eb0f4f81b9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a8b157c363d8d5aa864191d84100c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ee63d41976c5d35c263e754f2ca63e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h142cbfdc627aa546fd4d9f2bf675aa0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd66ee6e528a1d3f6e9f704c60185e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hccf733e2c917956ceced39ae72f8a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13663ba3689f0cdf16a74dd76290ac5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f286b51292fe259ccee200b715ddb5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a9b3551b70ddda09e84982f7577ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h344baccca917215d34b9f50daf2ed7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14d4497cf973642aa4b711b2f6e29c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdfcc741b744f40d7e92210fccd54f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h148621ca7501a41d9737e9f46181c4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hffeb0be0e8b2f7c8aa3583558c4a36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d96414fc054256873fdfee14bbab8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a7c163419c41cfc36eb1d5361004e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a2445d5fa3c103f24da25b0a42f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1249dafbf8bfddd8d6e3571ea3e124b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd770d3f4c48c6cc645e2957113facb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f90eb84e150475cb07ef9171822cbe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha0d2001dd500b357eff638878a52e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b8aaf2cb5ea36861255a5527b708fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5f240f64f7b59782bab697d019d94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c08dd5b6871eae121f42325e66f49;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd7b805ac826f411145e893c6396554;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b5bede69acb5f270cafe2a487e17c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138a5463344f2bacba3a0afa989a290;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2e6347a2861a5aa8cf50478cd38ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f7d2992ef9d4a2f44797d539590354;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4440f15fe2fabff5bd3ab1c8830f9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h177f9dd3b070f27ed0a79bfded39c4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h102070994d252db3e26de1ac4878386;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd29ce749e5956d508c8ea2ce3b76e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'had42d3f653663d1299d0bbad5d6c3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90e8f0d3bf34e24b0c98e22ab2c32b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a9a739afb2895670cefff122caf57;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bba879f74c849df16e6691ef44b18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb10308d4252e63794b50615496d591;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a6158c492bd4dae8367e741be930e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h166cb0047a13c5aa108127665e57bdd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h133d221708aa005c970a4f8af103514;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1208fcdf637ec58ec0c36c12f560968;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h130854e151b094262b8feb47bddc516;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138c2fb39ce84150eb0d29225897933;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h69a736731f2161c472e52127de8bcf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118e38e88e0d9b1fa356463c5a8090c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4e1e382c0fdc443a42f1f349713b3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1135ae54f207de119aed93fd95ad4a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9fd5e850b9fc7bfa3b896facc49e4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d8df30bce4f889a530edd64e20f98c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h650983760aee8c7a6d296685261e2e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d9c079a5c5725a2fff2430183f4a51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5c695086cf6234df6139bf5601360;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17a47b003d07b5f0e2392f96347f330;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h99aaa2fddfd0ce519e367c27db8468;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d81bdb07df71af29485303b6699378;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haf5ae92a81a73b4e36c9709546e4cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d78d9dea2c98c4a5463b2ab3d0bf5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145e370318bebc63a42945f250c1f81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7e4cf2034d540c9fb84f815fc48030;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ff4610e70a451f59982f832890a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1abf67767125315dc5d927e02d8b175;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha34a4fd6954b3f7942c85a98c930fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ded979857f6bc043d6507c77939704;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c1356f2e163d5ee22d1993f50c4d88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19f97e8b74a00979dff9646f2388d89;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138732844a95fe8b7e405d48b674c88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfeb9df5eca1cdba1fee1a0eae8ee5d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b18e971fb505c2a1a2f8c0cb48b9dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hacb355d925e70c97f4af8504ab58bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aefacb69b50a679b12a327aeba5d9c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cbee834e7b7756c9696cd8b9406e36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h170b21e9e1448bcd323ab41cfc89cf3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14bb79ff6e669b6ef7685e1b6210718;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5a405d0439ff45033f06f3c7f36196;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h130f3f2305537efc86f6771eb8c86ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf7c6f05452e296438dec84f98ea792;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13d59af5f6c444a61234b190f97ebb4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9c246f2eb4e49763dc25481bcb1f60;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138f618ba0752c3213bf6f4b746e2f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e65de03f8d9be059a13eecc2c40f66;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h114ea27c6aa57d010f00b7f99414ee4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h176531b0c09369ee95e5ba3315bedad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1edb9a532423673671294099f81d5b9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13e51b8d8ffe1d820156a0c9ec9a541;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1445d6bff3ccd54ea9060fe4eacc7c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c30c9b1cb9f53328a84d671f48e495;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d7bdfbd44e6500676b98a09b4f8345;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1faacb2bd4f10611630d702f6d1ffa2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107531dcf2eab406a1dd2e5cfc4d153;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7aa5fc1acd39b31bca0bf87dd36fa9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h167cbf41fdab93e8d1e9437476cdfa2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae9c4411cfab21be61b8d7bb9c1370;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha60abd9a50d533905676e3d15e4d21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d389de22bd0a2a2827d14f35474311;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h190b9c0a2939f83e3ca1e5fcfab47b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha25f4fe63b403c2b5fcf605304ba63;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b103f39772eff0466b97bf574288ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9088f44d2ad9a023a85b8766daf68e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c9573d08b48a2a341b8972881e804;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd8109e51908ba8da3dd65a4c04fdf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3ac08dc99febe11729538a55753eeb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19f288203feef8bb9b813cbf8ca1bcc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4195f0c0de74ad05a67de7cb02c26c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b1ee5af493ccf2b133cd31c749718e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h45ad212383c7d7d62f8352c3c8cae8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17fb79f238e59ebc61c23b2f7c6ef74;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16ef7c6bffd528a8b1b31a1a9427970;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b8b1a9f0cfe98f80acbd3ea041acc6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1926c9342c7c0fcc9cb72df2d57c20b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h113903cd25111e5cd9e23c95ee06bcc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15bea0e95a84ba739dd664566d3e7b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14e4d40c2d18c2ba12d6ebdaa18a454;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4242e86f03d50bef1301ee0dbb682f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1679aefc89700dfb3a05e7f7c317005;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5a304eaf6f867eedcad2467715b781;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e5fcb108e406f4d7f21ae02fdec0da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h72ac11f488a7f1f1a7782d1a6fa9d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h148cc3965aade9f2d4f16cee414b786;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde0fa6d74c3136fd5040355ab54c52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1007addb270a48f867dfd36ca8f34c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h172439eeac15e8aa83ee0eadce6a355;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1508d7c9190ff567e1a5317827e307;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c9b29029825530899f75bcd81c94d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb9c26d0da185ba88b4fb345b86ff1d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19bfaa8dbf281dfab22030856a8072d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a95a42606561d4cdf16d76e2e1d91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h155838c7c5ba3a26f89350d92e2780e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h24d3c270fc4c4b2c97bc5a461161ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h302bd7be703bda6426634988fbaf9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b408ccf48e1b722d179321113c6522;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h307813bab597dece7146c46456ddd4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9d22bd93571c51085c09ce57a328f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h152ebf46a0cc27588901d29e88137ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f10d7926f65933e4a0f644a595ae99;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1af02a66577d97170bee119a3e31803;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hda3a74aab95888230d5b80fb7f9e96;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbb04a256f03c1e26c4aea482d76a93;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h50864753f191118debb4b6017c4ba6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hda76d23079050b9f795d1727429bd0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8c372491b4739e822c389d53861316;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h769f815d2befd5682ab35bed11a8e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf06a32bc6911b788119a2dbf58a954;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157046ba4df35089fdb3f51bf7bffc0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h78828d59845b6f8f03471d45999f64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cb6afbf6ecf48288d4fecedab4f4e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ef264440eeccdae4b2f370329e7e46;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f49c1824d6ffb60e9c5f4f9095b0e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17d180c820d23f55b41c2a1008c5deb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h139a20c3df5383ec091605462a35606;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcb6c18de2572f88e0f8fd6cfbea70c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17006df93076f2dfd934cd5164ca50;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be66d04a1f9ff9467fbabdc6b9342f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15c38bc965358dd83e260f970c89a11;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a73a6906f20aa15c10d17e622a3696;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h673875bfd0b0eee2f528045591cd89;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c53b290d92492d6d5c849ed3aadd83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7b7a8d4d73c8a19652cc1dfd1e6e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a5b83d247423980399d3a124957a6c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f06eaa5f8191f95311084f3b81e7cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h68b89468dc328dc42e771d263297f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e413fbb2fc35d120c79a1f08e95a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2c04162648afe191d7cbb3aefb7991;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14a4bf938aba81d38d3133dfc347abd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd982917f17a1000f676064fa6fcafd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h272f68cdcd74e74357f0d4764dd9bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h696e557541755b03c8a99949095be4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8e6c37a3c8b28eb7fc8727ce016c87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ff9805d2366c872659e1f95e8b483;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haf3eb221e22f3f5a5aa43f95e22995;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfdbbbb4239b937b786e5d1cb00df9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h182a5bc2af718b688a255de458e9d48;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dcc6e6d2467f7400e52b4b06d2e4ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1adbbac23c9055ecddfda8331ffa026;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h135ca8de6ec51ec1b56b1f9b6bcfd26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd485cfd901d44a52f78db3ea2f0d3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h103f4ff7740e1b8d98e968e87c86038;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf0acf740581fe59df90bf607a9c70b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cef3e841e6d87f65a81fae0f7f5f80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heb41b02b31f37a6b6888700eee85b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11492f15a83ca3ffbf915caf5d92ea2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6b36c4682aa69296a8432409b63e2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1001c5b71ffc0dab0011e441709e7c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18d61b5fb39f4d13be586c94718687d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d4d7e41e057eb1f41775f9d77722fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb0412b68d1cf6b31f2cb2845ca2d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h906765c2fad1709b38d8747550d2ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1980475126aa464a443ff5c301d6628;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d667cef6207c38991ee4a2624ad485;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8894cf2bfb26be465c2e08d36d5050;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h57e162afd80d3c4669afd628dbad37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7a8067bdfab7b3213c05820727aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfa9bf81eb86e1fc07fa0368365be0d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcefb046af35c5a8c9ca1b3640239d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18e13da8876ef53a650babbe697da33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h79d7c645861ff3e399225ad65c1caf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ba19bca278c8602b5684cd9b0de79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb32ce77a4f8471208329bb7601b48;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7e9240303cf4c9719d95f4f4eb17ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he89a7396fb1ebf81b2f63da54c9157;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h72e65fe2f02e09ba62622121c87232;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10f315a68e498edfd02fd48c1227703;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f11d1f18bf7f0aaf0d3fcb9b118d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e27fe26f2971356ca96e424b8f2cd1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17a76bde55c76b3ee85f51694f797a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e87fc18c92eb1be34cdf91c9a13a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8097ea71553aaba7496541f84925c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc58887f41ed48f1fc3288013248ab6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe17e8bc772c45c54a93da394de8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1feb6435a54be74052247d7837e342e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h898cdb30d5270f6644ca29831ec028;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197480dac96406a742de0ba46bfb5bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e426a5362ce104943373d488178c06;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha89bf28de460578d2e482e93153f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hed370b1f02074c38d0abdd1283ce39;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1faae0e27d21d6db4cd075f35c4f677;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h196fc56177c9bb9f5dc8d3fb3327a0d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcbe4e83b0aedaebf5a26de15265644;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11cb47b0323bffd8f613393b34590f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ceb478b4e31cdee691e1df4a8e94a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107b3880b5dfa57664e7494f9521294;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdc8f5cabd5ee0b029e4b2d28d59554;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h729d10312fe9d5e06e42a2f6ab596c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2dce9a05a43af285c8a9e077eca0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19fa07f169b42c9d283d9ba2a17c28e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h680108a6ef5f22bd8f399e4a253399;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1388508f0d4a116b0b23b3beee26593;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12df691561b8e124bc2b9a1fd6cb3a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1009784eed818a92780c5a5ea131e33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1742f6d2b1bd53e5757eae99e427fcd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c00c95688e19203690778f3b5631a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c05a0afec50d1eb06d4a3579f3770d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h59cd6124e7138c5058ef578d32268b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13e61202fd115543f36f32460939918;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145bcc16f9eaf507643335ea0faf5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e8c5a418d51b60cbf204c82ad25c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e8acfc19b9ba88bfc7b53cba086bd8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfaa6b990612fc69d24306cc9669ca1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13be2ece12be990033a478e17af3cef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac6f08d961ab56e584b56f3fd067a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc7b52b1d74abc31a78f9671c60b339;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bc550e5ef5266cc38934b5b8a20de8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbad5c369b79b840af1a87d851ac6ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc1c1732c12ef2384c98a3a1b4aa90e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19703487eb0b9a3ca8153eee0221f33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18ccba70151eca2c253926dcfeef832;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hab76fa2d1489723d8d3ea0a8b06a54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h698ebddf33655569ec30060bd75663;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdc40266ed8a618241cb5ce8c7ce001;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12b3fe129eafa0603d1e39d3fc213e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197aca090be186dc48937b99d1f695c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5cf3fe29f23490f228cdbe265ae682;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8fe4d00191bc166af7c8e88e92a0c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c8a31eee4e6a60273d050cdde7016;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13d4b1eb739016f5481eb2171a9064;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd3cb2834d0c35ab7102ef5f7d83601;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdbe97e5d61123f043bacb06a9ba99e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10bdb941226dabae50107adf771404d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h96f057b2014836ad16680a1bd6a978;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'had40abb342adf399024cd2b5cbbfc2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b49d6712de0b6ed62cd49118bcaa2f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ddf3e247bb9cc61fd0cc5e2bbd159b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6841071b7bf59994760b8b5beb3a7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h25cc2739d17e6936aadf0ae42124bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h161ad1edca4a8e6743c8d4479bfffd7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13bd061b468bac0b58525515e9a2d3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec3ce27476e6b881cadedf91a7cd70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h73a371ec72bb41016d4b77d923d32d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14889c80512689f76f99776d51ee080;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1062c27fa35afefafd4853a4fcbbb43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1608b6943ce415edcf2286a47940df4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1373578315733f60f4735199d3be82c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb60f42a065fadc7ee9b7f8a6f106a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h143b44af6c69e2dc176f360fb757703;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1334bbfca7585fb06836f0db1f28414;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17ded616db4b88c4113a6825b771c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h126221c5f649d306041817f1251b35;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hadeb265e9be04a644f65aa655dc67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h181f2442db5ea99c32e5a1d0e1afb70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h940bb85aba6fd272add680b822446d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33e0c0d8ea0797a932324e66ad3c44;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a3227eae5ea0659c70b54d7d3649e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1879566320e659b331490e7f8e0eb22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18456351e2ce07be5b487ff783510e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1373fb45ce1c93fe33bc912f6d5a797;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4e8807d66a13499dccd6e298e0a12d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcc97b7d3d01313ff30d2d8e5fcae3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12594d24a45f1fa4f74c12669044693;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10bb2a06eaaded098d8f0b279ff26ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f4115d91e0d8b7a6b150357ccf16cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c8622538945c0a022ab45371d6e195;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3123a9c8e0035726e34b9305d380a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be7fe6c3cb8192c1b2e4281525806;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5cae57bc94584ba764e44af3a0257c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c29e9977e6375a40b5098411ffa3ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a813fc01d96a5cd1c3df038a097f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33661577adce8fde054a1d89e13d6a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8311bd4d7576de37a36a30586182f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha2dda3d2c5ec9a8544ecc88cd3b2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160dcf14b07c4de5ec20d25c334f792;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h143e65256e4cb729d1394f3f4274096;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7d0872bcfc86ce555a37ee00e4fb48;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec4ad0004d3f739e21dd0699de0076;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd8d98f704c72b4669a341a1e66ea80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11cc93a18b2360577d2b16de4c8d1e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e655ecaea95db090e7179512fee055;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8ec23f4d1f6b1d8c4e2b40579973e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4b481e4db9aa5956115c1500f642bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c50b4bc0d4ca0563ee0dc1927697c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159a01a61c8d2837d6f23f651b58c0c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10b66acadeee6d6ccbf3aaff58c1917;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h155e9e75b90ea9b68adb0b03d82d5d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cea2982b775bbc8f093da50a8c5165;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d574a549c278129c25a682f2356da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h644b4029960cf8b4f0c207b38f00ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hee9a5e1115e0e4244071a2a0e444a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce123d9e1829ced8f0f94039f3d4b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h628eeef1db42bb377ef3b4b8a04b5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a39ffed09173a75a6de162772b59d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h58db973426efe6eeea7be796f9ebe4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he6d888f8872545d83c877ad57aafdc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6bf3363866bb8978781dd032c9c81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f2bc6afbd096c5ce20f9e175112ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf2733bfbf73d6951dc4d6fd3f4bca6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bc67a11e27af70f0a6fdcc788923dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1717dab6f2a75317bfc6c5dba33d80a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19ca72ad3639a287cf2d6157283d03b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a6f4b7475f4ec2b0a580f7176d36d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16b7532c93b9abe01d168dc0ad5296c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h153e361566c98db247fc8d7a7e8e988;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h60b5865a7b604e687f74b4e9989602;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1625ecfc5ee1696fe8a1a5ce0d257b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d6f585fb738933618e69deaaeb2f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha7490cd57fb84377b683fdf617b3a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a213d3bb748add503379d89577e99f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc3b7261e9436a473a09c24f1bf602;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1521de7bca4d79b82f2b465d36a919c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a430fccb37ae8cedcb21587eeaa32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h22d4020f8d9b69a1bb804c8a3704bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3c00ab91adab027cec888872f48074;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aa04d8873e5c941e55b236bf8f7c24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f64bc7925b8a9566a295d555b5ff6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e158237826820f2a61d199496f881;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f0cbaa4c825aeabac5bc8a29bd23e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18ec73820a74a275af72b81d58002e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188d02e5c199d652621f2f1fac0b547;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1770f1d5f6ec5a5ecd691533eee07fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h40ef1611731000dbfcc36dddf184be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bde4065f45c97b5ec28dbc885c3dc1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hba2b43131767396f9b9e7418b00368;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d4d5aa9ff61f8bc6f77ad78fca4a4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hed6ad21d14898cfe5b052fa5813103;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3cea0f2e10aa3aeb808ae6d54a610d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13a0f5ed60a4efec3b41f521f0e0ee9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h144617484ba223c5bb35154b199ff2e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6c9c9f91f1214baacf28b9d0dac5b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h153e4471f7cc0e3d8e70967a9ac52f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd07139653ab6a1c090098053d95af7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5822a253c79eafda0e7df40fea03b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h946aaee962d5d6c60f2e2b10ffddbf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a49a78bd74e8a243f247519d32c295;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd9ac6004f02a25debddfac6efe9edf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17be7806414994066086b3b9fc2df5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1092800adf1eb3de02587d85f07e764;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5b5135f97354f523a6a316c692640c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a3f5c836ef9f02ecc899028efc2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h834a8ebb40d13a3394b371b2962f56;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf1ed684e451d5d8b226642df500665;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15145ed42ffe7497224f065a9e1e9e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he1db16d8b2c3236dc50f2c1318d7ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e081eb1eced58fbee16d3151d7debd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h80c606f6fcecac4d0dca06262ea157;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb0811028a8058127b3424a1ad65bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb5754aa8aa4bc9baaea0d1ff9e711b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb9b35ccfd2096f064c0e3d5335ce5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f3764946790263659d3d3f6c8dd184;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9ddf23da2e8ded54211566b8dcf0e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h765eb4b0db0d23264ff9d26e20d8a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16ac5f48816b95b1ba257b2154519d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h85cc08899fa15970b7bbbfafde26ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10303620d346867ea176b3564e7fba6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h32fbf8470b1c22e7713207a1c949a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10fcb260c883a0ad6f1b4dea65a9572;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf58da193f12bc162b74c4275f0f22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9f31b3a20175709daab98cec5eeded;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145aee8ad60e0d0f1e462558f29729f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcd7079e42be5f91378fba86767705d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7db7b26359af21daab5b28c4d7322f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a9f4b3afe01c92dd9bd3767e5fd94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5a66304c58bd240d073d0fc12ec42a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11a2288dc2195e2aacf272823ee38d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d24055e54ec08d98418cc12f7f58cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ca69984ca9b2fe1d9d09965b0ce4b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e44db99921e387af07eadd7a2a284;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c3ef619e8c24b2a029f0581d8cf994;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha3722bfb47da1dd110a52d24f7cc8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h55b89ff48204212c78b826501a81f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he049269f8f543c21a2f1f51fc3b0c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c907d086f21b2be78aaebfcd6499a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h194f3df0711ad6da24c91281e316efa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bf705f8fc401e36ad06a7896c68877;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a1336dfc67839e491fca9e32b40672;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he472b147660bf1e9a1f7529f4e670c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5a5ba44279f003fe7aa851d0b02b10;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h136bf584ac7658de7636fe11f1b06f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e8b27c12fae61bd0800a5ab93e270;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a17bdcadb67194226b50a380616fec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1036df70302d385209862c602c4b1c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a6379c88e2775d164289e902d1743e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9128e7e1581f0143e92145b81f1179;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc401b2eafa7a9ca1f0113b58e7874;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82ba7db193c2300354213ad769c47d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b9994935fc212c5b2cceed4254e6c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1016a0a49108c8fb3883e74401b0a90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h96378bbe17a9aa96675eb791db9654;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb898eabf6b93c6c98dd61765c538b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8f1d68e0f050650b7a5c4e9c890681;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2b10d1fec1b57136d481a3e5a9250;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11e8d6ca01c3347d4ef86e00f62de92;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h23bb01a0c5ff67a53267397f50b40d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8ce2c47c9671065e27adf48674b691;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9394acd9e379c3149271caabd3cc32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1826d6744b6e26e584ce8f87b6dabf0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c291d61443487dfcd165f4b10e6d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5f49a45cfb4303eebc17931e77851d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h420f415c2e181b9a3d6b9e7a3519a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a655151341b468b391f73f6571468;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1898b4dad5b5420b2e74fa1d22e42ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b06940ac1a589d67d5fd32b397c484;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18b4d8b317d6b108d7235aaf875836e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h119bb9d276f793dd4a3de7008d1a03a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1af0b9355cd075a2418eedf48975ee3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he7cd378d23fd51fac46809af2fdc0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h128c893de380792f8a761fec4140926;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6959e30e1e57e4ea0ced8e5803ca3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18455a403a814f8b01b4704413e8b35;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h176cd78d72a45f9a830364b8a839c5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa2985c9773e226699b185bc1fbc2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19895779c783c75e9efdae974601e37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h497bd977f1cc157ffcad05c8522cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c074034415ae60fac08c7bfdfdee73;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e50e3f1f21a8efa71fa94cfd7f79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd583db0652d7243ff55238673dec8d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fb13588db233697ed754bd7006268b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5617adfbcace80dc1e672b2cf02b9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dc715c14f275f50dba441cc410d958;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd25567650396782c10060820c965c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11b1dacf2efb06aaa559e19ae475be7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h30409fae45661b213ee418d21984ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fce5dcc0830ca8554f723446d7b34d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5ced8e3318a7cf01eef8c136ec1dae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c106121070b1652ac6ff54aab70541;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c3f97739956840d31d4aea6b9e998;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he6172b82050c0a4d16459d239b4233;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfbd74ee8f4afac995fe49b530a8448;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14352fe3a1320b1e967515f57df9ee3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h83172f9821469cb8c38c6fe8872323;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf2c6dd846556918e2b3d14062e8e56;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a42682ab60443d3ca2c25f8855b8d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11b8793f9fef52f941b3268dead228a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10d042f78c1243e9f1edd2cda2414e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fba3348147ff68bec8ea64ee20ac3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c6d41cb4e8c2b7ea8eec7d10722e88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h193f704fd9491f8f6f90b4986f4f40a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43122c7db4fa90919cc0cd6aec22e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1833d07e00aee8904a639861898a0e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7a2d4dfdb704472dc43ebe7d019be1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb9c586653b917eec3ef285a10fda8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba3df208403c203cc07d66268510dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb408f82d53e9af900b3f83e3a38ff6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18fd60cdfb7f5bb562b0b64ff34c2d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1209821dfed75f4fd8907ff42ed10f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb04b6a22fde78971ca516f66923c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1053330e436b3329eb9d1808eee2f6a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he6bde766b207c198b9a20a14a1e4ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c43d40fd889e5c1213c41dc35b0aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h77f77ccde9090f64c711a6ad2ef349;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e346064e1baa2b8066e421bc8035e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec6ce6d74028dc3cfd05f081eada4d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10dfdd628c066a04244926dc86c1b90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f5e42692f12b009a102b4daabc0f17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfd1c3d2c2a2d33e111aeea9ef35505;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h45f2d981f3f34ef150c0e0f4ba036b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac1c3116fdce81a7f915177817ee79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2bfd723d58f202ffdbbb1713e7f3b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h78fe02c0454314110e9ce1bd1b971d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h153fb9c58a639da2bcc4b80e129bd24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb6abe06db05e7cfe4c5224e06f1f48;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfbec1888e68ec7743466311887eff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hecd177ef274450d3cad8b7cea3ccf5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a4f40456f2451e8dab7a57338b8acf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h851948f79e95ab6b82be4ac8cad9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd00abc297b598198d802caf833494d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11007f327893dec0767e8cca24ee42b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188777c0193d13cd37810f32a3949f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h156d65f681088790862301fb8fd7847;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha0f0e49e3c918f605f21b791a502c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h59ff1a1b5589f12a91321fb0cfe1ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4c0badb964e5d1bd467ee39d4e83f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h25a7772e3cad285b64611aba82c6c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f4f210146fce19ff6c6205512dcca8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2d230476ea25976a88d84079290c09;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hecb2d8a555b97d4fa82eac0ed47ce7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fd49d24505c819292f5fbf81cc66b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14fd0d0095969792523765a348b0f56;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6003bbe839e32f522974b8ea047898;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6373db66cdbcf1ef7a42f69f9da514;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h189428b5a3fd8c1c8711083a0a8eb6e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e632a86157b4300bf80919a84a1db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf173dca3a495a3eae02b481619b061;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he8dde9eb82078e4c9b0eea8de5745d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h64df4066cb698583d2d43478f10d83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14b847141f44adb31cb61365034cb5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188dfb019d07bb4379812d5d00542b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h441f8bce9afe8abdaaeea7d00aed8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h563e1886d217eedb3b3c60b8b22d26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h41af3fff5521967aa38d4a05e57949;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc1eb708c632f97b6f19df72f2074ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1065010e96607f52494373a813d325b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdf88180dc77263d9122f0805f61ba8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9b4a0dfdce5e5e53d080920a775ec9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc9946a582c2a429def3971d8ae7669;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f4ff805679817e5f795f0843f77c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h96e4816b227d45f8de2ab07919c518;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cf42bdb8d783e8ef9e186a34f41e2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7b7a32fc9b31c5408d560e30a7e8cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h53362b6f20687d953137703d8283f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h91ed428f0e71a85780e5a1befc5d19;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha5032bbb135e6f6ed80994d9256cb4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf3ed30ab0a0f27f8d7abe277f0d2ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11621606d6662b47a86863398496808;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h557e2815eabacc3d5ca1f11524445;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h72bb31ab151c660db9a3612a10d646;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd7fe4220f3690dd2c253d5dd479d10;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c3d332cfd5540e4edbb50c8ee933fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1176dc5863cb07c09d972cf5b1e8693;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e77e8abd57734f79eea007f7c67eda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18df89364f9024f8fe21650dfd01322;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h53e0c922edac28b68a6c3d62163e72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he8f54ce735bb5dab511fccfbedd819;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5d8a3759b4914e79676aac0a08954;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18dc6809f3232ae83b4faad6c6c8211;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf9c6c24f44887da5ed25a87ced311e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17fbb6d8b5fc4d2445d01f72f41f8e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b8b94999ecede54f4205f732902d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf313ecf7d46a88d484307923a42e3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfc67a7fe7a38222bdf2434572edf50;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha3edfa02993eb06cd802bfbb83ce2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'had01dbbb38062a48f714a55c9321ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13471838e159b1326c4465eaedb513f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f0f3d7483f86fedc1ac7cd670876b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h105e0943adb1985b714bf96d889e22f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cdc574924056c1225c0e11a5b5bada;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c7c0b57f74a3d8cea70f84f3aa5910;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6b98cbfa83c1eef64891b7287bc2dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h85120251aba33cd4b26307fcacd6a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15ee34b332f455a560ccce5dba1a1e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e88848be4b065fd644e5bf5ad8475e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2206c8fe5fc0b1442de65623460ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fe0832ea96da57dea6d60ad4e1c392;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h189d63ef31748db8e01b955a86abf2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd7ecd7906ab08e9c6462028df2f79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f509ab79493051f50d02c5ed61438;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc76c8b82c84ec846654bcb7965bc8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a697cb5e29ad108dc227e30356bbbf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe6870283af63d8bd06d6535a35333;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1943aa0c2a7c826572272a9afdc602d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13da814a3816f4f002bf4848049d125;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ff43d3f15b26f74137b8b0dd030605;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h48412352ff0bdd94658d402df751b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a23c254576cdb4855cbfae53d79c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15efc8496a4d1d0e8cfef9d58f3caf6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8f4327b43990ad742d4024cb82a24b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h402b8785d89d16aa5cb1801296930a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1316ee79868471384fdd6ca38655aa8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18236fe878a7db4ad480aa8dd2f1f93;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h308249b33c9ee7b3deaa559f5cd12a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he966a6386308586da23e49b72f4c20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e0767114723ecd708cf3dd3beb3581;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12b9fd1bc03e77ed5d33084d19b05dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8737c1ae624f6228aa562f7cc12530;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbecac344ee9b2445c81147994e373;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43335f5378b5b3ba8842db62a6f01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h752dd591f9e9e37672cfa46896a01a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1013c57e28a98d5ea0a807a38493a8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12af8b2c798c75d495e16e054230841;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6bf0376e9c583c8cd33522532c44;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h546d421df09017a34bd4880ca14495;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h242a841b5033f3e557f5b0197866c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he03fad1ef2b69e4b898138755f912b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ae419daf685743a54ab7084c6e85a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha8d632c3f7fe1014bf89261f9c100b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h95cbe208b5b696caa09585ee226f03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1151fbe4ee9c6fa840d7698443d66ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h120af81df801bed59135755f27ba563;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1715fc39fb31eccf358460402a27c87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c20b2a1e1e97ebe7746a39503066f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h173b36cb6f5210925e0e323487dd80d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd48a23c7c4056698f29ef904b7b6af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h98bc0fa8ebf4a5cf5ae1683a0afddb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdc61a1a28f5c71f700cc32d85ea659;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5b9694c62d7a34f71b2642e47e62fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f61d2e59496ee550ae748396af477;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1422622c7a54474a6e76ef4ac545dd3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1af2b768bb5c9ec530ad64ccf0dd06f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha50efca855fca1e4405df93f036f64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h66ca215bf71a107baa5c55e2073df8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1108183898d5bd608c203e8fc0ce286;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f10ce3295271b8a1afd79f8ae516f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cda961805495ebd621dc74bfcefd62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc75812319b71265fbe261ae7d4cfeb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e215ed1505c5bb6b4185d178968d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ed00d0f85c283d1f7bd360473653f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc4e25756a6646be970f1105a64d8b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9502695408d916ebe49031dc8bc44e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfbf3bfd28bacaa72c64141e2e79ed5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2b129d63ce121b103dde6a59ad36e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43309b83626da7f726d3e5e9b11340;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfa9e6d4ea46bee59c173759a309955;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b0996a4820772c2e276b0d150ae400;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h135d7497fb90222a2b5251613f3485d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h191109084cedf91b9dac7aa920be548;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16a602891d4333f397bf35946acf362;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1840c9c5347f0ac9fa71523900b34b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h386b0cbe422b4c65a782c9a3529bc9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14393868aad8d0405060cce6c0ac535;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f377c6b3e019497c5b2670bdcb2648;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba81841a7936bbf7f238b50b35cfe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h961408143ac7073ef4d6a4eef2b683;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1540c94e6e7332bd985b24e0b0645e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h78134ceec15e11eeeb6f34f39af30b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bf79509d5c8cdaff53cc94f150a1ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h194a3416b5cbd7682553e507c66093d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18516a84dba80eb9e86417d64845d14;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h629a94f843f6721882e059acb3fa1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1279197c2f4dec92e3f484f7a69bb2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h134ebe9da745a2537debe3a42eff9b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12e75c66fcf6ebf59d7e822a829c05f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bcc7565a4a9301fcd1cc9a28720728;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17da968c44cb72947d5005913ced21d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a702396428e1cd7ea42070eada52d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b691edbb308ef0270d77390cfd24d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16e417427ef4bc50221530c4bc3a6c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10179e53dc9e89cd44fb96e1ae37328;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c0b938a7f25feaa819aea7e62b8bc1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b272fef99d964cdb9e02d7b21827d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbbd8f48462c4c6d992fb727984e145;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1786975bd95e3610613f1db3c0ce99d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h76d17c3df596e81ef28671a6e24cae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14ae4c4809044328891abb4a4f8a732;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd8a108afcfa5a34db892169ad3f7ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16add2e9481f74e5b8c761630707864;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7db539b736b75ca277bd601598039;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16c5f96fd25a6f22e1dfe6a991e9310;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4e0e910e0059d1ad7d280d5e1ae98;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d3499f9ba471aa5e3d4d11556a14a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12e6adafdf5f54c92d8c0dc1fbfcbc6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hef2f33c3608321b843cec676b68443;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c3e001d0be058bc282d97e05874f22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d3bbf55b1a7bc63f729aab367ac57;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h80fe032cd0796458e22ed15ec9bbed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h841c461d2633c5b2e7bc3fb0814539;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h56bc807eec935b9e1c3d22bdad3e31;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1050924d9078d2e51c54598cdb696e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b5f44aaa3d3344d053fe927c98b49;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdea156f68cc746091c754215d46715;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h80266c2d7638b3776302d777e3caa7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h202153822c1cd576a3051bf6e2962e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b9ae093866d3c13aeaca9fa825ba42;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb0ba9c25460d0e1cabeeb8270ee4d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h56d90cbb8f015fc6d0553ee315e65a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7e0ddc95f40c167672cb598589430;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h55833d80c0048034ebb63c4b48c859;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1da5b1a310afd903627a9171c59f24d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h57a31b64d4c0def094f581719e724d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ff5af513dfd1ba8e86230123f7a8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157cb4dd41c28764a39cd67a32d1b28;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6b05e4568c673201f5b0f056d99d15;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be1a06e708662e487f5f2fbe921f9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fb7da59876c1c3beea21a2e7c55024;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c159f9f69dee6b50b9145c56fe84e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c408bf500c46b428adb3677a524360;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c34edb80fde87a23899e961dd9b84;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18908b963ead138729f3a7d51c049bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a9ea033a0f3e6c5fe4513eadd980b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha1e2f5f26d052d9fc182e543c97b09;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fb810991c9d818c7601b5281abf246;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1092df0a1d258f8a1a8f37977659f7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b831fcae4fabbe7851626698a7726e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13e0334d348450f42d7c70dbbac2b91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha278dd0d1d4e0ab4a388d53156fbaa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5ac737d797fb368e7bb1d8622e8e9f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6470a91c176d8acf98096c5020cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf45891342a4157ac1d0b9fb83f1dad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d0780b5f8dbafdf7877d35901c28fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a14b8a786c54edfbac3910de4fc13;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc1ff65ae5d373362dadaf0b63bf3c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he8eaeba10feb8bde5468d5ac173b87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a1d38be14a2287a4c7b85271bf3d80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111a236966bbb46587a741d46c5a557;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb9535181b296b10c40c831ff17aafb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2c0782d89b658fffb1cd26f47d60f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9282a3f857c8abaf5b954a9e73647;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h115e5ec1e242c057de81f521b4a4ed6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1cddc386a098d4b0972ebc3cc00fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1de2fa88663923cebc6979a20b8ff14;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h58e34fc6f43eeffe762b985ffc6dee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h105377645acd3601a88acc55f4ce7d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he876f5ed35a0c80139917bc77ee2cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h357578d65aa96e9183ec8aa250d6eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h180fc03def5782e49c9ad531ce4c1ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13075dc331975f733b95f84497eefc4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1368d269c0e94bd72e933e2d54ac2d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10b4f639ea94268db6b4e02abbc22a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f44402ce734973387943e6db2b960a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6b6cd20045979dd95dc6c0104362f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f3b12064aedcaecfa3fd82109cb3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fabe5f03c309fd1438a9cc147c1315;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd4a68f84f8286b8722b205dc9b269d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h872769d36c69c1d8fd20b325806564;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a8982fd507da64427aa540a873716;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h74ec2e06810d7ad1d00d71c5ade2cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1664b1a5fdd1b796d46275bcb8c063b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h76c3b77fc347b3904aa0045b25fc8d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h117cbba562e67e89b74687aa124db0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h110985a74a2044b6043c8217505ca76;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h30e4c8b36bc064ba7ab4102f26ecc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16869f5e61265a65569e4d9f62f7a6d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb3226ea6e5c0f8c6eaeaf9777af217;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c3b3cc53e1cd505b022ad60102f7ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c46c61e7ca281cc6cf3dfeb77b581;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h178126b330545084b7e58ce8af7a8d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha5c4e3588105724d0d5e80893c8e2e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1740c2823f4d9ffaa4a162e60e51df0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hecc84558f9b71dc06de6958aaac7ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h186a0c4f0c76bc5601b15915ad20ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h527b81004c9559ac0d026ea826fc5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b9caae3fd2dc7343e9989c29b12c1a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ccc52b9e4ce6a7a61c3de99fc50e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160903c0165b352433ab5f9938e174b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7347cc17e6ec531fa2526b9d7cb959;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15c62f73126e843c54e2fd59b4dc3e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1210fbd7e07cc1a564e249c2a60da9f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e917b6ab9340b76313b156a2141cf0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f1b88c709eaa657f0dc8288618d894;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h565f4aab9f19c75bd2d0049ef6ff22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd31b211fd05f19580d2923dad1ebd1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ca218b62a83b8547261580786534e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce90887017f2b3f09f28cfbab65ec4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha0ed39c24dad4e33d49f92c9bcec5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb136911830cb18e0b7bce43a2edc3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc522ab4b95fd8579ade83b17462b1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h724e37ad67118ee64c33cbf3c75aba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc40d0f7e2a9a4daa8a71bd6f0040d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb883803620d23dd54146f0e2fcbbcc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h97ff23f8f08262c0a17d3043d7230d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h248703e8ff5ae9a9ddf7031cabd1bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1167ad6b0f51508a884d0b4afa7aac7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e1f9bebc79ca19b39bc8462f663b80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f0ae979a485e45b1c447088aa43dcc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9dc6d5a3dbe3462502f7d06ef3d55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4c057d615cf75b43d4abf8a193a2af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6cefe0e3f37a1c5120ef72a8822278;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a6c7f8b5078b28fe4e00211cf98c5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1613beeec72769ed61fc0601c58aa59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5135ad2832bf9e3a32cb804f7669a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c324792d0bb156451f07515e2b1a73;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17fa46a56d88ddcecfd411354ddeaa4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc018623b483011ff5de9b0ef93290d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7f83c14dc421c8e3ea212f879d1666;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12891a9d0647bcff60f377c71b2dd6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19c89bb193bdd01f16b78671e6c6d6c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h131e9d4cd688867a59a453f710e2abb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h353ad35cbe7920bc54dd6006215edd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188b09c0e09ba99ed9911dc6a568e5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h836e3eec89dc30e6f0dfee04fa657f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1169cdcd736954a9a790027b7f3ec95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb262cac2d7bf564d259f3b396a3b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc94960db38d00aabe0d5928fe43b2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h31fa67ecfd2000f9fa01c4ecdadd51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf7c53055b206cae9d08551e25b2ba1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h87311fddb91479aa990321371a46bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12ad2954440be2e706f50ec97521b69;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d9d7c65bab2487a9506bf34f511b15;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hffd4c7907445354757c1d19553031c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124a72c39fdf97c072f383aef6e517c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc83dd29e55fd18a68940f685bee43e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4666b7f3e1cb4fdccc7f47d27ca1c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h45fe53e0890938b3333978e35d067f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1acdec6ebb16595cf54820153acf91c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h147c1a5f7ee2047eebd9d90b54f2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c4671afe48d6301746e997a8c4231;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h23ae56b76af260dfb8c428d3138861;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a982e80a1213c6cedfa1fe3261d51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1025a45e09992b908cfee59e5c0bff7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f76658de00bff625f1cf071b8e302;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h31a80f35d118527fd9455c139bac24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5704ad5455f99dd9e88180b9786777;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18002a2020b9c77be5e9b9dfbc077c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15de042afaad222d48f9ec2d10f5eec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13aea1ef376d2b06b003580e44e8828;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h136d2ba4e94f151960a0225de0b5735;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d732ec1d7cf02e15d1ce2c30990e45;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'had981cceab97b6d05ad412d90868c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa2040e6704f7e2b7a563e83e866ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h225205d94d0240fa6aa8e3bf8fdab5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd191248356d4428a7c6d88fd5dd9a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d3ecc831d31b6c73d2ca1a9c81cad0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h231c144dd261179248035701848f22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h156b4b38018e882bfbdc8c7bf2354db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h48f1ec688be84b012360fa73d6501b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hddacbb3aa6e4b6a032f2d0c1646cdd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h28cb33fef6096d8a11b1c602177c88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb0a0a45ebec30f973f7012baae70ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17ee84d77500ce6da53254efd303934;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd96a8dee2fd86e5a9115d59dfc3bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e518e7b85f946d474ef048cf7e5db9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7818202de94a950a47f092f90ee89;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd69f43e9d54fc80f8a42670e1ecd3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fe644f417f0a63ebe2883edb15934;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16238188edcba0ea941d61b7149fe68;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h992ed873990a744e442c8e2dd2025f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4b4086241edf071f6624ca48efdee7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf5f6a037bb524e1631f0d38a6fb0ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cb94edf91e4620da8e9daf4a0155af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h42748953907e5795c9ae4f8e25fb21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1befae0a518eaf2245f9d0922697415;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h114e8f088dd96beefab759ca652be6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe8d7407bb4582ae405f1831447ae3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h108ff8da2d2000ff32869f3adbff77;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he3df0d92a5e0bdd3378e2639095590;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h179a59c98837bfc9a9cb4d018cfad51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc7688610d309fc223002523a1d85c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hadc1abcaf822d9c65e163420e61820;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cd1e5c5829535f1e0b9c5c1fcdbc2e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hded88f38745af0317d48623108521b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h152a3ef3156fff86d217f7a3e03cbc1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5978f00d78d5b289ce8a6ad35c6c5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d104d58da6cded8fc05508be36b591;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1101eabf6b374694f8a88953216879;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d981b58acb7832d9b8832980b2a782;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha4dfebb0c5b65f41cf231b46e868ba;
        #1
        $finish();
    end
endmodule
