module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [16:0] src18;
    reg [15:0] src19;
    reg [14:0] src20;
    reg [13:0] src21;
    reg [12:0] src22;
    reg [11:0] src23;
    reg [10:0] src24;
    reg [9:0] src25;
    reg [8:0] src26;
    reg [7:0] src27;
    reg [6:0] src28;
    reg [5:0] src29;
    reg [4:0] src30;
    reg [3:0] src31;
    reg [2:0] src32;
    reg [1:0] src33;
    reg [0:0] src34;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [35:0] srcsum;
    wire [35:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3])<<31) + ((src32[0] + src32[1] + src32[2])<<32) + ((src33[0] + src33[1])<<33) + ((src34[0])<<34);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb91d9c64673f69f7ef6a7532dc9feb4006d833086f38d35c47ed661bb4ee29a813c0a0d0f3e686a1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9ed5d060b7e66608915b636931885ccd64221ac210881dc28254d0b788b4ebe828b5c241744bb108;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf6a53170c5b0a8dc6f9c412d5ccd53a55c4643a280dc2481db39fac69d75de062379f36e7bebe34f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72f78e3869640ab1e138ee893f2902b64f0662d1fdf011553555f05493a32d62b3e2208315de75e66;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56909d7d35843e6d48be773de4c308c76a0a2fac1eead5b66939f15740e706ad800f854c32e403a2e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdf99162d5b8786e1ff6cc97b01151c71f55d04f8b67c419f2a16dca4f04da4f6d60be0349f879872e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98083c13afa89949b2df3268f0314849c54e38994824d07ff1dabef922220a7f26bff14634b049118;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e42af54a894d6734f5c047183f4b96f829c2c34270ab89e60df9a45e9bb2db9896303787361cfbc2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e3ea7d5a97470fb1bea227878290a69932eb3c97839fc410c67638d9600996b287943fc8bfd9c5c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38cc63ad844146ec0bfb80741ae9ee72e89e4c2965a2f4f1b17417220aafdf0b447da514bfd6278e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h204c4ad29f11760c10ae37fdf1a3ee29a6308afbd9be2014390a81fc06eb396da1a93618b890386c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9ea463c46946bd09e1aee2fcf13b1776d1e62b69c28a1e218bd3549fb1e60c77f691483f457b620f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h351a89f64bf1ff925c2a6ce2120448d8146cc7b95375e7071222fe2508fd89e0b9c6e3c968ad73229;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d30f3e3de1c99be69593afd65b3c35e4605a773ad4ff9e634215c87a04f70b951ad8a7f0254c9649;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd15e62e90183bcabda8e9e5aba0f6a58ebca444856f53c1a84b6a29cc68f8d2b52324d7c1c492cf71;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hacf6fdedeb3fd30d298f01c3db306bbe095126c489f5afdd6cab68064fca5a7e6e48eb3503f81f269;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd55de37d876d9546fdae14c36236196fdf574e7331e4493ba437df09fcfb86f1715efb8789d9b0226;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d7d8630cfb184dc006f71dfea0071f254d78ea21eaf86672c99745863b8a246817e76896efa17a07;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89b968cdeb2e6cfdee22e8a33e2c17dc669a640f33e4f9e2d2583736698e1b9a5f13c05728be2fb29;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60872d969e1eed9dfbd92f583920acc726a4211e762a3425fd5cb4b059a26add832e45543c8a32d6d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd48b4caa873970e1d9cab6a03ada23fd7acf31cd675f557bd9e5198fe455f17dd735a5c1797335866;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce577a97003a84075b70dfff85f7607d25e2aaa1ba3e3cc28da5d7e3b2187ed60fc36ba4ab0b49a59;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h979f8ce5140fec73beb37d7a90eb9e7e44d7a44cc0c0ff681cf5d6588dad8a6bd419b2fc7a4a966b1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5a8a615f2ae0ba6b0bda333ff7d6c6b6b6ea4f89b9cd54a3086b75468a217ade54e008e14a418a53;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4447545116f4efc9ecf873fbf67b0c779e3d567eab1ad14a3e0d4eeeb4f721859212dec79d7a680e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28e5fdf938f1340531302b891daba6bf78f54d2ae1def7a67103ac0354f2eb7949f92b6481a2d4a4a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95da97a723bb3a10a877e3875ea57aab216203430288ac3636a76732a5621af1724e9429a85ee20c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6be0fcd69e2db3d92204f64a62de343398e4ce32c1d5344f3b3eef50eec7ecfa68f18cf8462b3014f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h430760880e8ac6c8c3857214c33979152f5e8c5a8e37deedeaeae1e6d9701ce4698993c244a1fb3cc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51d2cbcb54fc2a1c62702e89003a4e01bcf8fa50594b840bb7798e9b82cb3bd9ae064d539ec2495f9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c3f64bd4ecb5c1eda7d31b225780c4474c14d912c30a602b83c02d395b26fd1698cbe0e2cba336df;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d031f959d9d02ab6e51617acd7866634d93f9543e5138136c8bb06b0b69bbff989f841a4d70d68bf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha63f6d861891682c23b29cf4cfb4a83eec3f51c97760d51bb88914e058af6e2717c69600ffaf70b93;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h304c3cb2c761166bd9860f9d0199742953c4616c998fe7fcf8ada5c88d5621cddbaa5f876c264b6ac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f59e11dce47c1a74f3e51692cf1df7800e47aa267b6e5a95b5c30a6a3354eaadfcde72454735eced;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc7f1c8e46dc37f01a90e1d8a52500c3f013761895fbe5a231efcc9753d2383d0a83a1d1d6fa8c989;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h670131cda5a482ac61f845e3565e3f88af0caecff01d2d7b37501ea22b2bcf960c3b11f7f8de57033;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2729f6086f3121446b95770d255586190530b05a60bdbe60bbaff715773d400085b9d99e817cacbf5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5a90ae86f6f64d6453fc229ab0fe7ceb05ba2dfe6bde0310e06adfc0ca37955b5cf017965f9e160e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84e918e838ef82af230e914817b0c83bf137f1bda62e50f6cf80421cac4b589ca6626290581fd679d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92bcfe7b8e89112f6465d5a4a91266c9599b29c2b6c2c1f28898bd91906a48532705738d8aad24e5b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37058bf2445361c858c76551efc219be32f0f0fe0ce899a7e14f76737351b4563603b4a5e9cc6bc09;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc480a8c6739449749a2fdde926a453a7850c45e94f8eb119960f3f395beacd4f06a1b140497134dea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4cd94c318f0f466d486d7c951ea6bc347e685bd7c85888028f2c98ef444554ad2f1e39d24b6cdcd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfcdae0894c502ab3777c8502e61c5c25e7bafd1c86165321c812ccceeeb044309a824dc6dfa3076ab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd66a59ddf10834acae4e58097e50305dee10ed661227c31da2ff04a00dbe7e12ad0d96936f4e20273;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb42da477323563b6acd173207acb21d297072a78f5db9010040fbcffe10f4ea0fc5bae06515a925a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd23c93a484b235653a5a8b880306bf2123b27c01e1b2bf4704abb1d43e66a622bc3c0f38625e574a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15bab80998e1cdd562fa5fd46701bf805f2f3801d8e2976d5792538cbaaa5eb898967b822e2452929;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4bd7b777ea759bbaa04771cb6bcb7de5efb0871b28d7856fc8e072f330d255f1ba6b55fc46fe9a46;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h274d0620565635d4d64fcd7c2a78300c4ae951a8bf2ef537a23400431bd318746003ccfdf1f2b326b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66f5a64a73f1c01a3dcb56b665ecfc2ea0231ba749081cd9bb132f9109125476f5b6c92bcd4e6013d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h372bee32c926e491155a901f130b9fc840bcfeef00f9731da580f12e6e148ff4da2b38c30849b81f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb93c8a1fb08ea8180742394c965df8ed61007f10f2024a2f62660a007d6ecadd912f5938688f8e272;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40322008eb439b4578584d00a97ee986035087272bc429be46fc037662a8caac4b7a39ef38d7f4cf2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c7ae433c676ac4ff682adba90a13c8493f8e3dbe8d9baafd62007687d64ba7b0aa80c848d65c1c25;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4621ba5ab6d7e2742bb231dc5f75009f86aed1bbe9e877bb48d257b0be3a466a4c8bd8b55ccf3b63;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfd1e21f17c879c8299f6cc433d508cb30694649c64b10f7d1d9e9e12b9590df9cda7de7eb47051e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c15e9cb8b3378a86cb9b1f2ea182f2490247ea2be2b5f0a5265b7a1cca18a04dda49468ad00a250c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfb1bad1cd8fccd5ad04938dd4b1feb15b1b1e7b54d0a7868e14c9628c6f9b05c4218024a556ab524;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73336fc2a831c830d01c590d2f696db504c7659c00e8ce96c641ce87a23af99e0bbeb42efa9d56664;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h792b29cafd955fab3ebf8ac39fc5af262eaa37658fc2f9c5637c3f6f3f0406ac165e1aa5035fa2d9c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda62ab0bbffd285893d8a48326b97cc7d97520476984b5cbda1579b1b09d36f15c29c5126d65a3b14;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2019b141ec643bc4deda2d64925ad82227e116511a9c66bd3dfe480994c5a3637aade04f6dc868e1a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4975f427bcf442a2dc6e92a9add5bb1053c5a436ecee2254649427b96025475d9e1683b768489bfb4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7161a1c2b98fd0a36a17cdf5f4a270704445c8cd277bead3dc6da02e20dc14af181ced246514e3e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hceb3500606ee0cb43b6d51ae2b80e4948f3f02e9e9c47cd7e182e4383d151433cc315698dc645312c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h844833fbcbc8d41336cfad567738e0d60d48bc88230276d719df663c73b47c176f13f4ed6830b85ab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29704f532b86591ab4ee9f8858f989965a2f07683d6efa04ebc1c9c659e0982627904702f34cdb0bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h293e7e396040d45a0e96d64dbb8e5c1a5ab30aa146ced2c4c4c4c17fe0cf51dfc057df8bca26de86c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8cdd7258def368740b12056e58745d29ace8165c347bf2a5982eab37583e7dbd2dcbb905b548b855d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h494c5440c94677596e7e4be550c71f2ce45692780be0314abf2c1abc109c03be306a53902bddec76f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf34d4ecb1d45cd51ce3bc4e4f79e264f2623ef7b5bd647de73b0ad56b17d476b74342b6405f77d97b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71976ed7d430cdda69ccb6e65430e8c1ff64bdfdba6c47583df24fa73e94467b6b48c42549f48f96d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c6ce34e0b859856b0566d1cc66eee487f0b36ecb03a32a7ab2750bb0e7ef4bccc26ee0b9f92a73d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f23ef188bf78776d47f271a48b3a9c01bb5aa6d38e1bcd8f32e1761cf04b7483aa334935696858e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5da7e59cfdc1bc5bb675a339390e4b70a9894bfaac9c439833d94a917629dc358fbbaf785a09b1fcc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h887e8ca4e15151c03d0192fe1a3a76a7340140141c8d4a61dc512479154c43a6156964b5c992146ac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd17f8d1a7609af60aa4cd008199a261cbd8e49a153f601c7f52d66cd3dc74e4c8cb4f1d064c0c633c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0a156c4f54438f57b6dc35242c0208c57e5713cd1f2c448651fe9bcf9c7e604522794e390fe5ff77;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a25d8aec8dcfb2945969283b0c2f3127272e2e68a70460917fb2e19d8670bae3a9a1578bc274f5f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h700aa0b7ec1257a261c44eba95a0eb4a1bb3fbb26a1008f757cb448a8f82756d53894b445303eaa1e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8484d5b5caa29ca323e77d5213ff112c662dc6dd9210517e604fa04104e3355477c2e11478fadda19;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde3814ea013f10f4af2139d6e61eb806ab2bd61ced6a26f618ed591c261c203e135099a93b4f16f51;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6ff5fd01af3ab04d27ff31cb53bfb3d721e78579c84094434b1b69f0edeebdd7dde6b6f5dad2e125;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h536aea7e2e0c42748f1d5e8cd1bacb3d96851494ff705757d9ead0759d4c98a7d062763ec19a5b8c8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habf196a09360ffd71a52e494d6136e548cdb0bb737e3a921d65638975af46369060f69c02535da7ba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2d2cfe57a61dc0b705d472f8dc159bbec7f269c5921d7c088f25eb0d7e0eef2c8884557b0ec1c0773;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd53ce2ea5c89432812396a36a58ae42b349f03da1e165db9c312c4c8e26eac6739c2faf353caa16b7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd06c4cb28837606ea295215ab403ec7e1e910f3e421ee2bd0441aeb7481d266cdfb02eb664884407;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc0dc4c2f198268bba6f6b64f2bd446ee4d9df9c94c5a5ae9adf488860240751162171155b83db7ea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4386eab654e2b1984a1ea80dc9b0f4ffa010cdf30a7875af7770cd9af0615a95baa7c32b2c2066777;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h416c07ee5c9e4e383a0df4a7dda95923ee1c27f651f99b63ea294f0bc2de227c83e5084eaeb1619fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d4661272b5bf82afd950d8192182a073bf40517115486022f52471478d0f2c16670f6f21310043f9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78681c3e410929d4ae9d4dd4afbd7ae443cfbbbcd627e89c6c8f94bd7972df06ee90da2d3c5ef131f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ae7838337ae4f405cca9e9876c21056ab8f2236a174a1c9500eda2203f16d17ebeffdca39f634af7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95e15383cac3509a4951c9f97b67e83d68d8637d44eb67fa5b2dfb946c76d82ddb038a72c10025572;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29a9352d3a9c74898bdaf52f817ca8878640d14eb129ba0a61ef3d6eecc720f875d672219b7134dd7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d9da3c70af3c53763a6bd0351ed92bd6bc3be0db5ab0de80c8a9da8a11c14c6bdb0678e39936242c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd106dcdf2892a5cd27fd29d8b256b86e02a5163cdee707c8c8200cf8f208c1a1ae82aa2675e08dff2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68b3579bed83cceafcb5aa6437a36d8ad76a8bc8e83fb8685c446478f84eefeeca006349c3c5c7752;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50b4994dfb367523cf1c1422f914472f45a51a45b8cb6a071ebe686f44bd02daae292cc193f408776;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4e19d8e0d8ef771e225e10946abb6f9ef6bb268a48ed931995d7d41a83b294b4a2395d53eb0c900b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c92c51b760cd58293375b1988256c7966779e0c47670f8be12bca5e7cc1bdd7ecc486052bb55b7c6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd32ff39c5536a81cb6246fcf8d0bec87010e3f94dd5cd6c48eeff508471983694a70a6c48ef817f3e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f9bdf8e1abe7f523109400655f8485d3559b0770a0b704d8855f54900a8ab4e845b31315beb2f90c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha343358a307d6b5fd9a803db6740f4f29a6260cd52c49bc7b4f141f27a0717799c6ed9ddd034f6cc1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae3e4c286988861df9e74f3494235a658cacdc15fc61d956c82a74abf254710d49cf9aec3717a7e20;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2629b97985664e3b6148be548d1714dce217bc5bd93f8f84563041bdc555815f30a84846420048077;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e89c4a02ac878195750d2f1e4baefff8ca5d797a1f5c38103f7404b0162d10aa6352523f2b99e921;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed16be85faecc8299a6ca3274a6b58173b3050017e54146ee9f695ae0795ba40456bca26bc99eb131;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7298b5c6122177b3de765de82a49ad63d3d764607a83f6685991c23578d716002dcb517fd6bc4bf0f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9661d496d5223557a23f4aa6287f4fc2e0c2615103cf0bb37493cec324d3e80a881936e93aac411e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a3ea56fe536038c4b08fcb3bb62d2d8c4ed42f637ef784cc2a3fafee0c45d2874672a3446ae3ba41;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h724f9b4651aff6d47e42cb0e0af0a251f7e824588c55cabbf9911f753446e0e9f5409044c522bf726;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f8a97be9a26309d4befe16a8cab89e8cbc2b70477d5960038f573b06787b34f894d83d06822ff2d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbcde96bbf07df697a035f87ad25a6a6c708da9fe96b7a26af2403a46b71d7afc9f2b90593fbd9c19;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7c12930e8d840f1694c97840fc37c69e1db6d98328bd647e1771a43862087482f67de2c947b879d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd13c31f84b540f7395b8e211d98e01768c649b67a7334378cd3ceff4e0e21003590a33b85f4bf990;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha54029047b86efee0245ae194fcf58b21034a349aae71fdf813327ef26849cf7b70167d3a07914cf5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae93df1f68aa8ed0d43e900d68fd9850d521b5f3c1579145b3d98f5276a8e2b2b0b5bd5796837f0da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd0d5a15d1d5727f8816488dab6d66eddcbe13cd492bb78c9f47645ee245500178c637d845da0829a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea574002bf559525c2a82021b013f77f02d97e2d8aeab5ea8fd8a9b478aa8be62a9e92eb98ad637ec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56a29b4f2f51f76ce3c943b4d2a5ef9b0650eacb0e8725e08cf4f2be7d247c4585e9f04d30f1850f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c7a7983067a8b1c3c93c1b7b5b0d01094cbfed724cf8977aff61970e422e1f1178162c067568e22;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9974b6d6a5c44f66d8bbf1f6ce661f34c3c64e29fb6319345592d50fa78a025b65c311a2b59135026;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9eb91c80b6fc9a25933f834560049aad88d809410c2813e6a74de95de7982c677f19f27a1f76ef994;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48c5c61bbea81c607b3453e1f930fdfee0a1a45f6e250200d5b151e8d76bd1b3ea005beab426febda;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1c329dfed6c1296476fcac80c912165c518206a0f1fc3a6bab852d8ac877fad00ec4aaa0c4c34bf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9dbac67940b2ca8dae334aaa09f535bccabd4731c593d122d8ddb42d89846b9f2620221f33cbf3a5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc24811d8719c1b69b16d305886c7b761765c31c42e974c3abee5ce91939738e79733c33ade5e187a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56cb1c937571d4b0ccdeee4724a0e8da694a9a7f585b6940ecc59070c8e2d6835c8d8ebc228eb8726;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31f24e7912b733c741c3312dc7e07643e684839d7bc391be985cb4b06ba40e41d1539d541f826d8c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18e90dab3b2cd0759570d2d406aa231b6433c430e6480b5e1d9613605ab84c61783a4b5900b5729e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf89da2c7cfce0850682110e04486f2136a1f901a2136c3f3a2378dca2782a2376c6582a1f3d08e1e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he95f522d62bbe40b1d6af844c42499fa3ef63f504d4bf252f1de104c09bd886ec9da60cb98f0e4c4e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7923658e78d7d039fd0d7d76d79dabe19daad2791a09dbd5dcf5114e8060760f5c569d5a1432e8f6a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9330a562f31a180c2c842cd195307f31f04e735558c3aa9e5417f2c3d5cbd1879a2c87f1c85205690;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2deb509a9029b217dadd1166b089677be4c21384122090e0691eff4e90b0338d1d425f2ee645d3e91;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2270a3be96ab91dade61c63e112a52028a04d0c3e123ec2b51bbb2c63847cea4cbdce33cb4f3b6d2c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h266118052e6ada49bfa9c8b09b454342e58c9bed8e381627531754135340301769ee47d27ceae3f9c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2609e70d316ed02569538b1c8556fa7227b4c26d606d2627718566df0129a8e26c99d7a55b6bc7495;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c2a9ebefeef9a180379d9c18dbf09ce363ee9a04659d960df4c7fa5aac9914531ba2311c5d795c94;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cd16d2ec73095f0e845cd4f2ed670b7f697ddaeb5342c95cc68206ca1e3fb7869257563528bc48cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83b4fd14ed2e1bdd555679bade6f4a58e975114d874c1ccb65f7e5d94e6d90706a13fed3e20a21ebf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2a8ffd36cab21d1eaabdd5fb04e6233b554bddc603c439dcbf1f62f0d4659014f41591ffff7f1e0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78baafaa6778c80084c5f87811897687214811f63ef3a1d1119454eb12e8abcc8f45f050a72a81e3c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c0fdb6fdfe8a4b0918a90d77caf5d4365bee287b08fb97312e9783763b356d6fa3ec35d34a627c4f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf749b7495bd7efb24862c5a2d6365a9709802ec11b2346ee9841d76a0d5561431bdecfa11fca94ae8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9abdaa8eb806d1ad94f427d7dca07252708e0121c5aaec6ed27dfa6b26fcf997bb9d9bef5dbf87624;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfc674fc17e8bda3d75302e312261238ac14c516b210c61dac93faecf0ee112fa880ce55b126e0051;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h840a2773c2c73f81a1eebb921cbda9eb0d84f7410d6b6c88b3d11ad68c8dda40f644067097b75b3f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3fdb3670e47805ce8e380630f75016d2401947c6d99a3f00836a3b717582f046696104cade71f37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d4d145f24a4e7fe6174068884139cfe6a2dee26b1c0fab0ea71dd1439d6acee28241bfe8b2126ee1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93d2dc99cd23cd237ec93968126d092d4420fd6ba542eb82d9215b227a659579257c2098aef09ff5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd51794d75f4a70710caf8fccdec51da4e1977fda098b34933358372cdec17f92f2a8d5a0d35c3488f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42f6a2ccf20aa997e17b1411d218f433c93071067cdfe1ff3858e518db1cd98f900ec082045b14965;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h309e0674982220d5f42f1bc28b87637850649b8ac9589c0e194ca5fd495bfc69d229812bebc88ce8c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha01b2dcebad919aeff3e70ef5fbff4699150b0436dc8062b651038cd586137dbe3f5e21f8ebdde3d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe3cc7b26d98c3c98ff29dfc9ed032ab8a1694b50ccb03e02f4157160398e3ddd87b431b627c80ce7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7e6242e6e65a360406a50c11fb0b2fa36d10b83bae20b89d4fa3d891aa34bb1ad769a2383dd22bff;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a8ac744c47b4ab479baf08499d556a96164709b628cb2119b6a5a75f169d25a93a95885c46b87a9c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36599649a8f7b46ea5ae87b0e7fbef6089d0158d0b410b4ee5cb4a272cc66b98d4f5685790b0a08dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c758aabaaaa0859226df7dc14762a362104a8f3a89807594f3647699b96e12f19c2b0aad069c1220;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61cdbf7f83b6fd182c2cfe874a366686acc7e6f317a63914b11c6ff72d1f423a5dc41046671b4132;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0b95a4dca7acdb75359815c0ff12cf6cbe9ecc5dcfbd91a547c2ad9f48a43d4f6155bfe844ec55df;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7323335778cfabe8819120418ad6ba237022723388b557f6d5a3a113f98d198e51fc6ab36c3e8b078;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d9674534569a31f79393004318cc426891246ee6804c25171f7b59571308f0467a43959145bea829;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ea0047233779c19179e424a854372c9784af8cc3c7361c81aae67b2ab43b8274b617509d2a339f23;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcca1c5644282c0ca8a7150886bc2372514ba9c59866af1420025b4211a02d767c1337779238391ea7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24ddfd747b09b974b0efd8f27c4fb898721bb785136fc708e8fdfb80970723ddbe71cd6512bf04894;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h825724c393f384e6d55dd6f28a73ade22c086485c997155c1b2d80fa88ad7ca3b97abb9103988e44d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62439f51e9dce446ec15a22d8891721b88eeb77577703f2a0886f2779898370a7b71d0a0ce622ae32;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77b643cf351d75fcea74bb67817d013d739f4e13f1aac6a2b4c7678f08348b76b93c76985df5bc179;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1da3ddf19472a084192f3ec0cc882c14b6e957cf8f42db70510620e5cbf058774d5b509a89d7b803d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ab31d7f2d2e14a71c9c28d1afbe1cdd2f980100a5aa6442ad3ce4fa6f91ce0050419153e42cd0a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hade2538a2957cdc427b7831ac2818914e64536a4432cebc7edb9b0331efa2cf95719dfd17631c27bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c341a2efe34f116662de3246d1467ff513981653e28620c639e9cca2e22fe1dd44906d71c73a832d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d8a7324c598c6fab954521cae56565368f95df23ffb267edc2dc5ef8f128adfbfe9a841347214a19;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74d38bb3a7dcdf0be4aee65603066b2ebb2e2ca5e8632ead12c01c7fce0dd13e342ac1465c42ea345;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8941a13cfcdb49395d2638701f706a715953b126c21287964599b48f3a82845601dd82e767842d394;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf90f9c9af71b80dd229b8675d869ca109b7aee0a48154aea20bfbfa906a0a8e51a5b5868888688ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5fb2d64c91f216dce9212f572019d8440ae11505dd2c58808761178ff2540078330555a1e4f7ee504;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h250e042b4228c86e4319ef44f4152cb68dcf397cfff11ae73f29398fe509daf6f9ce35360a7f232a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h863b366c03e771677c6d8ed6fa6b8d27bf82806f0c2ff57d09a8c6422d0e311fbdbdc51355596b0d4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd40d1b204aca245f54976ab6bea998dcf32c1bbfe8f4bac3b8603cf338b986c0855d6e33710b93c21;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf75204c7b624f3dba67fc35fb1e4a4862072ea8d244a696c0457973e7509286a54b98c5ba5518c26c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3c8277603189999320c3dd197d3c842585988076b5f559b2d3a7f8e79c55f960d90dbef25d29c135;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e92fc4a6189ef01b1edf66637cbe28939b79b648c62a3d52f7c91ffc8e496f1c42d4748b0b5911a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45e7436e5a2bc85f38dc6d32d6f4b1fe9a0706bb373cd8e2434e1c9b41de7c82765c502f330855f0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e8f85320cb64abdaa468c49eb4d207b02e4544e746148d91d116f19dd50cd9db92ae82ea5ad6bd99;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8499bf26fc801a6b4edafe947ff889e52ef23acdf3100bbb1d4832ff06da437d288aff0dfeb5a103;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he95c71c9893dc835b84aee9841b9b6127a5eec44e83c9346c4d9a635982e5dfea6fc62c553fc98fd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfda04bee4a4e318c1c52ed3c757ea5d7aba7ae0cab00b45e610183b483774fa061f1ba3e0238bdc9c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcccd23bc70a3621443a773b9dd96a50e62b9f0e8a0be8d0d54be89ed4d64b1673945c2d40263940b4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6271656d38f3f5047b4bc8d27feb821538c89566e7cbb3f218157bcc9054a5d6596bafe3e85f4cb8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbf8346db402be7cc3318383793b165da2974af0d0df18c098d6a95a63ba0ccbdd2f95651fefe0ab2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4723abad331449784b2327be872aff7fd9456a1dae38d06bb99729eb4b7fd588007bca1ca3c85b78;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c6fc19a0e156b9d7ad24d9dae3dbed99d0566807c441a9762b2347921e02b9af46d9366b89d0be33;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha10e58c371dfae5e4a48a9d822e10291e14be75738d6a23082ca26f2705a5c5e9bbf0727ab0bc9c2f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0206006dce7a2008088e545dc071feb5d76d988a554f698fd4212c874ce5d0902a7e05654e2faeab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1dc324485f952b529629de1cec94a82e0f54b3475a260d02de332dcca1586dd85f6e6925453633605;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1bbc06068eae495fdc4f004e320af8f4922ae2a7939322699e71e561d81f0800f162ac869952e2c3a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fd70021272a4e5b2766e79466c234a49c5c03e3b5568a95dacb2db1f50c65616112a269cb0fa0a8f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h726e70263c92adf69ca8f584dae023f5888e9b48d2019948a807b8aefbfa2de8d30e1c21834e41fad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha460b8a3b2854a55952d6817ade3e7debe37de12ded9635f05f551fbbee77ec43b4261c1e46b4ebab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6a41d3209d8740b4f00845470161232becd1578e7fe3f79bb6e7c60df77decc4e793f3aa4d9b4f71;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2bc853963d5e4db800ccf12ae3d0d07acd090a039aa902f89ffbe55ee0cb4c6fbba8312aa2e997bd5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbb1abaf18f6ef7bfa49d18b8679d156693f6b07d47cb949d536b9bbe3910de4824274797b256ee54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha355581e0dae6575a97953ab0dede186b5bab2ccc33f5676a05182bf059893ee46d8078e5f5744e89;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf22c6e9d714ad1e1b5ba33706f59b6d098999b78e2f8cc9cbf2d445e8a3a3b7b710f6b3a8a85ccafb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5bf1eb483db04425e5ad6063652edfeb55cf136cb7c8654ac44886689f4940534876cf90573e75dcf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22c3db2e83c5ee48c83a69d59eedf8d50395704ff554f7026716ceb788267ceaec7478570588aefe5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb99cdcff3e9b40dcebe8b0455e2ebba2cb14834de71454051e7b9f7e60c9fb5b9fee275e724c7e453;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha21ddc7b9b53e0d152b22b3fbf5ac870d5915ded8f14cf6355a3ad23697cea035e5f104f7dbb7bd7d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4163a83daa10da0aed100ac5ec4712f37fa32af75cd519492c3a7ec880c007cc915e7472ba470d22;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb096393fd5d9ad4d5eb1f3ae75e16446314f6e83cc940ad127171ede3155864dc99dff1d1f8a7799;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc6bbe85a4244d263375a98ad16c54e7df9bbc04af41cbaf9c2e8a2b1d683928ed8fd63222effe13c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c2fd22d9ffbed63bf471762e9721a6c068e2516e33e54c8833092eaeab444a15a8ae794685b5cd8c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63767e02cac12d85f2381992777688149a6f1550cd965fdc3a4f1e89cc291b289e5e9c7f8df52afb8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47943f1d878aaa1f29027643ffbf321365166beb81c23b178e20120061020b6d36f793b90ac3ea90a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69ac72803e4ba0a22f544e99c5df64f6ed9afd4f5acb78b35ec1e76c0b057672caef7f1110679c230;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcad270ec99e04d9d58f77be5c3e1aa43604baf042d708aeed9c5265f7de7f88e8eed9d6bb1827c1d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb5c3d3b32875590d132c13806ccd9c8b493948e7efdf97e8a644a8e0704205a33d4e7b146053374e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1f3de55b1165c4e0ee067feceba5457036ee49d2f715e05f2cd19f8be00342e7e458e0b3ee498441;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b2b9962339a558cb06574c4f9fba805777ea154a4e7a60f28672de14a6411aa88da56a42c5c54935;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h277d43a88b729905477e970d0419053c9249934a0fffb9292300e5e43ea58c609da0277823e8479a4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1177791e0645006c31dbfeeba327b1b83a52fe99c8cf5188e3f749d9039baa189e6d7fd6799b7dade;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1133aea58c60eaed46116f3aba47efccf3176e80ab12cf8ecfaa9276b41334f5e9c50542d1360c64;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6fba080f71a44703146d1ea1be77628320c16d52d7990dcac9793dd255b7da2b9ed3c71aa3113a44;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf92b7e66641d64a7a4e635d01bf408ad807cda40fb26332d21a64145fd1b209e3287fba533240e88;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a6fcf7903bce275e0be30bdb7c266c8f935fc2bde2fc05833ebb5b508af649ada4f9d8915e6fe3cf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63c4f60e3aabd2376ac7afbcbc97aa0befbed6509d3b132d0e0175e6d80d94a184f5f3f66adce471d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b5aa44c7ed81539ef392cfb2913cd39331ba36b541e635bd99533fbdf3c55b34359b9009d46555d6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb85d20c1ebad5fa767c90f1272735b5fdf895ee206f0ca8a22103074a84ec6fc2d0e0a9535f28d61;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2afe5e6684a461e9aa417a65c294feee42bcafac8f5220e2a4e11e234cb78cdcec44687d8cb9db65;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he17a3d600535a508cd72de462e940681997c3ac53c6c8f2770a15ed56bad557c74f446ca550e91675;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0da26fededd96bb8626cfa67db4b4acd575c898e92aff57fd184013a40682061b03012e9c83e7de0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f6937940257a5809d8e162e55a3741f639c780e76fa880f5c2e58b964b584113861b0e26963d16fe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca007ae88d086f79fe0b325cf7e656203452b7b6f58fe00d7475432709bedc0bba4f703413b693e99;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h908dd29cd78363932a7ba86e74d6aae0782aa5ee4a53219a551932e47b9d8a7baa07b117fd7fd8c2c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d3aa12573a93abe5b5566c0a962cc392cadc803a8d61336443341532b32e3b35dab10ba3f7b00d1f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42ffc8ef6e41edca3ef6c7f6b46d981941c409bb235050f00122da03315ba5cc47d66b403ea41c094;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had96a3f2d9707212d2e0476590ec6c54b04cd2eec687acfb84853b091d959b33641b2110108a33703;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b81c42b1bd0778baef1369f19b641789403c30b765d2e2f0e7bdd77c0bcf8db3d7d93e2c40f7993;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf24a7a2aedd56a08d24cef9b3a5a0938d4fe5dc23f08f3ef4607235b33ee3bc6bff4456ff11e3009a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77371bd839f4536719d650d4b8d0fb1b7d2278070ecea14b573342a0579121d74826f2bebd5d55ce6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31bd7fca4d56350277457bf0d15e459a73a61d9b64bdd09d12e9ea4f151bfe219af31f3891d0caf75;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6bbe49dfac48c30c227592fcdf97ffd4a6f3a90b12959e44f0b549d8d09d691a6d7809d7871b66ae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h717450cf5c1ef8e4ea36e38b8343c1182208e01503695b18ad058a2295339c03e1eb392c78b81d9ea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha549f892120fe92870b05b6933c90a829621aacc20984a4b2705ca9d07a5979bec0ba73979a6f9adc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f777b93cbe388bf72e119382c09fa014a51c17e8dd0e70e53f1c5516558799dcc55347a318e51552;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7336bf18b40b288136df090b379a949c2f13be063ac09cbf014c82f88306e70c510e154802a661b44;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c798484d88cf521edb1b275ec7ed2a68132dc9775d0d04fb885658393b760acb86b1d8dcb0a41748;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c9f78fb81253f273a16d5d921b55053d1c3cb3a3845bb6b1598919b41a8df0617a1d016427ce76cf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbdb0a5254c2b368cf03bacc488642dfaefdae6c36747a020a698e7e873839f5e1bb414685a9ce3f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30d5d55531f3fb80d5fcd358fff62fec7e622a1381985b2b2e443d9a30c8010dfcc442f51197be4d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44241cc8e63b6a9fb94914e9ef10ef5321ee22eb701bd91e835e409451fb24b14eb2b99256f51d8fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7852ef3d29e843082a33158904911588ac80b9e27685b7af214d87bd87d696037a7743c1126a85180;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h135f958c3046e6afafe02b84a2f884f0cfddea5391bea2eb647719d68a8e2982f44214d8a1bf2a1e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff5fd3c283e6d688a6ab918ae484ad31a28b8e1425fe8f2e888eabbe75823ffc2563716bc07bb3d2a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd90ae82fa0f82abebad068800a0dfde44d5d86c0ff1b80ab0f9cc21c21a6ae5e66f0fa019e350c979;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bd6099cf1595d413717fcbf8f7b3fdf642baea88746423d73da4833c8c63f801df3d2ade55bdf07c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f266e7262db3d2cd095391a45cd272524d66409136bd10b0e43f1fbfae57356562e2c81c14fbd73d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fa8a550317545c87bde0715771293171fb926b6af6152c45e0cc9fd7e9a5b666c59f31ae294b8942;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4420bac1c60433be8cdc040ec369d15926d56055c0b089149e6cf9b5bb8b313d73d6ce32e7b022563;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4dc8d7f3d262a452d7b8ccdf568f3cce0b0a997091c260367ba3407e5090649723dc1983f7bd5da9d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48c9404eb760accf7c862552744ef9b74b2091ddade5878b9c519a489f6a7f03993bb405769e7285d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb3bcdf290df97d84aa5e78f9c8895d65c5332f885d8d303c628fc3407d4c80fdc22a51ea231c5274;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0c09589250d8d28151d3e720bae924a5c35a2e9e641085eba34f5ed47ebeb647a7254d9ef30d80b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde2c2e882b9c99e695c8f0973d591cf7bf0db0ce471099286c0020c2290ec2073020c0383741e3540;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12326d23b9b02088dd4b4d6dfc8d718ff0aed200dd8f402be7c88a6226b31b0ccbafe7ca9a9073007;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bcf0e72dbc9c2af17887bf65d122070673b83bbc09911c8946e8c519f894c99b4faf1efdb1ab2a41;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb12020753363f87ec2ee8723e5f0ee11be359de37e3b5ee2e38c347cbf41f9b8c4c4ccb37735f8757;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f60e17372ad6de4fff8fe16acd83d6eee42fd8f60b069560880de5d8bdbcb7b059f09a5642d8d96f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7288fde4c956658876b4223318c2ec76246b2b93c8a72802cb60f7ba8fc61fbd02585de04ad1ba84e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69545909c1b15ea1a7ef7bec93d98e60a6e85314a556373e632070aee4c6daf5b19b115c693bfa184;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6aa29aa0a80297017973dc7166ab514497db8b5cca926253d2a93c4b27a053a6d3e836a9793b780b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5d2493a9812f8798d5530e4388b97a8b8651a335989017819c9ed191a5628224499ee50342c60999;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h587946eb6eb9e83d28d7313f4265fe409ea64b21c4edb93592f4130620e582be5fec1036d755efbfc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc4f9a68d4d8ab97790789128370789acf030d4ff209d1486a50099b004498115e640799205a5208b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9965c42555baee3a80fce0a83327c4c3d77a524971f83286ee0fa6609c475e397cbad38d4da92087;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfdd2493f18014bf876f06cf4161cf0a7407d1b35d6c35f785c9d7840d1a559b9ef7963160ccd4ad17;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d5a85706a500b75b21c69a1c213c4b26c87d96f872dc5ae12215d7276c30e4cf90aff0b25d35073;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2deaaf0d2a84fa949e699d64a80aa5a24f6825cc2f8a07e019b5cc60e61e94224a9810d092fa93262;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cf992565740acc6702a3c737b79ea9a835b0267c4fff25a6183decd8615972fc8c35ac0c3d97d256;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h562082ec87f439ae69b941649ccebe9090473c43bbebe3e820fc0db210c7e91cf51e17894fc0e26a1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97c738559c602ea91f8fe154d4f066241301a5244c323c11c58d16e1dbfb1de7863b09209a0f4c780;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hccd2d0eac6ddd7a2b46670f18b5687034c872842b73aad689a91df77ca883bc3be15de65147ee2578;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h868b8db44ad116f863305105172edf24224139def591c5a7dd76f8216010a65624a8db6154847050;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7340bfba52b1ca10d3791be47cdf10d35927d6200c2836dd12219d2db2fe43d38f2dd61010901e469;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6cc50b3cb7ceb7af4bb87f9d30aaeadf14b221b80e1ec158da77d3968d826a7631fd705f4f9464b8a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ea79a34e564951bc659890d7f8e1c0b1188e11d9921600309e1a13e8b9f77d08e0ff09280c4298c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4f92d537dd81c3e7b0f2f430de22df8e59b114400305e6a7fff23626f6e00b279688c6112bf89efa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12ef813909d49d8a9a2bac7002f0a9b1999c3f213903ba0550f456ebfbbd4a2041c4815b9db3b348e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd8330dffe8b8ce3e51df331baf9ee000e735db09f4f5bccfdebc4818c27b82b58e66bb1e7ab659ae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b833f5853470db9771432a8fc704a7c2366b30111d77a4dcf646f38c8bdf2fa65a896747d4fc7996;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b17cf13f19f0de3b2683f1e97aca670029d04b507512d5d1a80ff3997a47c9150ece2d8b2b947fc9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc789d8f9a27ed8959c494c4351b3f7b215874972f683193b74e5de1cafdb6ea008423986a28c3fc15;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3097e395cde82cb235b53024f5f13e721b2b3aae2e1fe67bc4502e7949d83611e7240c20c80e31e05;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha88885f66d927f240b7163628c14385a7c4d7de439e86bcf7277b6c3f8127f60792eef82eaed51a3b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a69f4df6678193fd7289647197b9ff6f614a2145d77593b37edad7dd187e94d73bd1789353edaf47;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8fce97dd5bbca49e15eec1ae919df71e3ef7118afd0d93dab2759640451e775d14f25d3b3a21ee2a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h376a1f678a2b1cb4c3661ae7ac806214abbbdfb196b0682fe2b4f556a5d3a2231d00103319b66f08e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h682f9ff2d5e6d6819d1309f34eafc938f67ca482d0bb12a7359bf64a09bb0572e1053aa23c78008bf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20b69a162afc61d7fb3dd6fc76765d422067545c23b115a5a3a99851b91c316cbd44a6437c01ec330;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75ce449acc934675d2a1e8943839b6f1cc9d1dd0882f2dd88a85e6634cea515144509dd58b89b659c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6746761120d51afcf2506217eab2a6ba71ec11920d88257fdb2b187b2872a2e2ce1049c6a9d96de66;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h556b775c8370cb19dfc1f6230ea506ffa0a07679d98fae4c8619667fafbfe0de7bd82955807a11ec5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89e4018c3e937df69210aea1625b2c2748cf8ad378080c9bda98a627feab5051958e9121c2129cc21;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63e3abd64b3504990511eeacc344a4892443ad2e30897f2cd0e5234d6f4926ef5dba50a2b54c2cfd2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ab44f3d6426aee5d09f8349b5d97ba8db0814d86b39d77d6e8c1bc85536bdb4bf0fcc3905a303168;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8f6b5e3976298d7bf74369def4d523de68006753a99e0d1089aba1ceffc6a1aba6e062fa0116d4c5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c40ee7753ba017b9d8e12910efba4b7e7b15fbd54cfc822b6bbf05339925c6400c19b97423f65e6a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd56936b3366102168e518e6356fe8ef1ecce129e58e3b44bc950fc19e999f92137d8530be59b75bef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1971e5e0591c660821f5367b5c55cfda2f90d5833dc1cf82d0e8c055753a2f97f8e14e1089e39033;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17bb5fc519cdc2b97f6e6405a85eb70953f4cc2914174b2f912da5f506d35b724fa36c7cbd2163d02;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc31ffd917c98aa8a6f973d674548310d9c4166de14bbc92355bb4eae79c122a8aca17a013b6c0a5d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfcb2d29979f47b4f0b16221a9a338376654660dde59d1b4326f170ce4786b8446b9c19e591a5bcc80;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a5d67b6150f374279e2d4ebee51650c1e49715d3f777dea494495f0f2689570b238bc742419b06dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68cf0b1eb3d54336dde1b4c6dd00da89ffe3e513bd99772ffcdb82e69290f370905fd838954b805d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7841a86dc93426fa8e9fcecdbf5ec729d64838619e0649e65cba561c13b24c34a0be4c28cd873855;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99975f67975953a0bce16c06a9919e218c39094ee05c43efc1072a5136198ec0cee4b1b576d34aa0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h618af987db7e3dd6b7867170bf9fd540f53dfe904b5999fd87a404b3e14bce86cb98d061b35b8fac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8b6b639848316f8855b9b8494d43734fae72e46745e945381ea0827a5f91b5cd4356a17a5281ceb7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he55d07fa2e75291ea4ed6c8601ead1be7b6903c98e8cdfcf65dec7b087f9d0e2488ac56aac581a457;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1aad5a8d2bf19e1e81f1d64561dca2128b3fe4bdd0e72e7ed6998590def9fad7f9c8d3331bfbdd01f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee601597be221e3ab63402b81ca29900685e54427629c06c379456317ea50fbf9c8f1a1551cb6b401;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba2260f44fa2a73d9fbe54dd5f4fdd2f300e5a18e59eb9256a9dda679dbc37b2a96fa974244ea7e1e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35bb3373e8b3d425ee4df290661b6fe7169f3346674ffd7f4f13a0fe15611d8f93adb25f2e3539095;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7819c71714e23b8c8cf8e71649160bfe4c018feb75ad096907ac2fc516a0205b463cc68cd88b0e5d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50b2c6c1fa2bd9a51120ccaf16803f0fbb594b9121382e678169d9033a70aa4219685d7c8ed81da62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcdf67f343e6b1e62f30da0883e23b78bac585f29ec8f664d4a14ab99b7967fd8526600dfe74629fd0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d995642b7b7986a303abae1be73a285cf284ac9a6a4c1ab550ea3626c9fe168d84a345d96c916206;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0aec48e17f3304269dc17f397310c6fe76c7622aa00fb09fa802309d3dee8dbb35f0a09ccaaeed69;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha14b1916a6fbb16c45d6a3f59c6620566fb428c13ddc7545b03c861f1bef09384d2f12d0fcd41b636;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d1ad627860821fe691d397e51a2fed36e139873a7e050aa92dd31a03dbf18af726bed18d60b1a293;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1258fc9f1ea4a718a26783e2024a944f1d639af359c6047721e2c2b0f1a62cbb605343aec2187cd7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda405acde9087e4357242837ad48115c0ccc892382862d144baba1ccbff1e3f08655574475d2f9501;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f10380e195e5651ffaf28858a78b5641269d6ce3a5a2e43d7efdc59cbf97f91eeae1c59e000a5f2c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3d62e468e72d8338f68942eab9fc1408aedcf2b6ee49483024150757917e15701b38cb0720253918;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9c8a6e9be5d12cd2e42df215b919dd73188f30f8b83f56ca80dfe96a754f79c9b87a718a3026fd45;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff014aad580f97e5b5ac721f9aa4a04252860c92d4be65859ca2226e0f48d7e3dce91d43f4c3135fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3092f8aa52b70ec4513181e0647e3bfaecce0121445b08e718ca913aa60256f126f058451abda18f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he30ee3a8553abd9a4041eda5b242e398674dbb1991f868af65b766dee073b392319fa6194f8e5ed70;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefa732d6347cdf820ac784fbf5e5f62b1f966457cdf4486402af587e1f7b4cf1dd76383d7889c410d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b40d09e5d15227543c534b9d0a2e5f6d5e9635e777b3c4671359ee81039a27e68048dafd7a0fb39d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h764c730ef4f541279bf90bf23757fc79d074eaa8b8182da95bb38390243c613b72bd25125753fb4bf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39ead52e630b02fe0f8fe2695d481f49e2820c49839294a99491a2234564bf9a77c27d9c128e8d6e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf28ddc3bc9c5a51161959ae1312af6725065fe789dc04458a7b58cdcff087ba51a37be30fb1d956e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6e5949e917c925ba03c62a04a805d9deaeae6bd11b10679217b006d722c1864239d71cd8eb5833fe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb8f9987a7dff2a60e7d34a47f36dcd67f5b7a306e56e7f75b2c3e143f5bb8c5caa2266448530f40c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce80b6751b01b7559b92a3df31c114b899b0a353c72a767a132813bd92ccc8a503364c769bd0db9c6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6f6c4fb3d4394b9a880040a162d24736b9731d9e5b83571bb5fed63d3123276d9a75e48b6325db05;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d03dcf1a93b979c1900e3a12c11cbdc0303c0b3fa24da6028962b587eb19c267c13cbbf0eb4256f3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab3fa7f8cbf980ef7b4ea161e2f7afe2dc3b9fb0e852e7905579d559d8f531895bfa447435ddc99b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4b1631d658d630c62490553c01920495db09466cf306653f52ed588f98b5942c282a9306162641da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb54088547dc78d57a1d6f6d527f1f919d4defeeb9ea74783527ba979ede71cefb5350b76c426d3402;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e1b2d106ebd5b099eed1cede791f9f42cd6f14ff1b4e25372faa4f7c0ba6806095ce0cd3f285d3b6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61da12833182799864d18727dd76d75bea459244275e0bef55db9aca661a56455cc5da57a5cf2b6ab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c452253f1938936b856f0b0ccde6d80ff53531fb446fcf75fc3f109b5c1b580ba8a9ba4f95b1b071;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22d3ed7fd333a39f8192ca17f354237e2036df7facb83578e86ae2222083f7507524f08b0a101a18b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a0677ecab0b10481517a6f64c4e693f713d8f9cf296756faa392aaacc64e1bcbb60985c952ef6384;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a991674cd5e1d0b0cc1be4eab6b4722f0a8d185abd859f2f666f07c073f7c84e6b8fb6eee0bcbd7a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84a8756ce62385c5c693b265585485a04b5a7129b83c2aa050d4ed8a26f1e22959b23e2c7721ee87d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hede149ba6acd130766debd3d9c141b88a8ede46ff589bdcba6bf3dc05c8b41ba1934c849cfa2e8ad5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b6777d7990b2e1896ae9068693fc3b278433fffb0fce5d11966975147109c07878396f43b2889b18;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3652dff21d9d06cb3aa92c36cfdff45a09bf5beca453a482bfe6c3067868d05ff9d5f8f66d6bba16;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d61b3f180f2139434c89b8d2fc8610a73500b25c8c80b164020a0d76b41ac0983a8740363ae3d3a0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86f9544a6f9276c2fa9e0bb3990f35ef98c8bd66824984c5ee948be6908e361becf472eba4e11e259;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2b399a92ef493c5e60dd3420d6a4c6e50395fe8f5f8c446129f8f265fdbbe53c819532c94d84bc2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7e158a19b405af7824f8bac127a5dee5a0bf9bc5ddf21a3af42b80a12108e490264b79c54444f061;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h297f0c54474c1ca79051511c4d7a94c766230beda8a79e109d74228df6752d3d6ca22b9c9f05d4250;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc1f5269945507f8bf97ea55ec647b305717fd00104a812061fbfd3804904dc7a249a577231c3a4f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9024df5bdd82402a58d0a74620c0754880d383e2a7b50bead872241b9b3c90d711d44bb071ac89ccb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed57624daccdd0ccadbc2ec44e6112d7b985349b817365d3d8d5da3d1f6e05cb6b5a2b00d09e52e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h603c8d6cc3ba5d46c05727aaf72578cfc83f23655033bf87eaf29f2637be5065b38e38508948d3dab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2754040ea3291f1d5ab2e6b4e7031657c3ff8c62f0b10c532811a7ad3bfa08dcfd6988c9b0a916fb9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he021ad1858140ee90950b6135ef8c6ca41088e46cdbaf2abf836a3ab4595554f236cabd999c8cbb3c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d2fe592a07431a9600328a7e25dc94de07d20b7a3a506bf83fa2b41b2b6fee76387cb227f3c7fcf0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1e8ddbcc02614c105abd29f8c0616b36a555b79aed1cc7da8f24ae1e1611a8b1f95b1e7f078cfcf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b972a9496acc2ec6517e363f55031a7afc13307a256c84b3853b7b86aaf207eb468f5faa96c10cb5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5191308fe6a9d0e53c7de6ff368ced2b8bcd212ce088fcf366341fa2bf935dd5659ba6135ca2dae98;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f56b6341d398a8c10cfd47d8381bf677311d73e0d884ba8ba8e29fc7499cfd4d4bd64f9dc185f688;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf010f789604374baa47036892745d2d8f2532f69ff4eb153cb29f1c76d61ad9c4551944e582881ceb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9eca58eb35bea3dafdd93e9f46bb35e2658caed54fc6d45998e9c2ce223a6ccf7b82db05a883ac68a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6a1188a51114c0d40dd20d82f0ef58cee2dd6788c63bc5103fa75f744faee9b840a0f2fefcfe6ce4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea29306bde573d045bad68bdbf038b8b22487daef2d4f6ee81cb13c5aab4742f8eb0842dca6e36164;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbea8e1896c8b75e1e9700d06f08118993816b4b51e4ff3ebdc5108a0f456027bdf8b7f98a8b6da937;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a6687bad5d5232db3bb54dde1792a618ce6e3642eedfd9adf4bce1a39766659f3fe071e5a8a4db5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97725e67b640b27f1f850c4f08f35f8815d4254589fcfefb0741023e94d656c8003c5bb576c48fab3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49c0d967862dc8ba3bfb9524ae8b6b830f91323313d278a50bb4e03bf335c5c4947faaacb215e7709;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5dcbdaf57322e2b16279a9513fa6084c3c2bbe2919178e4ed6fd1036e646070259ac501f48a926f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1d8d7c054a2b1d561f2ce59bfacf1f9b6e612c0b038e80588e9b38c505ac9d767a937d35e76348b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9353ea0033d254190cff8ef8ec2b18fd71969888cc2169150eb8c36753288fe5da8bf3626a52614d0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb76e7af68f4ec6a5c638874078fc2d69dab480b1664d1c17f944c76b5cc2d6ba1ce74664eaaac885;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1cb460fe6a969efcac928da0e5601a5bffc52bc12bf85a6d555efa5fb154d411d7f79ee8f4362b230;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3e9499bf67994cf1a03c1f97636ddd2dca14a55b2c3403ace04da2fe3c6399f3b3f30f1e4fe53357;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc34da1506e0b644fcc90639e062f38f219f56dacf4f31d4ee3c17f6a26d9d156a2f860616489f2b90;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h324ef5ce4b83dce09e4653efd0ab2d3c6251d7770c9c63196731f2e4150aed79b59e962bf4ff1f730;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb628a13394ca582574301c13da88453aa27c7a781f02fe3e68c58beccc3cf94c8a23f0f3f76302304;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h530fc9047d050106cdd573f0a2c27c02c8ba3c2ad698d1d430d27b8f3f32c7b7d3f26f9bf4b8ab06e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c868c974b5d907be3ed2336cb1a17b7353753c0bc76a10b623bfb361d716efdd7a5e4b26b227e08e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23a4f5b451d3ff7d10e9bd8cd9e92b91cbf25b0a4371bbb72ab384728ba6015da13a44ae5c2a2c58c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcab77859b70917966e98bb75825e81801500d2a9dfedb834697b57b4dce4757d34e4bc23932bd570;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e344bc0b156f97fdcfee742c555dfa7e3053c96132afa6ad76559e5fd4d54d787c658a9163308e61;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1d86bb311c723694e79ba006cb23aa77948ef394eba20e5e936657c3df34de5630e82a51db0c72c7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f420fb03f359c4b5bb52f69be6a9b7fb9a86681c55030cf3fe485b26e7e58f52c5d743fdbb231903;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h625c441e17eb894c6df696dda7067d0b438219b71edad9951ca74b1bfa4054fe7c5177f6df4d34378;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h491f46a74ca08a5512fffd881a062c05bec05e3f4c798b03be83b9ca5db188966c8b6b613840c0a54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce93aa532f4f429ad6026046450af37a26ca5a8c4b2523276aa7a0f3dc14ec34b1d5e4d79fbd17a1c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h716ce75eb511d80934aa7d8018bb51ed2798ceb5399bf47b8d5abd9a1078ab2a275ed6056196c02e6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f2250738c8f36e5c91ee153fa7a00bb46b21106747f40781195f9c376c090f8370879a961b634a4f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1fafa22b92d53c912350c648bb0bfd0d83cfef843a4f42534b5bc1bca0fc055779cb21b2512d3fa1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h315e3ae65d82b27e2f9fe276bc9048b9007e32e4ce4336d3fc3d8d947564d6b116f47564ffa65eeaf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3fa28c5535f31f353c2e337a22293e130635fe3c2745b923f95500c5ae0d250c3b9e1c66b706f09bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64cdbbc00e7ef0660f10ac350dd42250c3495bb07095c608a997ca383fd33c6365de0d5b2467ae091;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h513051f9b363d8ac1211f0c1f41d9746de30155092dfa030129377e8d1c85bd4a20b3cd552728408d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1f15023b3e20c8b734fba412c600219ec22ff6bf28580693b2573da0a26c04315d2612fa06982c07;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbd248d2127ee69f30b4efc76a231909d0aef34a311da9a18b43205e358a46c764c4408a893a8f0c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a8d891d185879691a57166fa917716a2ca701006aea6494d0453840a292fead2a0866d6c8a88837;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf83180bb5975770f788425ba5d38bfe3be4bb435cd23a196722718f4106cde251da13760335632f3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40d75690cf049ff6e1b0842d6e1a8699ce1674f8112bce9f9b901c91e61326d4c5debbda3a46c1d77;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5509cf04a1c90a717212a7a32c6176be3086a94a4b422dbf87d2b1518bafce867d6beb566418b0f9d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bf9a5f74360dc37ea4de96951210e2fe13e99e9d8589c264235c74eb7274a891a6280c7ef3302462;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h819da3b0e697d86c68493794a10a6e7c0c31689cac5f42f908a399a3a173f7539c2209593a44c45f8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41055fb9362e133032bf94226eaac556f4057dff9e08500ec0b724c31cf290b7db053b53af3066a9b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he66aea550928e6ecc5b07374a0ea4104213f5e446dcf912a7e1b76dfa53b199cb535549d1f7f38678;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h793b9ae02c895b9e4a4a700da87eddd808e6eea1ed592bdf07330917d722455680ad4fad81d32028f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d0123d19cd41c7a932cbd685a47209e771e687ccc9fbd27c728ec758b423db1512aa51308539a99c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f19ae89b413481ba9bb6e93c0fa40a6d4eeab0d70d38959450073d3d66d74c9362ff4992d6f2edb1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fd6619ab44241d9e4f634e9dc01e8b1ae00430cd6c46814d8c17cfe9569cb9c459dc3cf73015d91f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4fdb6583cbb85cd0a03083ea05db0aa16f63b9659da2b6087d939bfcab13c95d010f0ff051920334;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ecf9981118fa092fea497300bb551bfe9de4bed1e7fe2474aea530206ee44f0b14e3408d62a88f03;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a8cf26d4c8c6be17a3a312a961bddd12425b326da3a854efc42b5b4b45ac05b392b0ca5b488566d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc518818a93b4c28c02b96c539fea47d70658e1b930b7cb271538aa303c03a2662d46a5fc91b367bf2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h317dbabf8068323df330c24b460adf3696c5a783731dc54b24881a1010521111d9e6652ab5d9b34a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf8a9e4056f347dce408bd36cabbd13b19dd87d810df5b6a107ea7db849dc0494dbef83ad1888b773;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h766622a5067b01beaece5fea82795f2398b81d53378965b1c681b3ec8a632c1b60a4dec5ffe14c2f9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb20b2761dea6a8d68bb634b70f814083ed8fd5fc5fb6fbc49f1a9b0e1a104d4bc1a4e859da443d114;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h358efb5276b0eca6d5f702a3cc44e5415e0de60d693ddb01fa53261c9aca946f9c8ecdfcdcb53afee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4567ed12f3c2beeb36eb2348f318383c0abf88ef02fbd97460fca8f630d3b9d14d0c03a23da282985;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7456983abcd4c9b3c06e6180a0d6a3783b37c3d1639f499f9ae3bde0498e948f94cf6a02a7d6b9653;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h603240eff3c7fec136f1c9c06dbec955b304957efd380ce2b45dc7fe7d792110505bdbebaa71c13e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6203a356d3fb1e49b530a82e4c3ca9936867656a78b55848824061ceeebdc44573541b4d2cfe5f048;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6740c4324b30cf26865ab3858c159644d8d5ad354280b71abcb891ae7db7b626927cc668b53a01270;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b1e4acf6d36f91d4bef490fcbcf11cee843d64bb136ddc8aadeb6f2cbf401c10e70cd148d16081f2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a186db5e4b7c264bd98f9609dc682632adcdff61dfa891a56c6002b5222432d520e13152efde00f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a8b8288fc8b0f4f429165f96e5b5d09094e732ea4cfd3a80ec500a980a60ac525710f44ff188d392;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e2b52a346c338bb4c7375064804a52b707c9a2794e2fa3e40cdea2688478a166907be040591e1ad3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb7835afe73325fcedf4ae5babab6f5fc4a8eeacc48b17449ca86ec60b92f5021d2d5ce64f90ed804;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he427793246416f0a77deb514f1d06166375041d8e51d2314661112d57ab739664fdc5c38836018a04;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3409c966bd6626a110d1ffde657f70150695cc075278533c9e45e7b3b086771ef9eca450819188873;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c79e7aff2a34424b67cab7132cad294e50b30d93524b1aaad940df6f57a511e925f1999c163840;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h586e0ed248b2ac03386da8321cd11e9e80f91e8c90826819e6d694f1800d733e31538a3e2ae7589fd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6177dd200b7e312786a070f5398e03c5bac02fb92247b337c45b16eee11ee562f824b9e1caaae3b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6824590d4496dc93ac48a7156f86bf44d57ed705cf3ecb9789eeda0f3f3a32b8f910daf3e69780095;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37da92a834042e16d82a9587d6473ef0b6b24487d004329a7c2d236659aeddedf4157fba8485b014f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7e259b55c914ee5258230d68bb7b1ee8eb6b30aab6f9423a258e60c21f021705e85cc2297773bf64;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc83669e9ede6aa026023dbc2685e4a3d8251f0c84650a1f369aa844ec360ccc8a31af05f3b3a3196a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bbc27dc33d0a86d2685612e9652d02eaad1b387ebfdb2f2b86b300802b5118b17d12ae4bbe5c2cc4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5f4dc134f3555455c47aeef9bed460d78335d4b21a37dd3a650187eba71c167ee6b70cb9d8c5f928;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8953347b4e4b5325d7d3932958d146f96cd7137e5b6f32aadd6e25eb4517d78fd802ed966ac936cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h644d0dc3d244238766c526fb1d141893b15b17fa5128b33b027e3fdef12c9a162398264a9f4777cce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e8a3d06d148a5cf85ded44748bf6342cab65edf7ec48dc98530128461bc2f99df3904384e1e3ffc1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74cf22d9f7239014c94f0c575fb5273a08f32a77606afa6cd32b5ee494aefb9575015213c61b151be;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha963b75f868ccafd6c4a72418a8e8eb14d3f108a0a22ea2469b77985c069a0e49fd8c82cc578b8ab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf63af66989c7bb60f63af1b8e7604e2acffdf05d9614b5bec6bac1f2f8e0ba102228c2b2765a8102f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b9a1b8a59b9e49e041c66a206d92648ad4e6cd43f60c8497d6d0de7e08d702fc1c1ea0d432922aa9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8525745ccb928772598b277469fc585503c454bc27115ca04b348983b1999f290a6bc0ccb2059b2f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c8433d49b3afb3ff1240c74c8fbd1bfbe087fa5f795db5b32114897a735fccf92789f0b9745a756c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd46a880e49d83b33b8b8b15c91e4b68976089d3ce508d379687743d184faf8391fe1120619619992b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1d541afe70a951c3e065788f60619f7e33ae7aba619ae8cfc00703cd281236c875651c60b064c742;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72f9b09609d5c3cb85bf4d8e051208652789d2df160e58ba65a2aa25d5f70b1a85f1fc3c0a4a0e3da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf54e11f642d5589a4c4771882ffbff031e9fc99811bb9cddfd7512c4c4e407fca0787299499fbe51;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0e2c046c616de18a8287386896c6377a1a6686c3b580ea52171846d75424560438a2e6709fa01d2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf35b3ef6e26ac0f5990893a7d6bcb05a38a205458a78cef8b6b7b74a4dc54b94391a6fc0c6ae6c686;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9efb39e798b70e364742663c763bfa85b8f7740d58bcda8acf6c0f09eab7b9f24bb9b68d4c6e4862e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e894bcebfe69c4cb61c7fe43756e60c43d898545f91ec9e557da8c8bbb601945a43230364b3e8bad;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffc0c901ab97f507315df8394ab4c3cd9f762c4c5c0bed55b4d57c0fba842df8474359f72a18169d5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1fc4f4d1818022f9ed2eff4c59bcc053c4f63adbfbe26811a258f927f7445c9c96ba205605f0d5fde;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2e4f3b1ef63505342feadb4220d1b9f6e85a8edaf0f256b5a317305874c8834323bcb7f07ac50cd3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fcf0d439791d76f494ca33aa50333fc33c300c7324a33fc32e3078bf0e08f77c4a9133e65542834c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf282717e68a6ff5ee81ed65af39e6ae429480d1b9f8ade85bab49844f8c895615d62406263533f6a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h863602feae5ef9069a2e17bb71f428ad1044397acf749e91613dd1dbeedf27869be9e4b97cbf28d62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9c551c23fbb03af1104a1346b021fffcb2f92da23215a3a1d4f85188422954048db64d329b71f1e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4d7c842b28f7a3c71cc32653350bbd1b4209ff72293f24cb02febe071a16967076a63c50e93f3874;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfcefe590eb055e750d24fd375fed842b0f183d06f1a7d3e336c3f00d7d4b1cc9117115c26cb41e98d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e132b917acb13a78b8c22fdb03f02afbade9ae638326fc144cbbb8f08f9f6de7f701d00b8741474;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60f762a2225335413f20df30261e8bd92f15e060985ea778a3bbf695044ed0f1dcecccc16a79ef0a6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1ad34f0f4832fcb66c9acaa908d9b6d9c76a0688b711249251ec383261ef2b6dfc6a44e192f1ca48;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heda3744a6544febdb6099d8bfa4d6ad80b7ebe752d97eef011680c38aa9251c74324af0956accbac1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26c14b6fa14ac5a5afab66626e0566e8934b497620e967cb864f8110330b00940271d6c1dc64d7fdc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfefb1e524578bb4af5509480fc536c2e67f2f6f563e9855f7eede081fa5004f87c6e79fe61a94f75;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h730b6c7d7d198c9b14f3a7e593f1993b266526b82a465ee33cee725991ef9cb9f65edb43ec64a6ba0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12a98e032e8f0fa9fd81dbee6a87dfe1dee215e51c9324b1d108dd968349654ad45dae5e2e3fb79f0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b368d52d8601a62d8619f521ce13d31fd38e389f7ded9e94a5e1117f3431f7deb7c2c94d0bac7fb7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf73b9fd4bd60833e675c6cd9620b12c7080c6824ebb28dbf23ab21e82bfe774ced9002a57714bfe3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h661579a0901dc69e6f103581d054b5886ef36e633923b70005160ebc40aa18e4a06ff688ceb1b6775;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h867ae4327fb9a84f30261ab10f8a2911c2517ccd1069583e3998ab55cc1f6006eb7ae1a7e63b5d44c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81054f9367f4aae145b043de0655036de91456ae8b02b96bcd6a508276121df9bd0e5704c9a5ea97b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc95af01d143b7afd81153a796216b1499a30676ac0eea07391f22f53982526320bad6eee6247a494d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10930c272dad2bc05448703f5105d5e2ab4da93b37fe771f2bf84b7a65e1cab9c03e727e3cb6a6c7d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h554f326ea16686de4bd8820a198efb1ce014b308ad89940dde28fd13ebfd989956d19bdee12818eca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1443364e5c90f7f892913a1f97993da10204a5123756e8f4433959cba9b090164226728f8c1d2b6a5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4cf1ac0ac9795a52e8e7be60ae3b6fab0b22d049e708273bea2c048330a99127bb921e0f4db6d69d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb5a8fc9fc97474a3ab7004bb47a15a587dcca1d7e5d6b1b59e1cb3810901dc244705172f5cb327b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h935161feaa3ff53a33b163d1fc2aa3be1c1586430a0bdd60ca112169791af3adc1656d3be4941d6b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6aedfc5e96e926b5d31ef8fbd135398eaa3eeb8b370027c6a762684e8942b794e6843c267fa1d8391;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h825367608075ede43d5e4476081aadf7388910bd0f4a42ed91ff5dbb5a380c515821b92e2635b8fb1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h716a697919127603b8f96b80d1fd2c16f8143172b7ac99602a2ce16fdfbf3eca346bb58517eef099b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9b97c360047ffb037ec71b1af7b81c0dc01b4c93d07d4b7ecec8718ab8019dd74b5b5eadc49acf7b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb825cf106e5a5e993f12e08d88ba3dc4264fc188a12bde3ce495e2fcfb63866ddbd0838f1785ef3a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8b7d41b3e6bc27d6366b644df4bb3107435d706e2d49b91e1c204ba5ce777ae0aeff688360b76ba5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h990ce9ce81585f6359864ea46b34c1e44b558daef0316dd065b227532391739b8e5fe861096cb6ccf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd78aca7674a266903ba02a47000e4d04ce67e4bdb2b271abf4f1df012dc862cdedfc8a8725b1b5300;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7134a0a9062c35d1e0eb94dba6345e16de8a3f82baa84e576466435fc03c5073493239acb09f7bfe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ccc139faf95fe4cfd4c90f79c1a36710e93a1f81d24131d2d76c0f15dfc0f6e8aa4677693afcc1d3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2bb5058251c251ba7d4eeb761c78256ede6641efda74a818750ddcb4906779bb27493b869e538adf2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0303e34755e613fc374e29fafb402e2bd19bd27243aa3ccf20237749c05d76290388dfb3348589;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b34bfb67b8eb91bbf6bc95d8592dfd18e208351a2ca8aaeb695b37fa4a0a259faff5cd081a2d7d88;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf1c73594661f83d98905772a1b9b22cfa98e405207d5fce3fba91f06bc33bf54055671bd1a54c5da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a754649effee83bcddb15fe2508a3b13b58ea15668b35d288ae3af41173d7683d2e1188c4e7e84bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cdde1f931ba4cb2db43045e8fa19ac6b15b18ff61d2f49385543882497d9198b6699bb92ffb60a33;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a3ecb6d9694e45b2438594f944b18df4add7e7647f525c4df621366fa725a8b7e33711b049deb71;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf5f8159700067488137dc362278f6178fa5ad94e87efc5b6df178c29821a17350c6d62aea48cb2c41;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a6fec8fb5172ca59f4e32dd0b5d16512f0343ea4105590c560930da027cb0b6bcf9d0dbeeb66db87;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb3fbfa0b2614f8217bc99ea70c4f9587c771e54712aed02369fb9f9b65c2d0ee30497333abc7f5e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h951dbad6935157c3e1fc764db716808d8038fec2b0a3edcf6e706ca8da59e1404a8c817789f7b36cf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8ece1afb148bf92c86bb6f1db7993bd7c8590d526d06f89f7d9ed26374fe366170c3090e45ebcaab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e2063ebec11ff08dfc969a8c042c6868fb77547b17b74ed07dad328ed02686929ca5df00b46e3183;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10e3d811a3da5f44e73c8ee1b12a453a4c3b41c9eadcc0e1927d0d934b19ecbef85db4d16d713ac66;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cec0351c997aaac964365940070ccaf8e00ab8b715e250cf60a852b3d2a36f76d7a1897aa46c2bb3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h588166500fd4d6a8825ea753fcf272ee70862f253cb056c1042485b525f10d9c54e9e0331eaed0ef2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd02b04396b6de938708a53af93ae68601131a9b515e0f25387eb0a6af45576c72d7a83426bb7e8c0d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc97dffb81bca03d07f90e89440244108dff913f968bd0b5ef112a22d3068513df50d2404d850dc520;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3de74151c55b3cb4d8f4a9c4196668cb38ae587cf104575d3dbd8eec442fba583b0fda884dcccbb1b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6cd8776d421bd38fa1b2593be228b9e195455864782bc7c848a45eaf534ea16d1c626128a05df600e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54bae37f6c267dd1385fd2f3ae4fd71065885ead3405d800e9aca15df459e8177d3a6d18ad8385c3e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2d5bd04bbe7b53d70bf1732595583bc0c4f3aaed858c80dce26ea3f58bf98cd64a89058b704ebeceb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf381e1a4b1c2dcf88183c144aa011905ffdccef0558235ce21627339db0c3dd7e5722af3cdf332787;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0d115ef2969eaaa2f6c865bcec4c0271810760066676ebebad0f570520bdce5076ace5b4d27567a5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefb2f39f75a875d7ebfdd62209840cebed29c87e7a3a3944cbb464d8fd8ed40f94f3596a24e38bf85;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb20a87eca408ac140d697c8a1dd0f853c21931cab470f15686fac4d246c396b3af4525f254df64df2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha84e740bee55f68465082acb8bdcea1a2bc1e586e237842768011661ec52e9ccf139dd69d2aa4a188;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f90621c7aec1fab5c667eedc7aa1e2d64ba62c4e9c5ffcf263b3c89fd311bb9802a8de83f3341ee3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcff77f8ce59aff6a7595369f58fcf52806ada8986defcf166b1f5b2d2a65d9cc28515ecba22c8831;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb96b60fa24d01735068d84bc702f45e22dae241025e1b6b3c4b931e000f395e53bed469b4dda7798c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h893a34c931c7a1ec5e7b0f547415610e5d52bdbcd79e8809b087cd68a6690652e7e2bb9be42466aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23182c268a130dc208b2367920dea8900a1da89785507516ccc87d33ca2ad5a111f3f55020f58ba9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h333f479dfae24aa2297513ea444ef0408cfc9fb049ead8554577a7cd7d7270460eb8bcdf8af02c4da;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4156f76ad3bf719b6c13e58e182e7a68d989250c106f9e37242d6d17067132871ac92b456235fcc85;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6ec3d7517be3477fc29549953bac142011c2b688362eb3bc59a49e325258c622d34ae29ed808cf7c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7fbe87d616d8cf07f76dab2888d20a5d396ef938776306652a0de69069ad537de5b0504993b37054;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61712022b6461d67d9d23b5ce962e39922cf1f59a3de086b870bbca02b60d74d5c15b54273a8213f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9af66e896ac7c8372d60a2bb3529b371e52fa1df3831fa32e4b56922b36c62ab9a1c03d10de453d69;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c1c59e76ebd2633e88c09c708b1a9b80cebea6c3f4daf72ca34b203e6875297fd62c4bf6a2469c51;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0488565d1f6bdd79962fca3770801fceec0d83473ab4877822746a3b8197f3d143f8af5eed723570;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e3cf25f1ac3de44ea9bc1e042fe68b63767bfb1aa3eda4ac7a207e11b29536164b532517ba3348d3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d2c5beaf30b823dd57bd57fb001b15e7c28e0efbfc0b7b598d5d05f48d547ff53294d9a4e6988f26;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77f8b12830c8f6e7a09d6bbd19805dec5fbed936ce87f435d1598f25e3b668070c6521ced0d4df1f0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1be3faed5b1d5937c5ddc782b6199b6be59b45fa130e73acc7d252a1febce7e39e47fd65933d2cf29;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbc7935744c78ceb626a6316e0aacd9d8f9d6b0118423862d3162cccd81abc60cc585f6259e11146;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31e0cccd3b3a46857a4b82bb783332b2381808def0265375b2fffe456531fbcb25ccd5b95af22c92f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2ca37ab299a9ab4ebe345277143de23259fe2a35649a5f983e0ed6b830c17e824b4c212ae8cc3f2e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he05d4f05ec70fb8827f3f4d595602817b4b56e3670837ee28ee291b147ac799f1a7055dbaabef7fd4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h880f1a0b6d112ff5905577cfa29600a600987b2974745b5afea3ec72cd556870bf4cc67806e30002a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ff863a78faefad32e83b83add6cdc8cd5b6ab8886bbde19ac26686c0b0e1b295d22fe284f4fc2b4b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb28a155995af1981d743bebb5c92ef4b2818dd89a2fc1dcad9512b247f7dcf85624e3008f7715a6c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd71089ac3f7a426414911d094cd0578fdf23686c04a4e7f2702fe9ea21af6ea8f1fc96d52b8a5ebd1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4a89157b12a464a385236cc7cc9e4a8967007c3c72eb9974e4e82ed73dedffa61179f8e8275de9d5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60b1a604bb89045de570a36f7a6f92f50994b9fab14223d0f37e88968976cd3fcaf59ac584e2380ca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd610e19fe0c314ec71f49336dda01f7b7c6eb52469bb596b26df6d366c1b5ca06074aa8b7ea9a11b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c06d491f2b7560eb99751395d7742298ce8ae3d4057f7429df20d87a974dc6d18c842e5ce49e9310;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h638c9412d423c4f36f432136d2d7a56225e4fb6edc6919d79f962641f7b2a90c69da25068b2d2e813;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e19fef31a0f43f6a49ffd92eb2f9a0c8e9a1c9d7f116ea6c22e42f53ea1309f82b3766838a916b0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5dc5ac10efbbc887da6be8b0718625f8013db6ed5aac6f978899aa40a135dc01a9144e3f3403dbf5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf43a2cc395d2e86aa42e25596bd6fef72300a013ee933b2ae218c22f98897f0c5be8daf71411fb7ef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h378943c0bc0163e7a4fc272c2ab6e08955d379bfd0007e679abe923317ec00ff94fba80562379b636;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a33a3c29cfed7cd23f406694fa520156ca2b4b3269f912bc334234232e34ccebc1818e6c3c218d54;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11caabf4489d811ddf0fb9839ad9c0e386ece404a98aea5d8b224817f54d10d7b01cab425cd83b876;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cf6ea1bd1da8e19e66b7e0b3be831a9c8f2a4d35f510757faaec2dc8cf0a60598fe8d3d108c7b7f9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ee4d89ee75d2359528cf6d07f0da3c7738c2972949ae74206b8e6613b9ae15dc1091ed72e52150ec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfeb14b6ab02cc9d56a0bf2e9e09e4d88efe6238bf16e31d122b971ad60bbeecbb3e94691f6f7aa663;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h918e00853d3960a4a178c3afa7873a9905e572ba7e198a1b49704895ff7999844d0aedf7936f9cbe8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37850c2f3d1eba6f853078ecf3211ae448ea850fd1e83f783c1d95b880d65f1f270ef31250f4c4167;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6837cd85839c56f8ccb146f8f1289c3cfd2f5ef417cda341635c3f9c2ff03414f62e2ee17db3736c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e48838db6a7045c7d0d43d945bc9cfc1e56419c59410993f8597da125ec8caa0f5a1d5887cf9ea3a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h155ca5963156c0da9a9a6a54ed8bbf8487daf033508830db13829ef2e87ca336b2c54d84c746dd65d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f14d72cfe0b2ad1a9b03bfca3f98ac280b67b4da995942a4003303904fb4d2cfd8ceef656546ac5a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbbe1dfcdc150de9958c3f595679d7c67e50896f63ec72fbc0849e2d962d2106d8186c42a361e06fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha580b41e67826e31541a13ee7b8f513bdc4c7931978ef823a6a22243e401746f966ad94ebd31e8dde;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a980998275037a7204dab9e91f7b230e8a7594684acaa7a293811a34ec8d10e32ee93d2421740f21;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65e11fcfaaf24eb36d0953a5c010da470588b61ee230b3c0df368840fc2f7c550030ef96c24a7d753;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75f7efaa3ef1477462e5dede3dfa8da90ec74d1c45d157d95155750cd7f5ef22c913511a0f4d2be50;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6eeac1f6235f3fc494dd2a7c8af4d8b3711b0dc0e07823668cc115fd58291deebd1136b4ba8fdf177;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24230cbc34c2e2e980cd09e58b5c3a5d65d609d93eb2cadabc807b97ebbe3b5d4361dc7099513d6a8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6119ea33a92c3d043f8250f09f113422a122355be55aadf2712c77eed48bbdfdcd6f0d527f7b2e2a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1d3bf8586c29cd1918edc3d82dffea436408cf5cebdd7a183414ac639783b1d6ef62eba3896a57ec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42cb4ee585acdf8c15ab8c662402e09535392ad66e84d44d091b4de7967a76e8698b8163248af2abc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38f63b0296c33601d68b73607b20fe8f060423f54041d197277105a78ebb61ab9486db88537cc507e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74ea9046938e196b8aad3279eb1517baa7f796144d894ea6ee08c08bae195215ce34c0e6cdc9b6e17;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h379801990b1873470be07dc605faea5b1688855415345a9115c5b5cb83ccc5176698911e54a6081e9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b86872819ffb02dae8d446ac7acb4c2c804026ebc6dbd7ac3857bba285e91ed96abb0ac83157d5f0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h703566677734f9efcd18054c086f8b99448eb09abaf98357ead030e074d30ea5db8823e3c7f822e5e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca9d203316fea5cf9297eb1650b61ab7a1d5b9331e029fd53b574196b3825fab755fed216f83c7367;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefb9e3ce6af94ee068dd629716f7e2bdd04c6744c2330264589bb4f359b320ad33f1523acba1ce25;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57be0b0fd3b1ed5f35857b78d734c994cd31ade2404f02c8c8e20d5c8a6f8efb69b2fd180f1e547e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72d0314810ea85c5db7164010ccf70acd1247e834d04af89c625eb8d60dbb587a29bb0cec6ac43bf6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae80644b9345381e0df46abc717dc275dec784c91d170437d6dda1c8f54fae12d7202c641c89dfcfe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52290191559c75d0342d19aa7bcea7a8f70595f8ad8d84a16d829c80e7c86ccd88a8a9f263a518de3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h54e61d485736b4ba1c297eb156b818c852b2322c694e8cc48014045d6635fb9d5ec89ea5a350cad6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8612b5eb30c2c84cad49b04a7f11d0f32ff51b4be69f6e8e2a15b8ebfa5a4ceca8ccf225455299cb9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h290e66f8e5d10b3a9e93690db31159b7255e286a080c2d6b9b8bb6af1712e649c08f036b999c310bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87652f38d99b7e80dbdb66eb065b628d43ea917473e794a46ff4c725db492b956a259ed06c996ba62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hadf9bf7816ee1d29d0255a6efb20eb9145ede9dac3e1b36571b7906d06a8624d85bd4c08a57b06824;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc85157aa56aca97bc5c22f09dc240be110b6f9013afd544e4316cc1600611c3b02fff04ba6e16bd3c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h800cbb71695e1bc508aacd4be0486575e763bd3a705ec6f3f6b2586663758f6f7f07db45231d06183;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3763c3ccab5235deefdc020eef0afbbed4354c0e4f6871e9596ac9821f0b0ee1ee24405b072a4de2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h362491f62c2c10768757074a979c87e434699961da911ca93da3fd72c8b4cd37ecc2045e95194684b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6867dbd341b7750a6a5601ffe51a46e758ee1dff1116b5a34588326349db18c622a1a3f7548104f52;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11a84ceaa38aa527a48ec9f23c6ad252f5917786a3769fb32a6b93a7715d24518cf1b77d16fd9c17;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7c6629f6e0d8919b3ee92b924cd0daeb8ad07830db483d11f9f62a2afc7b8d1360ade1ba70f689e6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3aa0ac867914a98c16971469159dd8381a601d8b31dd21fa70f0af6154e1a0e1a0112ec08b7245fd2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7aad726c8b0cf1f0202de5667e3dab790aec161da16628019f1ca1bafa34d431524dee8eff7505c26;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2a943b71cba0b84f135cd7151876e5b86d488b4b22faa099fdb6a9427f453aa377b3aa6a5e82956a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c7c6fc8ee83d39990afb38607c5690bf3a81d2b38119fd4efb6fa0c5c8c9f0b8d07e525506c5cc95;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab69df39511b0ee0d6b12f37e3432acb07ea8023f4db4220db43f7aaa69bd01bdfb35af95b0c339dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c207834777de250a76bbe0ee4f11e73cd698bc5813d239ee63db6b6e7cd4d38bf68a45ee22417fa5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd6a57881580731a49e9201ab4e778a4de583e9175f22982263917f5fa84ba1fa70932378d54916006;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1719b8a9620deafbf6b1aae6231fe387cd69f6dd0c8ee97fcb5573defb248e6ee81ab72bb92a375d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h92ce8ea176ba7ac824ae59b752ce52cf764390ee8ab511a1760d63afb129310ddf7891a8c4bd47106;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf7e14949caee28a5479628c55affe14784a558674aff2ab18558abf0338da36ffa951b7c94832c57;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55078b0081c158ebc280d7bded24a44339d588014302f75d4e208d8ae9ef588e094b7baa40fa10c76;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9273e4760d480681a82b156c62b017275ed5407c78678cb7bb43460569ab5ab4b8a7d0cba1a14cf1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heab9a3a280b6d8a9f7fdf2146406f29768d3fa07e632ce40d3abf26b54152fce5102205ae969861de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf64e72ebb70fa8e76658a708edb75fd8f8df856320b95717b5bddf1b50c21527ee4416dc78584bf56;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc7acd309cb1a284f2bd8ec35e9de2f59975f7d8721aa406d1723d1398e88502ff88e274b6b5e15c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf186c1b1a335721c4a9d3c79ff4599b50ebba368e6530f1b1d4002fb208b7a3a619fce7f7c52eb558;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h375602a0da9dcae935d265ec2c811e3cb43612989859770fe1e17dfc97dbb664b34abb3d1d5e012ea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h436b73b33756581c319f3fd65338b9d17134689a49f8c5034ca2efea3d8cbb1e4ba0e9d4c51479dd7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f610d90e936a7c5520537bd74dc78dfe4d1fedac5d57fbeb4156d43af49e7a3615fa60e5298801e8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1cca0bc2b9cae221b8771dcd12d6262ab9fe00845e478a9b79ec22b0d33ad9850c900f2a8d4c2bf9f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h874d946ec2ab000217741a8e49dbba488d9b0625408e0ec5ac1c79ce475d64bb840977564ad9ec47d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39f7e447d5b28bed7ac5b016b11d1108a11facc8e103b4a31ff5038d75f528f849eb38e49714907fb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2772a34a810c82caf7c65644162c49ee09bc0eaa0a38c75ab47f2346e4c7a139e9edbc4fbae5ba4d9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a5ef1325d17d18ed326a289d8fd0303582554f3d002bef8d3edddec7919d954f8698e79ada841105;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcd0186e94669667d0a8a7e4b4a840b7cf794cf21ac06ec40ed1f454ae85f7e44dd6f682b8edcc2a8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf26b5d7088d0baf4ec09bcbaee0768075e0806a396943559eb7c5e4b15342af2b3071377f5eaa5ab9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc4520b25a434b4210e494445c5c7243d995f411e5fb327b1d14c963f032d77254aeeb4d6a58b4ae7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd83b16cd92fc334d5f7aab0612ecdcc9deaac91de3b66507fe873aa3692bee5556e3def5e136ffde6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he36453b2c63d28fca9914d7d4103b0e902ee60170965591499b7dafcfe547c4770af2d3c0d843194d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h669460c1e85f6af8c859704924d366d2602cad3b7c0dc4300608c6fde55118000c9ae6c41881bce1d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h119e8fa29f806b0235e7f26c07ee5a87d1c0702dc95bb7bb3e30a71d0e35243db816271649677f4ba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7b5edf924ea306094b0a321fcb7d14e54196cb64972c140c58bd25339ce4de1c3062a8a42622ef2d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d38119b6a6a498010a6900c77e87a6c187b9c6ba2b341352457017a2c1a24c2597e62360a9ad0cee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0ede3c934c2c42a87b63d9242ce6d058ec68debc18c516d3d8d3d60b5182d2f43413295b545d2ee6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb32a5d7c424861518cb29c2e56364cdb34bf349b2e5e768a1b5c9596bce96fa46ae4ebbc858906cb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87be888f854a401d04679969c3e8ab471100e33e6623ae9a19ba92555e2e88e52e27b75baca448b09;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h412ea6209fbea2da3eb987a468767762f1ce2285c997311f642741ccfb73e6d1da532ba57c3daf3d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h957c3f7134ee0175f39b40039575805ea7258b1b65b431257517c81ec615defe4aefdd5992be8747a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a9f0d0e3b46fe045b63760274894f35de780ad6d0465d23d73acd4b2c034ab3f0099054b41ab5f3b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24678fbbc15ddc48a21197028bc198b8b162d5f11066e0f7eb888b9b5600f78f22142dd9f5f69e17c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb94b7af0cd0863c5b0e0823227357760e329de9517e654bd7dd9e038366adf269e4cf7e4d53981eef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddec669965c5f85744a5170ef57428e14d514a240366fec3111f2737141819f459d830a6d5eb5be7b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28a71732bf1bab80c7f581ab326bbbd6480d4cc0028c55bdfe5fbd92642dc915a0291693b8ba6b01f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a54b2692f10970115385a4217c94b3ff85e6676967dce886ee2ad597cf3559bae02adef907ced9f7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7bf7a0ef5941b3f2153d7cb54a1d57d65e821fc0b280fb654bc61ff9d3baed3a32aff91061899ea0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40472d1871c12e6c5187d92361ed2395f7e157121130f74e60f8c035ab92f98ab697ffcb8416e5a91;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f741bb6870a6a058ee33d422fe7b21313145f4b949537ddf73872aaff5db3f823e3705c9c40d2c21;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h932cc2530311b483c40a16b4d63afa52c33c782d535c19ad4a70cc5d3519b00c4f31e853221325abc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7611ca8b5f5894f0eaa7b2e5a09f92bb6ac77418a440ed315d48a37510bfc3833e32631b15a794e85;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49c816db04319a9ffb963eff050a703acdd64cd60f414874dcf4be3b8cd90755961e1628a5dc6bd6c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28220eb0a480bd59ac4d9581157a29199742fae78747eadacdf3c3296ff8c2c917fc1c85b9cbca315;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6767066849fa516d36510bd9bdd68fed30771f4454c50c45152ccc475d090af1344b9acca826d5aa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc80b0e144ba5eb261c8d59b83aff10a2bb21b042cb72cbf81fff70fcba24c0081bdcf452ab8dff87;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc4525a5e37d7db3ed95dac1aa27c206451e91910261a8043a92b437edc66acc152dcd60ea515e75b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87517cc013de964f158554b2c04806992cc950fbecfb06df09b420bd4d905deaf1e3d999a1509f71d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a7251a71dd2b750916671d60b5882b45a28b3468dd390cd15990cfcda05c8c56964a654a2e3e3d25;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2242b76de19750e925be118a52b8810abe4b705b59165e9eb280c949e096c6ba874cc639235f94f31;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5ebcee00662c0bb1426fe6569ddaa9ea94a57ee8c8fff0652ffd4c9a5352556169745c03a0c08b8f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b17ab508b7add573d8eef9d46a16390ec8261264eaecb23d2f5ef98e25fc7fabef48e4c9d0d58d19;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c9b58562b060446c4c65f6d5ae851e45933aa133ad3e9fd591536d08d2a3a10d081c40ac0780bce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd78dd3bf58f143d6013c562061211a2cafb043a74488eb486f4e2ee12a29130e205a9f4575369fd99;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9eec1734cfb9c4c825318c87bb7a1a44a520b3448d787eeade3fddbd30a6c0419f9a693180f9189ef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a342fb39ae65836c853cdf675e18eb176731a88579c0e9f33f6857634dd6f1e65151d8eecd7bc190;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ef5329010783447be3d15555dae166db1026de69dff232f474f9713796cfeb16a64697220e81fa30;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc43c109989045a7dfa041ed540a45a9b692d27df5e58999ea57ae0f8b57c67b98f11ff53bef66bd84;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13a37e8521a7f1317b29eac77a8455198c80b96b7f6dfafe8b2107dc9f4bf3bfe3b81257653d5ea2f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb53770aca488fc9581ef112361cd420b191b3d9b4aabc5fffeb5108b100579495d56ee76eb174049e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ad99e39cb0539bb5607c6244b2714fef5b9e3f0ef44ff6093f1b977cc0d267d68790c70db70449ba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61aea7c1c26c53ea096bc1c7abee2684c1b504e2fe3bd2877bea6cb16584b9a6cdb4ca1c73c8a73d1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habbb6aef8248eb779a58d830ce3f9d54349184e45584dbaa2214742e6742552a56eddef1c39b7f217;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h312911020364d241b229c7b82082823a137a21e97604d77c50d142891a58471866d5f0e24adb61a62;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40fe875e374ef71f115c985f9ffc3bc549a9378cd19d3c8a624ab3b6f1ff054dd8df9dea4b665cc81;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf59e8567138bb728b93e03bcec3ae1d75b434e59fd406e650766e9675784419f2fb906063437ad895;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f8ce81c0e0e7610e4469139495176981e4b6d9528e06b983db2484176d60223af583a00497c6f8f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21f9f92d39df0b43ca90db6fac868fe382232ee9cb7e9ff2b9c78c16fda20124530af9f8be9eac415;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ae709f399c59d2d2c23610741628a3e749ce975c18d10927989207b38f3122a70792e6ea39b12149;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f756247b157f61f09f3ea4ca6c8f3159e4ab9558845ed001b8ea9f2687fe9f71b4340b2a18645c6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f5cf9fca8a9fcf68b4b6c54243bd072c94fdfaad521222b326bc8a40229c85a00a56dc8b985f6435;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21fd6a63dcfddab71b853429f0020bb2127c81379e469e99979aedff6c64a9eef79b5d710e5a567a3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a1509e3d78a20447a8cf620e9cabfac289d48741df98be587d10df03d471251a3b66ad2d13bf0fb2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65d3107ff4e68f372812c0a58fcfbb239d3dfac91d892baeacd0ff75e75e4e494fcb7d2e633e04be9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97e82b07efd00c5c075e70eb745e9553c8f5b1aefc8206cc11d9a92617d95c245093215a006302f3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he04815ab12d3c1029a20c922709d8640b8f7b23018d4c011866f5014ea3be7f375bcdbdc8f7cf5081;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf20a6ab0beffa79abd346a8465c1ac455e234dc6361de94586fb8c70e58d6c6e50dfe0fe15a0c18b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6eda7ce9e65ae08b3ed9380b47b88de91e98e26dccaf3c61a42f9d1a13c98cd3c4afc524d9a54296f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76fc6d1171e0783d561a864dc57a60930d0aefa0a641293608ad695d5e2a04318aab57869ea5c4b7e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7181b53c7368880636e3f3cb0ad18cefb927e1891597688b4b1fe6340786982002f6377dc38d93aef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff0d4a4d7e4e2b954819fd87a8e476e1a407d784c4b4e6abbbdc6a0399a630c3fbf184a1854797c39;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd45aa59fbaa47d71290e334e5fd3ada46da73ad4cd162f01aca54e7c4db467907e4f2b606b402f63f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h669f761696013b62028593c05024a953c819e31e48aecc5b550aca3460669d06c7c7315a44c2bdea6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5411f0eeef1dab3035bbd41dd0ad2b611aaa1ff6a4bf8f32e725a9af2808c72025181ed7292201f2e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb22d6ef22fcd3b4ded1ec3b99b103d9f66688a64bbb3b154ba7b233471de877186ed2c0ab79065665;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cfc87dfbd3ab849fef1dc426a8a76c52161cf945f0a34afabf88ae201fe959dedb555c0f32797e2e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc94a9898eb2bc05717eb62992d74da44ad963b97d89478950648ac56d881e2d60170f8cb55a0711c7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1832c76587a84b40302dc1b977fee3e96b64562830f4f8936ecbd9fe7da7061d77a4555460df281;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1d058d48f29e8c726fc61c51bbdad80344999c1af8b6f535e3d8c36d54643ddd748cb8d0c6af0e4f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7fb6091f4ab8153a376976a94c1f213ff902d0cea4fd40d7d522a006005acf77eb5b34bfee9669829;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba12d371b6cd4edcba65ffff8a2f897a7f76de0ca162941a404e51a7f84ed389312a12e7c983942b1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0000815fcbaab1591d9a56f27664dbc00c8022adbefe491d64c894ad24594911b194c2084b42794e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e7e20e64eb5c5120953c5e38538b1818a9872e3711a2a821abfe662a3ecb9f71334a0f6f75ae2633;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5db74aadfc00766e6b8d39f6d421954154bbe834b5b77236dec11e8e1b4a83919f435ba6bf050777b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0e5884b5129deb97a531904bfd1ba03c375b1b215c9cb904d9b678ca4dc44f55a4c11e0b6ce7dd7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1e71e951424cc807f0433f6c5fff0e81f5e81b53454865ecdf7e5be801d4402cab8e09bf61e9bf3d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc43738995c604663f72c31d31b4d53669f38277fa2c2c757dc759eb02b8556b356bb9e6839eee5ee;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h150179b1ed73bcb7880963083dc0319ba08ea3b37fc6560e1742e6407d1abc6f4f7a713d02d16c1c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb369488e4b6ac722ce05a431676422406ed032ddfb978a4e364b3b4e4111f9c853d30324d19fafa5f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9aaa923087046e37d54de28a2f81c7794be54b54accf60430b1249119689b8d978cf9886d32e50d00;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc6a0d07f28ce1c2fcbfc11718bd9afffd413bacc76a35c617244dd25e9d02c2303ab258e972f068b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5643f1c23570cee5c42261f01bff6aba4b7779f8c651d8ac9be19c2c531a8621a31cd48ebd57da04;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ac720f317b02f901e5902dc21c86eebb1b5589f627b2a3ef8d3cabaa1bec7d980aa2d8cb17bd39ae;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebed73692e5bd67d7f499324b423992b739b2ed9b80545524233bb7ad9145a0d3157b04e60ed67197;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f414a83a1310c09bba9de1273e13715a996055377977b872c4af0bdf662b7dc06e638eef02e9a352;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1b53e8c6d9d1a5952a23c5f6dc4a10f7d9e98be4cde031b1528731673585c5467c4f7e78ea007dc7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9afec23b4e056239f6805e4518fc1a093305ebbba91bf2053e33849aec54a9d2b264f5cc4941d6bab;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6954d394fcbec683991a3224065771b0075e31a3163d57ba3fd049139e6ee25fc9cc270896c79062f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac08a997ff1a2ea4a14530d6b02a045e5fb26e9d58f6193ecbcd8b32f81359f80288c53946c889577;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1dea055e1a5e05f2da662d07a2f623baa16bcc06256fa82c9bcdbd7c10b26fb103493907440143cc5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e8fb0492e6c383f8d15b6e452ccfb03856485fb4a12d7ff81b9b769cb368d53279d82d63996d973c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h524e2bd90c04b9bcbce504e975c6bcfc29aecc69142bac52bd4a8859cbcfa6a1643db0da921384534;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d369e3165bfcff626371634efea6853c48140345b5f8dff0a53205a4ef7745fdb874e818cb665099;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5bebc1c4e6a83eccb2ef8c1181d0af47d721af638a89c5a59e68cc24e0f5d4b2eb1932bc4544010a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30358cda4ee95833e086bfdb798a13974185c224d786cafd0a48bbd140aadb4eba88ae2946e123b30;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcb52a1d5fe702e339ee8c0d620da0edde03f4442d270573274eb241ee63975e984386bb4ade7c4c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51e5237a19f550b8a8ca8c3b188df016d72a584ab5fb53fc789c1dac08169d1b369ec42eb624a9344;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5264849373f130a6091c74f0ba22f23ccfcc97d08b23e3a3134575790e10e2eadab7402cd4c434d6a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe8172a2258927c81d9beceff4a826a0b4218dded42f738bc58da1ca0d2015464099e79e526b2553b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h803b4ae2b148e5d36c25e5cd161b7cc5782e11def5de894a4045a308cf22c138e8798fd2145a95c5a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he77f0d5ab6aed4e45138609ce972bf6da007e0ce6dba97da85dc7a07d1a5da8f95c6bac9924f9eaf7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1df4f862b563d73e8eb40a4d76c8e915a4f9514630112ca462848b60a51e1998a39ba5cd3e5a74aa4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a599432a093680e6cde3f35b7603e0ccd696580e603e0b2330382cc37cf98fc53eec98d9eb99e767;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb53f697923b97b2fc25242998e0bc21c04c4a22f8d64a400cdc4a45776896718febf010e88a31c7dd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4a6950a7d022cf242a46ab88b4a1255428aae062194665c41398f7e9ee0f96844714415e6fab941c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha97f52bca98b9e09295576600c76845fdba7cf2fb06c50b584860a9092a309c9660c0d89dc3576239;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab425abdfb3c75110438fe0f9f8b890de766e120b32912517bdbee9736ea126e57c07145e791f4bd0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h742290b38c5ea5cb63543bc38766bdbc1efe84009e20a1e8609e99f9a47a20ae239863643e81d5978;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h576c4dff04452ddedc2dec5d4535dfef03d42fb8a619b30f2f38d51c14588ad0ee5621d6be113a124;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5efd5e2ef3684ffa792b93c66e4e220160affe08e70e0f43ba2fa57ee1564f71dafe9a6e6e0b5eafb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2cb81bccaa7bb2421bf9fc64a61ff519c5e36c37aaf13650552f167b15ac4eaa7ed54ce4ccaf7498;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c4d2566cbef8cfd6981a625a3ddc0969c5c2198903abec18092d31052ab360cd084fc93511fbc022;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h177c407a9867207241fcb2f100ab9e9f2c2e60a4f553ebb80e4112c1700a83e3d0cf4f75fe93ac12e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ba116e5e420d4fc0b579394abd9d5ccd48c90814251005094d95709e2b9358b5e75827df711f124b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9081258167bfe6eb8c4ce8d3bc8513ca1418b3fc9fe75b5c641c2f19206e022ddeb35385135138824;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50fe8cee4e683df2aa67f074e731e6a23cc0ecfca23c3559c44a83113dab2aad505f4b6e833f43f75;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc99c27ef9d55559c8e640683b26706f5c207a68951920708cb5df2ec8ade65ba4c6049566405e863a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd2f16726accf924614102c42a18158f7c16f9207b2840e7bbdef6c402c21d825f36f1e01be0476b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49002ffc8a1818c7a91c7553c8d37e11a68612f43a01aade132b1b439ae4d1356043e901b09cfc27b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb58dda1137da81a09ef954c28d9a0614518feb1e4ee97ffb0765814aea339851c91a7059a57c6f03;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddeba9a1ed5f94564b4fc4ec200d9689e03071e294f6b2e25ebee2e92c2927b035316a6d8442cb8f2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ae8dd77267c608e2521ba75cc36da23bd893cf9142bd76d1e328342baee598899ca0bb05a68e46e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4206dd84f6f270e726b079ef75b15372adb71f142f8df33b88407f49e54c5b9e68cd2c0f46df84ea1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf0a35de0df4e623954d28b097ddbde97ba0305e230126528917aff57a49ec6ae37ac6aa309e59d00;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc939e1cd8140af5b4375812dae0f3cac7587f1cccbb95017a50b0fa448db5f7dc2a6bc96612549e3b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ecb787bbab472190a4f1e2c917000a6326aae79ccbe733b1178baf4a486fdb992b775dc6419e1500;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbc2fd436a67148ea1ea5044776b5272ba91c7da1d36e70750c088b8d4e62ae52ec5733512cc04ea3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a1d13a32f95acd6bd56c9d80397d43567ee056669b4b3d0e4d4c5898d22ef9381e09787ffe3c5b89;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17ca2c36e39bbc8bd95eb0028abedd9e9d3404cf5f2a88d4e8505229c2615893d0f60bf60d13cc3e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd727670f70aeddda57e872d1098466aa366d4ed5880b2308f660689fe1505837616d7167895fca711;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf9a31aff4a7e849c504e554c1411e9c37b856d319ac13d19f0e92011b4bba5d45a1ef3c622f04495;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5634aaa1602215add08cf16be897dffebd1893d2ed1311bececb8e359b9283f9e6f23322a248f8414;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64f515b5e41e2ce2e4ef2eb172810910d0cdb98df19564e3f602468b7048f41de6bd6b46142323e0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91505aaa7097f3b0cbcbbf90cfd49880880863d86a8dfe4ddfb8e8026ef9abfe9d96f57bf6d7d5b9d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4baac927d0eb5a0bf862e71f10351a06f7e5d87fb9d0c559ca114467f9361727b3b00ec6547b5c7a9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1695e335a904f7d4d84c6a5f752b4566d7fca2447bc262a8c5f3ffdeda58fc3cf791e382b78f8bdc3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h500a7a2b66bb5c55ac2ce9c8e1bf8413f7cb6f3b5f613fdd7b8280c635eb201eaef874c74f9971bd2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb5ee08fd82c9e92e541c49a25388c0f61984dbbd8a5114a5031c0fd415ac5bcdf1ce2f32baed6e8c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd415eb777236580258a6a888ea63df1c6684d00778cb0d0f54f3b45ddc464dc722f9e3d38e8e26c94;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he10433e1224e99312fbac4fd925fa287f9033d63a88b062f1a5413cd18b922e98159c776db761e111;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1a3aa0ebbcd8d8d2fdf64f499ebdf4ec9c3aeaea30f06c36af22ef17d68c27713fc6a7c6381e2b0f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6ec99e48f3a1e3707f53fbf19ef5eb41b3511a40119a50a7f11c69bc9e5af5e55b2c791bdc4d216c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d210b7404a04623554e5880557138816101804bcdf1cd8f280d78312a52912213b9bf3098947f417;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf26039123aca47e05927780713104d46474281d7271a89e5f0127dbab90fde0f076906615aa6d709;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5087df46c0807a826debf0ea9feb4004ea2e68b1747e43c43af005cc87d877c693c0d199113b44bea;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46bb8b42acb439bc6f523895a20ec47a3b286a0480d613c876f2a4ec03df86f1f598cb0a9d5ad0c37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee83daa72fdcee7824e25f3614841d333fd88579e89c43bc3c56c40c0299f3a331877ae34a64717f3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde2a5eb970bcf64161dabe6d967fb80ab46cb91afd3308d5eebe423469179a198d42fd1b43c923e2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfa781c45b53fc77f0b48b9064e48f9d9121cc39ade0703a68435cfb1b7f77b5e0f1296a15a17f7b4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37419c36fd97528ccf0b5a7d813f43d7a24205ab3ae7445234a69237fb14928dc12ab6f8f36058223;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f3bf89c94a3dc98218e6170520416e5086b5187494dede3cf01ae0bd003b6f5610d9b3560845e751;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c44d631035a5c208e755af36c1ec20ccc48831f8fbdecd1be978f29b832348d44c0256428fe2a01a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc890cda838972de533e5173b45619703630b217ca86e1ef17ce0b14ec0960f339b1e70ba6f1aabdcb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfecdf5a901d0dd562e11cab10a748a394950e3564eb8d21c45b6ecf822bf22e87c31eb8b8ff1f173b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90da64929695e3c59c8fe6f92cc08e8e038a9113c7c31986fe1f04a6c0c34c2e217f321e9496476a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9278aba8e1a87d115919f03663d052b2472cd6dce774ea60c3514d952d2bc9cdaba3bcc701ebec8c6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9556833d39e3ef3b2c7f141b792646446eba781f097938338fa40c73745c27d13118b7c8c9cb9ccd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6aee6c6d24df592fcfd399176535fc9c9ae9e0333ba8d5c61b40c64e8e3dffce492881afe0e331c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1db58ce17d893d4321720c882aa78d796cb853242343ced8c8191edb22d6876ba38f0e1faf09a2e43;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7ff0fe5b15594e285391425e686bce58c17d1dc555d820800cb56329d324b2b6082aeb44214e25f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60e7e46a4bf89323cfea859f6b58cd1db4e9ea58a6cd11d11963333ae633307a21cb8d2ec167a478a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfead030ece34b9df08e6193cc49e1c0b361f184904c007c9df1854b056785e5aa7b5290e396efb802;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h100293f160df665b75e0d15dfb325e71a54396273acdbcd33d5f3a64dadc22a3b39e61194612f9ff7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b15e67a4c69ba293b52266d8848cedc118b26cffef28f7018044252d18d60c9e4cc184b799420fa;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37cc3bd8dd81d2e0464cda9bba9f127b03179363f2db25c67d90cfeef4fc255d4f8d83e032c7c0723;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78dc9b23154b2aec2cf2eec24ea0e73c16a8d133aa4081b1e7c2ce8e47d9747ca045be6044446077f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ccad6188d48fc54e07f4d323255238ed4294ac57665140ab135040501955eb43fdb306917c49a307;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee0f0d547e7453dfe839190e9b65ec76663d612b9f13b7b66fedf985d953ba6dcf503f851237e3f57;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bf46e122a18129148f0093b7041be1f18347da20122c31b2e864920fcffe32c5c67e97570adb0f7d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b10ec54891e93ffe8254d41d6060bdf45168b041716647d393798d93f70299a24984125c6156604;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a3e56f01c65c4a67786a225fcf63459b60fd1ed81e1b1feae7cd551423c394d4b8f81d15a2c3515f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46044b1a376ead065e49c1261eeb9c0f9fb39a3efe760242e19b6a6b1c3c129e4604b07ee70238770;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6bd902055a38bd7728e899014230c4dc8afa7f15edd46918847509016657268e6b5d6a39c7972e283;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6b81b18a6215a84207d6d68b5805d220dcf0c2dc005210f4e67f742c418e9ebe3fa096f7d2963da3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56c65f7295ba64964b16775c70540129ef2e7c793f3cc49822660ca0381f0660cc038279b4977c2db;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h198bcaa3feb68b50f893aa834fda53b1ba8ecc51c4f52cddee5319e6257bc028bd2e27e9b2c266355;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c928616950f672f5e30badb9af84a9c15b51db02a8fc582a8f9b16073360a53179aa4eb99c7459f3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea5a4bea8a132add6ceeb02b523f478c2dd809f3e88aac53706d01ff214377396974ae5842bb6ca94;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c1ab904ad5d0d5943eaeafd32196bec7f90d6d3b348eb0355a4a13eeb2e16e8a30b51fc0efec9b7f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb48d1008e937c1d0df07118edaf022cc9a88a192c12c949562ba26f250c284b26b391bb457cfe140;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he694ee7acfe8a501ee96a3f72f4d6c0ae990ac22317df763dffd60e8645654da4168e9b1a2e350f4a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h172168ceb63c9b202e14484b27134400830a9e9484fdcb74ae97322e6327d300e8baecd7901eafcb0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53818c0ccd3e66b57793ab1a64bd0fcc6a98b5ba0672394da1ef954caa90dcb6e834a49fd47c5b20b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h880572962e7ddda4d7fdd83173a5601f38e54cbb3d1d8408aeb8d3364c85ae7c5f62fba6491125635;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac736c715beb3fe7e9f204c2a5edcd2f147611c361f2f09f3c1496b9bd33de10f0f50658152b61560;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94a58fbe652986b1a94ba5ffd63af05df5aae7ca78e93a98d5e2d9578078179cd53fbdc11a734c59;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5fed2d03defd9b59044f504ba5ab7a88a6cdb0648f14da1f4494aa1077c44cf6dcc3059c5cc8deb64;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h661630479fa2a536310ef30a71f4921d1436417787501b71a9adb5f5ba48f464aeb2435be7210f7b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfadec6d17ca2c81a2de79e4b2b7d43772fbbe787783dd1d8510ca98ef7001575ac400edba9cc8d862;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3fb31bdc0b24b38d67180cf426247fee931af09cba57e74d8db9a24804266c56697b0fff0a2fb2159;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8073d38a81ae52887fe541676a4fb0e442f4686ef9cee15c3c37862bdc0b07ce20b2636360090583;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31c62d8b20426e656f70c5cacff03c5a93f0f6baeaa6f3f2c72f3a2efc4d903782a2a7bfe2b4a571d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9dd182b12e018776aa6d0074eb703c1a52dbe92c4f14bcb6a84415ad93bbea08216f612385a58e16;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddc6301dfc64c5c7d03f748872e0bbb8ff163d78fdb04418b5e2e1bda75e4ac87639c1cbd94412238;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1340ed17339c4272e50a133f46e9d5e1b9d036b8bd5628b63bb386a82db83073405ba0dccfa9b3a21;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b26cdd30fc4ed633347ea52dc91b4151c2e2ff04c8483109f858a2ed8c4d6ca862bd2c4e7eba50e1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98807d17689eeec6242e0c11ef6d1db7e8a86a26cf8606582256e266344627228f37460b1031105cf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha174557fcdeb37419e932f0197a521b6f57911d02f6da301861c975d22d5794011a96c10e3151cd3c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc89a386696ec43a9cb9846adcda10c643d74a90614d9dd2ec5143db916a1bf04030fc568e22f8aec;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff4689bf98d290b8a1a30a94e921591de7e72e1c74166f808cda4c4e10cd5ea10015bddf52fff9ff4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcea0ba2a65747f1b8745cd090dba747498388d1d3bd8071a67a75bb6b1f72a9b459cab703575119bc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9712dd9d2a5ba10662ddf5e33d92c8e96df170e36aae96b9ac7e7a37e44d9a0fd7ef32a760fe0907d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19ead1b5e41323a77db08d031711d325588d03d50a772b26ad4b0bd9b585a0f1d9d3828cc2101a748;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ee70e121368328651773d19e2bff764ba0513c77d18c714245147223f006f4d2c17a9186202546fc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f3679530020ebe4c3c95abadcff0778b679143eef13f08bdfea0889fece80d9f460e6cb7d318dbf5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7f0a77c90f52b799b4bc9bbfca3afa36da35c274db3c3d9460b085e252de487acb87ec39ca03fa25;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h515b5fc09161739d849712869ac7eb607eb360849b2b2b2f09a8980b958e68e46d4510394aa4fea65;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h917b6cc24b3689fcb9633377681882a9d892493627879644fad5c4e7aae489b0fe66eb8f7de5ac383;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8bbaa552cdef13128bbff265c96d80879464205ce7416098571cb7a1913d6c0d93e238974964723a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h690d7d08112f9c17b17d72feaee1d6d07585465749267760898fb99c96fce7e6667212dd03e2a04af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h610bab7aa3623d08a1de2466a7b45012681ccdacfe6db0ef31d79aae176d55ed55bd0315e4176e3e7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h302360ecb033495e5bc0035b0e95c3b18c4e293530c090f8b06438bc1c78fc050ca4da8f36282638f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf6e34c7203e8d3452da587b17dbd5f98bc73df75ddb188775a5064535cd6cd54b1f26cd010b3bced;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1898b598fa12c1fc6aa56f7c33d87b8ae6bb1d04ce2a17f540ecd92eeb8fec35ce7b82912292e235b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ee8458358d2472f8445507930a4ae69b05c5f3978701336b8f98accc91251d54c529c33be0e9e725;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50eeeae7fe65c9b50e9d5baa8b74f20ad2bc9bf2036b9aca6d02b876051eef52a08afa967ee798076;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h38a33acc3252777dfb688b7a19f824f8def600fbabe3e0ac0bf8cb696f0dbc0df6b34db9fc2003db9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbb5ded80f5fefd5b3499152a3a839407d34d3468725d4ac661585e902413c46707be8658c7de39f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0803a861fee471da7e450cef2b6fc4244c49a32a2368f6003433c3ccecc57f3e5ac6c0cbb9a4f032;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82ed82c9dff04c419e463821dfa3ce2a3d86fdafbfb39b0e0ac115024f7da09a2fdffee380b1b99c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75a80497ba5a5c6b9e9fe8f54e7f8bcd2e10b99693276588cc27d949bd271a4990ebd6c267404310f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ca3d9ed22fcdf4290fd407fd6d87024cc1dbc6b84ce646212f2699de2612d73b719d9ea6190968a2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28415697a89349b18bddf0da601c2add7825afccc0d5d45590d5885d8867fe5a4717be00ac6442f4a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56c54835ff5ca5e948d2605726f77425a557eb5cd3b38a663968ab380561aa0bfa64162b6540cbf13;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b6c62c0fd206e8218f457f4de733425ce3808ebec2ad518784ba74ba97a10f3c5c5d6d4ffbbf10ac;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57d624364ed4dccac2ca963e4fbc70d7eab4978235ecc6fcc2a484a9f6df5cca3c0945e7b21417087;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9277d56dd511b04411af756cb2c11eb05879fdd11599222a6bce4aeb79d6fe9c0b203c87480701d10;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf49fc5260a9aadce15e416d06f013c9919ebe60bf60fc47c76ca5b80312e7a6b56d4a126539175e2b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3150acdc2d52c6b25c404c43b9c68191654c82bce580cac1d55c599aeda91d2bcc5cd828c4d87ca5a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8be1b23126db96b053eab3b3489711e6f8ee50be5f3e2323a3d526d7815ec1f1eb5fa86988f7f3eb6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h122f2a2c97e00dec021b4d02c70e6521d0ce037a1eb4ad0d1460f259cbc8e9af80d092dde3bea6501;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4851d068748a525ac8599a75cce985d6ba442e37e286b3489f62530f8fcdca6bc4c145539246a69c1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8146db6ac3a7fce744947b0d31288a27360ee00a08c995fca8c4b7fe4ae6dbc62f42f38fb637498ca;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0f707db23525899bf9c19581057e90104ed5de438a82941151cb1f5ca20f5b47a184eea1f07dc491;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a20407d6de55ed651d44ec05c738682ffdb7101aee728f5394563762e725c16537395278022eb76a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heff399c1e7750fa490d316ba32753fa262e2fee6c848522e35b6f9d979398aed854ca37f1c7d67a80;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73be2e8164ebf68895f95153405d88bbc4f5b86f1a145362d60aa209fb47258445445e6e9da529c87;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9cd75f5e4b3d605ec0f0c70f068c1fe04246a40c0bc0a81e765ef7518abe45ac6463e340170121437;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cb436d49f1959ec400c927af221be19b5f9a383de7d8429b3ea7870eb3c54fa40acaff329dd3a607;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc55183401b7929705178fb256326d546ae5b484bc4acdd88486d329ce9bf3d8857d34a8a09b610286;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h269aa76328c9759dd7af64f6368f16df7ad0b99554a6126968fb6b2859f48e41c5e5da8082fa201bb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb4028fc39c627fcb07d29765eaf894f673c18f5b23316c1df5cd385fb472fb076bc53b5db77c0db3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a017a5f6f876ec39efd51690f29afc9a286af2edda542af20bb271a9220013e7905bec32066a5239;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9dd07a84fb8cd40326114875c75cdd483df1eb419ff873e385383e550be51374cb41f73b0095e3519;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf6cf1021f710aec8e9e00ef4157b3ee6ce45f8afba4b888fe6af162b4369ce38b21d006341d8d90a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29cc13353998b4bb758aea211fe9381563252e8be69172f54c8a7954b00671fb351cbb7e942da7d68;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9237976f7ed34153ab84382d6585e60c583a59cd5bb073a5d2a23ace76b0319768f34e9d6a8708b2a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h937676075abb0be31a709abbe9fb3fd941ae6e997dc30f0293276cc5f414cd791c9bcf6976b00c77a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfcd1a2813bdffa0e9c3bcc055376bc007732b5a38b49e834b3c4245263e751486be242b532ff87916;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h906a800c8bf166042aeaac34d1ad81948b3831e1d2cec36e0862814af875ba7347ea603a60d7e9b94;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39f7855446a99880665ea3a97f5e654e944f4bfe9bbfb90963c1f4e904dbd18ca2a1ce5037c9a2a7c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h693f9d223b0ec227059e37b0ca87051533b6cbf9d909aad45094ec3f68d4d8acf6342a0da0eefea34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29a85b5cd9aabe17bdb4cf61c972a4491a0c79e4868d48219ee07b27fada98648ec715615df8f6471;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5af0f3be6a7618719c5614a1e60765a5b36081d8b90cbc5dfc5a35e789c92a098d63c77502214a0d7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59d7c1bb7fc08cd919093a394bcc2b1e5ae19aaae0738b18e850671e9629195d02c9cb865f304966b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc952a83179a6529cbb19beb8b8d0fe47e8015dc729b4fce837d97e796537b9ddd2c38dc898c13e6f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc278d059b7cdba7f9130288ef4768f6026b22ebacf394fed93f5d98546b58ace1e13ca7669a6b271f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95d01e56546a0fb41cfbca282a2ae5eb6de36ee1b42ee4184b4c7d22bfa4a2285b5eba5e864596619;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h752db620685c828f1ed95165c3dbf0be2038c8d7f7d2e5b74397aea0555b1b48db989b0e597776702;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f09bce0fbcf8846ea2e6e8e0124f4e6e5e272680a1b4f4c353d17c1c5afb21c5b985b586673856b4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h387fa160deec0745c8f3063e888785805df88785bacc291a2844faddca7d6c5160538d4a8182d8f68;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b0581078386b0eab96495960275779d26bdfcf3408887f1f8ddccbe481ed567a4863c32f04245cdc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f6c0731f4f6a64e0e5bc357bcfcf61c38656b8f99830ddc4b1cb4eb8cf9067523a7168a5442d9b34;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc443cd9ef16622f3f8729d3fb86983f50bb41707fe64eadd49b124a8f4eac0f6c8c345b1e70c5e9b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4a4cd8af02ca60df83f2c174e421a519a1f5a3bf61c061e31d221c897643b1f30045130351f9bae3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h604240ddf8bfd20d1445bae2722d515b92c3ccf948fbfb1011221d68b4066aedd5582ad202c0e1ef1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24e1a90df362f0c87dc07f49625877e0fa3d9cbb59c5e6fc010293f3216bf1021309075177453b3dc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd485f97115a2fef12b14d1847f30a7706e325b9123f30cdffda6bed4a062ab14ddfd27d9983e81032;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26a626ffaeb086f24523cb657c4dc247ede03a774c116e595303b047ed2e700ebd8cfb6f3c09c43fe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e3f00aaafdcdcc31b21fc09f796ac5e253a161c56461a41916f95d2e40f8b588f7eca3182684b04c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca9e2644147b102438a25a8dc2e3fb7af9ae4149179293ec2edcd474475ac046c9b2cbcc1affa3074;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30812c1c15c3c90ff19d11322ba059d0af5c415172eabdb926105af8c17a2ce72b54d07d25d71700c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52b287e7d47724d0065e0581722ef5904465fe65795984e777578e2959e5524d3335c8c19f6e2a788;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc65ee9a22f1baa31cb80096689d275d95325e4a4bc5cd4ae6e33e53c286e1bb98bf7ebaacaa5d65de;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15b50c53de45fe34b8874ce89b8b9f3c7d184581e348599580695aba7712e36fd8142caf1054557b9;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7677cf7c0b2691352ccdaa77ac5b500072c1cb2cd8e8fd5e560224973f65851ca24b9b9c0dcd68233;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7c35d5ba181c5355a354897f3f1798b6c48dbabed1056c85fa004549877ffaea87cafe6c3264d322;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac64b83ed16efe0a40d330a3a61f3a2d739e5d66e1adc45b24dbbfb35dbf80c21ce1c31e29d31bb37;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64db91520e771f9586b81ff1f9a14316f6159ba50068ef0bc8a8c2df1eb9e55b6e578109a7fa02b95;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4351e74a4ab4db88dda5514d46f476257765597f8b6c6e5a968473cac1c7a824f86c3224df87c8f2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5520edff0fdcacfe799fd8f23294e81f0100bb6f5c83e7d24ad48677d927366cfc225dde0bd049b3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h763eca454668d6886eec0af4c374ac4eec0341c8bc69dde310df1fae97d63e9d1883351f22080291c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h597cfdb54d03dfdf952f9eef0ea83b7533aa163c390c72172c016ecbe3fc019173b7cad274124dacf;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3788b81c941c54e0c1a9bb34a031ac5f457ee98f45452aa8d3bd1f490392d30da26d2129c7c3ee247;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h390a80685539fad283a0ec65046b6c0d7484cd6865a77c9973553269448cbaf59c1d0b4375f463929;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c51def7b608c64d696454d2467390049b9c4195f0a6a972a12e6f73dea2af7478c929ad7193e9f7f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c42356ab315abb4352fdc43c43ae24443403c2ac03c1eddf5024511c8e527fe04f59910054b708b6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9aff7e4fc38a7e41cf1c68baddbc6289e9cea9f5dc5321542efeccfce7d94c3b044416bcbf87143b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd709b6226415d34b549478de63f2b72502899cc5a252361d4b4951a6a038fa259e93e177e9f34ad0f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9bef957e8ad3e4e8d25487fa579c8406d97ec6961ecdcecdb1ade724909c4e63607283612cfaed81f;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55c3d6fbde2c2275db0c8c53581699a748a414e47e7e97bb34778c2825e6e56ec8dc4f0cff5e794ba;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e66b212ad46239ac5a44dd76b50059bf9598941a753be16796d5461adffe829ced6ea3e23e48bdef;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfac02bd2d6f6d52485f44e34d19d12381a11a7d426946249f3a13365b4c60cf1edfb1bee3f35ae607;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h216d001c2ae99a3fe7d911713ea715d1e741f9be29533abf880398b19fa9e68188623765345686217;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78b73850cbec97364b7ebe6205270580504777d10e0e2faa82a3dce7cbc9004f95d7a044155f34ed4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef1fbaea4dbdfaaac27da4a5b95b24d440460ee221dddf330ecf37623b45385d286f534ec7ccebb0c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44d7f6bcbea2280373ffe63d4e7771d80c04b102889b65fec6ef6572982c3c8458d15a21c5007108e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdec6d8224dd7cd9c51f79a37edf635ee88d6cb680348e07e585e0caa774b3ce9dc83f21157b27cc22;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bb62134463a4eab4f06362f3890a9a0b4e553a33b8795a2ebbcd8fe376544c22e5d42c305b957dc1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57f1c7e1a475e2e8e1ca9d23fa66b4dccba7fe28dac5ead6b59183ebc0b7c03fcc6eb257f5ee6a057;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77dacce3a0b4cb0b011ed3dcfddcdf399d03ebe6133921cfe0cf0f36add589fca67e1b35f42f04285;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d3e280c3b0efecb2581b037f3081567cc19f34ed48dc9ae68bd17957d63cb646b5487d9c2e7bfd56;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b0836c792b2590f927a7b2498ef0199f1fa251ba54538931641228b5332d39d91e059c85f48d172e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57855648917ddacba964dcd970ea0a19293b220d102ce6a8d48f91d8a65324a2cf3b3df7ae396c4b6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82d0d5c85db19f47b83c7fa73511ffaf38a3db8b6fde0baf24c5aa173b3271c879cc42a0782b78819;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbb884d63675d457defa45f23209868e4d02b37083882b07b4eb93e7efde9f877ac84637bf6f8ee9e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedd4d586f795f26fa9c1fc7fb7f8386c68cae1e4792e2ae4dd6e3027d3f1101eb951b5b1e0fd57b7b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3956090253d0f33ade43449dde4a6e5f581115d2389452fd3c3af335c487c2b2181468b8666ed3fe;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bb217fa29c9df711786c1b6b2439b026f5f8b3a4f06fc872be1bf651b77246df55ae284ac2c7bd12;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h33cec544a5f50119636aebb1e99bda903f5c07064b29c9fcaab1c43f5a5b45f128414a6b3cedf8dd8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc404c38bbccc2cddc9d992978ff5da00ce0fbab898f2053bea8ba0f7cb148ab2f1e9cd7af5a8c379;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h133b8a7b3ef4911c4bdbbac47612a184568a52a50311b5cfb7d0a01e5f51b35173196b966d6416864;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3881fd5f5777e94fcc440d65d3edeb85848aacc5811316e34da7fa1fd85faa16f8eeed90f10e21da7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf415585dd8ce11fa3c307a38b96f5c36a37163ed1791d919dfc404b52ccd15659536468b00a7e27e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h169490edd5335362ad917ff77c1701c46cd9f9432de94bc796b6733766a7bcfa9cadc37acdb6b50b8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b9aef8c7966b47411699a25c76feb7693d75753ccdd42e393f53846e42546a38b84e39e8bbd47a14;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13cdbb038cbee5b830f3363a2846c49999da62efc12e855160ecd94c16e0624791dde2ad66cff2b0b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa10b12e6fed38a63ab8c67461f3d6d80e14232546d61a746f594fca61d4bdaf1372da8365616192e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca3e3b54e2cfed273b28561c88cac5588f1c6ddbaefeeeff3e9d783ce403e201a83f7841ceee683f4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93f90111e548d102e1071c3b1f315439d6b7f91d955171798d3f3ff2c877f49a8aee195c7c3443e8b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf682449fda342632f5370745b527db33798a9b84e0977a20d739d53e5194b1ff3a8a452f68ebdbf29;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0b525be1ab1524b111eb46fb764d556e6cb3d48c8614461e571cd25dbd3adbfbe7beed8b42333175;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0f592d27fdea9bf9d52f8f3fc2555a78b50bce09c44c6cc9aa4eed52ab9e771fee0eb73c7f71e3a8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b03ee69c67e88621ac2b4738c7e4018638eb11b7f573a6e930b9d4aacab4fa0a18af2235c0aa14d8;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d538fa0f703a2dbc0bfb5ebb206d161dd32cccb4317270dc5201fb65e67baf8c9a160c4dc9a23dce;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10a4bf2047a5a6f352796cd8b0154e8149e7dd7cc44e36c79308bd39e0efb0254e25e80e038602bcb;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8967049a5b6d4dcc834ed66b7aded30d5cad6fb66fb9662d0f4357ed6bea42a4c110e7a5a3e800e24;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1974a89c15ea6f356b7336b8e37cd83ec7aff53e063a7afb1c4463ef2434c8a7acbac42ca9321c955;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h603f9a03be809a590f43ddc23f736d313669b8b3a066734cb5f33422d2aaca65235e60dee3446fb5c;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1aacc00b4865d20321524e8034cdf35debba9c992c05e1e7a3b42f74e6151c155e48da26cd6a3c03;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h286efce13669a71f83a3d917a8df77fcd7a21faec278999f9a664f60393a80be8303c15f695e97f9d;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6012b75e4a305e388c1a99da3f8391ab11589d25d316dac5904db30ffc3f70369e5efcb893fc776e5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4add2d1e7940bd5fcf2e538f677e14ccc27a7b6de8dcfc52519f4a1ae13e484c8e817a012c048be2;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h476df1d1a4196cac6d4243591ba922fc2ff23166135d74f8072e2687c2ab04a14f3c209ea7957436a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48b3b0a2d34d69fca1cf53c004eb4d0c0045fc6ef7fd205b30293b01ae40c3ec0611ec13363acd674;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83101154b4bb6653fd16d236c0ec5107e80920f14aeef4024b0e3530ef13a59d575d44ad3dacae562;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc7c97f425b6f92123abc70b0bbaafe242f3d22f8b89d34644eea44bc16dcb113dbe2d47d298a08c4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha736e18bccfb33326a3a3c218b1d4d458b8655167ccccfa37f0635208c6d2fbbe2ea5c4f2af1c8695;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae4fe279e417dc0b4afefc45fa3d37da5e8539bba7f21d47b5b66df2a85bdedf44491ce14d281b313;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ec5ece0925623cbe0932eac245631ea2da821c0c0739ddf35498163d20d3f21f7fa397ba9a98fb90;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1461b288735658a5425629ac0cff3e7cd25385857160301621a2bbe696cce30d7f9bc4677e29aeafd;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he784dca008f7457f81ca05f3a7ed267fdf748c4f1939e82bd723758ae75717078e78999433289081;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h756059a789994ed74ada7eca0208cdc1a577794c3e8c898ae1b72e28effb4855f06cb2b605c574481;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h458d29221ab979c1fd641cfd7cb3d10bf9782999017c4d87d3827417d6ead61f8518c5c4b56a478e3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd68acc76ab546ed7856fc3ddf1fb2d148b1cad651aec478f48c7e804a50ce2dea7ab8dbc4aa391a8e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4d9abd028753e635faa8525f48396f275357b91e160c697c2631716b3f6239e87c44fea7f3d1d7f1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11f0194e1a076302d73a21ad49bdaca4416775ccd25112c9dcc5d0723bbdf70ba17cc6d3b0111d10e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32faf663e069c9c1bff63a538fd92038d44c47ee172a6422a5e8fd4d63d1b83bd1ea094c64404813;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e857086a71ea6793efd705c759faa4c333faaefbbfee4cc76bc30201f0d4dab5ce87ea9f074d736b;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0aef074b0492e52b42ec5b63fc252017ec86e28d72f1b92eee99aae14bcb7bf67437ae9a73a0ce45;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c71d8f270f4390a2ddea5c1b9285051420a93dcf3e4040a8a906e274892e1b0f2c20958a6fd1d237;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h161c68f581798c19a076f32e3afe9b6060093c4bcc300bc52cbf6dbe5d8326f1e96b47cea0a8225d1;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4adb9cfeb723daff603926e32285aef11957d7e13832db19f025d222a8c94e7df7eeac7c1065ccf0;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2942c3ee20970dc20e5727cdb0b459b8de89cc01b0f53196a557dcfbbf33d5246f4f573b34627b708;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93f56a34f11df3b88e2a7105187ad9fb4e7fa3785aea342f9ad670ede71d49de0ce3f0ae2cae9057e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d924c2367b62643b04357d4eda84dbf28d7109d4ae7ee3f714d5b4b1d7f15205b453cf7ab33be263;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4ded57e7d2b496c51b5e797e96bc33fe7947c50e19ee53b63ab5752078cb570930fca50a138d526e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68651c09349b0025ec16eaf0322691691e218bf1a4d57e1a03d678b5e7ec9b6a83a2487f48b5b1bf4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75957a5e719d5d8931f2ddfc456028389a0f0e03f2dbb6a3990f82ce42eabaeaa5543a48152dfcaa7;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7548167cce5673a18f752920ea3d9320b9507601215a0d35218b00580b38ec506a033a00c7da348d5;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f1592d133f5c9526b4bfe9bee39874683193deb87c2cf44481df33faabde82a84188260a647f982e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97ed388a42e4bccca00f702465b26cf78904989b4174f12cd7c6dfcc1392461384d3640a7640dcb3;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3f3aeca040460b8ef922768118cd25b5751aa6b003da798f9305e6350fdec8541a8bbcaa04e61bc4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7c8856e7ad715830d5e0c51b70681a7347da3700e00ece884ac3239abd7eacd4d2d7da45f722d5af;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heace750e80b5c84c59676e42bc13ebe3529f847e5aa09ebc2895016439ae5fd949fae6658a558f82a;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f93d7a76b6d6d73439919bf0a1127fbcfc7f27b4cc95ad5490721c32f4395670395f822e53c6d3f6;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52e1979274ad436cebc8abc51683da9fa5dfd0d36ac8024a44e7dab3a54e5163f088f6568cc1e3f61;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5584638897bd60c0660ffd236811f3f220cbef3f809e283c80e312cae6490e105752ddf5a12f77b7e;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6de487247f2c291c505ba390c571911a101a9b4595615688e9c83aca2248edeec661c196174265167;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cc975896b9d8aa07ed7de26be9d980a1a3ca3a708dea0ea17fdbe70497b3620448cfeed950d770cc;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3184bd2966aec8e5b2d6470df6abbc77fd51aa3e23a9932947b987e72ef90222810e96a01df410e4;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96d7cbb39e846b382da5ffb9f76e9bb5f8efa22e37fcf296a961918b6d0c78a312a34a1e25e929068;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65a0e9d29087f0a5ae61d0f44c1be3f518996e3a39350c56f7c1741b3a1924f9ea84b4fd8b9e42101;
        #1
        {src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9755c3ca0b96ea61d2421ccca26d4d7c1e2c25000ba4324fc19175281b43163f41c103a6ae5f0203e;
        #1
        $finish();
    end
endmodule
