module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [15:0] src54;
    reg [15:0] src55;
    reg [15:0] src56;
    reg [15:0] src57;
    reg [15:0] src58;
    reg [15:0] src59;
    reg [15:0] src60;
    reg [15:0] src61;
    reg [15:0] src62;
    reg [15:0] src63;
    compressor_CLA16_64 compressor_CLA16_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67));
    initial begin
        src0 <= 16'h0;
        src1 <= 16'h0;
        src2 <= 16'h0;
        src3 <= 16'h0;
        src4 <= 16'h0;
        src5 <= 16'h0;
        src6 <= 16'h0;
        src7 <= 16'h0;
        src8 <= 16'h0;
        src9 <= 16'h0;
        src10 <= 16'h0;
        src11 <= 16'h0;
        src12 <= 16'h0;
        src13 <= 16'h0;
        src14 <= 16'h0;
        src15 <= 16'h0;
        src16 <= 16'h0;
        src17 <= 16'h0;
        src18 <= 16'h0;
        src19 <= 16'h0;
        src20 <= 16'h0;
        src21 <= 16'h0;
        src22 <= 16'h0;
        src23 <= 16'h0;
        src24 <= 16'h0;
        src25 <= 16'h0;
        src26 <= 16'h0;
        src27 <= 16'h0;
        src28 <= 16'h0;
        src29 <= 16'h0;
        src30 <= 16'h0;
        src31 <= 16'h0;
        src32 <= 16'h0;
        src33 <= 16'h0;
        src34 <= 16'h0;
        src35 <= 16'h0;
        src36 <= 16'h0;
        src37 <= 16'h0;
        src38 <= 16'h0;
        src39 <= 16'h0;
        src40 <= 16'h0;
        src41 <= 16'h0;
        src42 <= 16'h0;
        src43 <= 16'h0;
        src44 <= 16'h0;
        src45 <= 16'h0;
        src46 <= 16'h0;
        src47 <= 16'h0;
        src48 <= 16'h0;
        src49 <= 16'h0;
        src50 <= 16'h0;
        src51 <= 16'h0;
        src52 <= 16'h0;
        src53 <= 16'h0;
        src54 <= 16'h0;
        src55 <= 16'h0;
        src56 <= 16'h0;
        src57 <= 16'h0;
        src58 <= 16'h0;
        src59 <= 16'h0;
        src60 <= 16'h0;
        src61 <= 16'h0;
        src62 <= 16'h0;
        src63 <= 16'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA16_64(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    input [15:0]src16,
    input [15:0]src17,
    input [15:0]src18,
    input [15:0]src19,
    input [15:0]src20,
    input [15:0]src21,
    input [15:0]src22,
    input [15:0]src23,
    input [15:0]src24,
    input [15:0]src25,
    input [15:0]src26,
    input [15:0]src27,
    input [15:0]src28,
    input [15:0]src29,
    input [15:0]src30,
    input [15:0]src31,
    input [15:0]src32,
    input [15:0]src33,
    input [15:0]src34,
    input [15:0]src35,
    input [15:0]src36,
    input [15:0]src37,
    input [15:0]src38,
    input [15:0]src39,
    input [15:0]src40,
    input [15:0]src41,
    input [15:0]src42,
    input [15:0]src43,
    input [15:0]src44,
    input [15:0]src45,
    input [15:0]src46,
    input [15:0]src47,
    input [15:0]src48,
    input [15:0]src49,
    input [15:0]src50,
    input [15:0]src51,
    input [15:0]src52,
    input [15:0]src53,
    input [15:0]src54,
    input [15:0]src55,
    input [15:0]src56,
    input [15:0]src57,
    input [15:0]src58,
    input [15:0]src59,
    input [15:0]src60,
    input [15:0]src61,
    input [15:0]src62,
    input [15:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67);

    wire [1:0] comp_out0;
    wire [0:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [0:0] comp_out67;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], 1'h0, comp_out0[1]}),
        .dst({dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [15:0] src0,
      input wire [15:0] src1,
      input wire [15:0] src2,
      input wire [15:0] src3,
      input wire [15:0] src4,
      input wire [15:0] src5,
      input wire [15:0] src6,
      input wire [15:0] src7,
      input wire [15:0] src8,
      input wire [15:0] src9,
      input wire [15:0] src10,
      input wire [15:0] src11,
      input wire [15:0] src12,
      input wire [15:0] src13,
      input wire [15:0] src14,
      input wire [15:0] src15,
      input wire [15:0] src16,
      input wire [15:0] src17,
      input wire [15:0] src18,
      input wire [15:0] src19,
      input wire [15:0] src20,
      input wire [15:0] src21,
      input wire [15:0] src22,
      input wire [15:0] src23,
      input wire [15:0] src24,
      input wire [15:0] src25,
      input wire [15:0] src26,
      input wire [15:0] src27,
      input wire [15:0] src28,
      input wire [15:0] src29,
      input wire [15:0] src30,
      input wire [15:0] src31,
      input wire [15:0] src32,
      input wire [15:0] src33,
      input wire [15:0] src34,
      input wire [15:0] src35,
      input wire [15:0] src36,
      input wire [15:0] src37,
      input wire [15:0] src38,
      input wire [15:0] src39,
      input wire [15:0] src40,
      input wire [15:0] src41,
      input wire [15:0] src42,
      input wire [15:0] src43,
      input wire [15:0] src44,
      input wire [15:0] src45,
      input wire [15:0] src46,
      input wire [15:0] src47,
      input wire [15:0] src48,
      input wire [15:0] src49,
      input wire [15:0] src50,
      input wire [15:0] src51,
      input wire [15:0] src52,
      input wire [15:0] src53,
      input wire [15:0] src54,
      input wire [15:0] src55,
      input wire [15:0] src56,
      input wire [15:0] src57,
      input wire [15:0] src58,
      input wire [15:0] src59,
      input wire [15:0] src60,
      input wire [15:0] src61,
      input wire [15:0] src62,
      input wire [15:0] src63,
      output wire [1:0] dst0,
      output wire [0:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [0:0] dst67);

   wire [15:0] stage0_0;
   wire [15:0] stage0_1;
   wire [15:0] stage0_2;
   wire [15:0] stage0_3;
   wire [15:0] stage0_4;
   wire [15:0] stage0_5;
   wire [15:0] stage0_6;
   wire [15:0] stage0_7;
   wire [15:0] stage0_8;
   wire [15:0] stage0_9;
   wire [15:0] stage0_10;
   wire [15:0] stage0_11;
   wire [15:0] stage0_12;
   wire [15:0] stage0_13;
   wire [15:0] stage0_14;
   wire [15:0] stage0_15;
   wire [15:0] stage0_16;
   wire [15:0] stage0_17;
   wire [15:0] stage0_18;
   wire [15:0] stage0_19;
   wire [15:0] stage0_20;
   wire [15:0] stage0_21;
   wire [15:0] stage0_22;
   wire [15:0] stage0_23;
   wire [15:0] stage0_24;
   wire [15:0] stage0_25;
   wire [15:0] stage0_26;
   wire [15:0] stage0_27;
   wire [15:0] stage0_28;
   wire [15:0] stage0_29;
   wire [15:0] stage0_30;
   wire [15:0] stage0_31;
   wire [15:0] stage0_32;
   wire [15:0] stage0_33;
   wire [15:0] stage0_34;
   wire [15:0] stage0_35;
   wire [15:0] stage0_36;
   wire [15:0] stage0_37;
   wire [15:0] stage0_38;
   wire [15:0] stage0_39;
   wire [15:0] stage0_40;
   wire [15:0] stage0_41;
   wire [15:0] stage0_42;
   wire [15:0] stage0_43;
   wire [15:0] stage0_44;
   wire [15:0] stage0_45;
   wire [15:0] stage0_46;
   wire [15:0] stage0_47;
   wire [15:0] stage0_48;
   wire [15:0] stage0_49;
   wire [15:0] stage0_50;
   wire [15:0] stage0_51;
   wire [15:0] stage0_52;
   wire [15:0] stage0_53;
   wire [15:0] stage0_54;
   wire [15:0] stage0_55;
   wire [15:0] stage0_56;
   wire [15:0] stage0_57;
   wire [15:0] stage0_58;
   wire [15:0] stage0_59;
   wire [15:0] stage0_60;
   wire [15:0] stage0_61;
   wire [15:0] stage0_62;
   wire [15:0] stage0_63;
   wire [10:0] stage1_0;
   wire [6:0] stage1_1;
   wire [8:0] stage1_2;
   wire [6:0] stage1_3;
   wire [5:0] stage1_4;
   wire [7:0] stage1_5;
   wire [6:0] stage1_6;
   wire [5:0] stage1_7;
   wire [9:0] stage1_8;
   wire [5:0] stage1_9;
   wire [9:0] stage1_10;
   wire [6:0] stage1_11;
   wire [5:0] stage1_12;
   wire [9:0] stage1_13;
   wire [6:0] stage1_14;
   wire [6:0] stage1_15;
   wire [5:0] stage1_16;
   wire [14:0] stage1_17;
   wire [5:0] stage1_18;
   wire [11:0] stage1_19;
   wire [7:0] stage1_20;
   wire [5:0] stage1_21;
   wire [6:0] stage1_22;
   wire [5:0] stage1_23;
   wire [7:0] stage1_24;
   wire [6:0] stage1_25;
   wire [8:0] stage1_26;
   wire [6:0] stage1_27;
   wire [5:0] stage1_28;
   wire [6:0] stage1_29;
   wire [9:0] stage1_30;
   wire [7:0] stage1_31;
   wire [8:0] stage1_32;
   wire [8:0] stage1_33;
   wire [5:0] stage1_34;
   wire [7:0] stage1_35;
   wire [6:0] stage1_36;
   wire [8:0] stage1_37;
   wire [5:0] stage1_38;
   wire [5:0] stage1_39;
   wire [6:0] stage1_40;
   wire [9:0] stage1_41;
   wire [6:0] stage1_42;
   wire [5:0] stage1_43;
   wire [7:0] stage1_44;
   wire [6:0] stage1_45;
   wire [5:0] stage1_46;
   wire [7:0] stage1_47;
   wire [7:0] stage1_48;
   wire [6:0] stage1_49;
   wire [6:0] stage1_50;
   wire [8:0] stage1_51;
   wire [5:0] stage1_52;
   wire [13:0] stage1_53;
   wire [5:0] stage1_54;
   wire [5:0] stage1_55;
   wire [6:0] stage1_56;
   wire [9:0] stage1_57;
   wire [7:0] stage1_58;
   wire [7:0] stage1_59;
   wire [6:0] stage1_60;
   wire [5:0] stage1_61;
   wire [6:0] stage1_62;
   wire [13:0] stage1_63;
   wire [3:0] stage1_64;
   wire [0:0] stage1_65;
   wire [5:0] stage2_0;
   wire [2:0] stage2_1;
   wire [4:0] stage2_2;
   wire [2:0] stage2_3;
   wire [2:0] stage2_4;
   wire [4:0] stage2_5;
   wire [2:0] stage2_6;
   wire [1:0] stage2_7;
   wire [5:0] stage2_8;
   wire [2:0] stage2_9;
   wire [7:0] stage2_10;
   wire [1:0] stage2_11;
   wire [1:0] stage2_12;
   wire [6:0] stage2_13;
   wire [3:0] stage2_14;
   wire [2:0] stage2_15;
   wire [1:0] stage2_16;
   wire [6:0] stage2_17;
   wire [4:0] stage2_18;
   wire [2:0] stage2_19;
   wire [4:0] stage2_20;
   wire [4:0] stage2_21;
   wire [2:0] stage2_22;
   wire [1:0] stage2_23;
   wire [5:0] stage2_24;
   wire [2:0] stage2_25;
   wire [6:0] stage2_26;
   wire [1:0] stage2_27;
   wire [1:0] stage2_28;
   wire [2:0] stage2_29;
   wire [3:0] stage2_30;
   wire [3:0] stage2_31;
   wire [5:0] stage2_32;
   wire [2:0] stage2_33;
   wire [2:0] stage2_34;
   wire [3:0] stage2_35;
   wire [2:0] stage2_36;
   wire [5:0] stage2_37;
   wire [5:0] stage2_38;
   wire [1:0] stage2_39;
   wire [1:0] stage2_40;
   wire [6:0] stage2_41;
   wire [2:0] stage2_42;
   wire [1:0] stage2_43;
   wire [5:0] stage2_44;
   wire [2:0] stage2_45;
   wire [3:0] stage2_46;
   wire [1:0] stage2_47;
   wire [2:0] stage2_48;
   wire [6:0] stage2_49;
   wire [3:0] stage2_50;
   wire [2:0] stage2_51;
   wire [5:0] stage2_52;
   wire [4:0] stage2_53;
   wire [2:0] stage2_54;
   wire [3:0] stage2_55;
   wire [1:0] stage2_56;
   wire [6:0] stage2_57;
   wire [4:0] stage2_58;
   wire [2:0] stage2_59;
   wire [3:0] stage2_60;
   wire [1:0] stage2_61;
   wire [2:0] stage2_62;
   wire [9:0] stage2_63;
   wire [3:0] stage2_64;
   wire [1:0] stage2_65;
   wire [0:0] stage2_66;
   wire [1:0] stage3_0;
   wire [0:0] stage3_1;
   wire [1:0] stage3_2;
   wire [1:0] stage3_3;
   wire [1:0] stage3_4;
   wire [1:0] stage3_5;
   wire [1:0] stage3_6;
   wire [1:0] stage3_7;
   wire [1:0] stage3_8;
   wire [1:0] stage3_9;
   wire [1:0] stage3_10;
   wire [1:0] stage3_11;
   wire [1:0] stage3_12;
   wire [1:0] stage3_13;
   wire [1:0] stage3_14;
   wire [1:0] stage3_15;
   wire [1:0] stage3_16;
   wire [1:0] stage3_17;
   wire [1:0] stage3_18;
   wire [1:0] stage3_19;
   wire [1:0] stage3_20;
   wire [1:0] stage3_21;
   wire [1:0] stage3_22;
   wire [1:0] stage3_23;
   wire [1:0] stage3_24;
   wire [1:0] stage3_25;
   wire [1:0] stage3_26;
   wire [1:0] stage3_27;
   wire [1:0] stage3_28;
   wire [1:0] stage3_29;
   wire [1:0] stage3_30;
   wire [1:0] stage3_31;
   wire [1:0] stage3_32;
   wire [1:0] stage3_33;
   wire [1:0] stage3_34;
   wire [1:0] stage3_35;
   wire [1:0] stage3_36;
   wire [1:0] stage3_37;
   wire [1:0] stage3_38;
   wire [1:0] stage3_39;
   wire [1:0] stage3_40;
   wire [1:0] stage3_41;
   wire [1:0] stage3_42;
   wire [1:0] stage3_43;
   wire [1:0] stage3_44;
   wire [1:0] stage3_45;
   wire [1:0] stage3_46;
   wire [1:0] stage3_47;
   wire [1:0] stage3_48;
   wire [1:0] stage3_49;
   wire [1:0] stage3_50;
   wire [1:0] stage3_51;
   wire [1:0] stage3_52;
   wire [1:0] stage3_53;
   wire [1:0] stage3_54;
   wire [1:0] stage3_55;
   wire [1:0] stage3_56;
   wire [1:0] stage3_57;
   wire [1:0] stage3_58;
   wire [1:0] stage3_59;
   wire [1:0] stage3_60;
   wire [1:0] stage3_61;
   wire [1:0] stage3_62;
   wire [1:0] stage3_63;
   wire [1:0] stage3_64;
   wire [1:0] stage3_65;
   wire [1:0] stage3_66;
   wire [0:0] stage3_67;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage3_0;
   assign dst1 = stage3_1;
   assign dst2 = stage3_2;
   assign dst3 = stage3_3;
   assign dst4 = stage3_4;
   assign dst5 = stage3_5;
   assign dst6 = stage3_6;
   assign dst7 = stage3_7;
   assign dst8 = stage3_8;
   assign dst9 = stage3_9;
   assign dst10 = stage3_10;
   assign dst11 = stage3_11;
   assign dst12 = stage3_12;
   assign dst13 = stage3_13;
   assign dst14 = stage3_14;
   assign dst15 = stage3_15;
   assign dst16 = stage3_16;
   assign dst17 = stage3_17;
   assign dst18 = stage3_18;
   assign dst19 = stage3_19;
   assign dst20 = stage3_20;
   assign dst21 = stage3_21;
   assign dst22 = stage3_22;
   assign dst23 = stage3_23;
   assign dst24 = stage3_24;
   assign dst25 = stage3_25;
   assign dst26 = stage3_26;
   assign dst27 = stage3_27;
   assign dst28 = stage3_28;
   assign dst29 = stage3_29;
   assign dst30 = stage3_30;
   assign dst31 = stage3_31;
   assign dst32 = stage3_32;
   assign dst33 = stage3_33;
   assign dst34 = stage3_34;
   assign dst35 = stage3_35;
   assign dst36 = stage3_36;
   assign dst37 = stage3_37;
   assign dst38 = stage3_38;
   assign dst39 = stage3_39;
   assign dst40 = stage3_40;
   assign dst41 = stage3_41;
   assign dst42 = stage3_42;
   assign dst43 = stage3_43;
   assign dst44 = stage3_44;
   assign dst45 = stage3_45;
   assign dst46 = stage3_46;
   assign dst47 = stage3_47;
   assign dst48 = stage3_48;
   assign dst49 = stage3_49;
   assign dst50 = stage3_50;
   assign dst51 = stage3_51;
   assign dst52 = stage3_52;
   assign dst53 = stage3_53;
   assign dst54 = stage3_54;
   assign dst55 = stage3_55;
   assign dst56 = stage3_56;
   assign dst57 = stage3_57;
   assign dst58 = stage3_58;
   assign dst59 = stage3_59;
   assign dst60 = stage3_60;
   assign dst61 = stage3_61;
   assign dst62 = stage3_62;
   assign dst63 = stage3_63;
   assign dst64 = stage3_64;
   assign dst65 = stage3_65;
   assign dst66 = stage3_66;
   assign dst67 = stage3_67;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1]}
   );
   gpc606_5 gpc2 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2]}
   );
   gpc615_5 gpc3 (
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage0_3[12]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[2],stage1_4[3],stage1_3[3],stage1_2[3]}
   );
   gpc615_5 gpc4 (
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10]},
      {stage0_5[0]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[0],stage1_6[1],stage1_5[3],stage1_4[4]}
   );
   gpc615_5 gpc5 (
      {stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15]},
      {stage0_5[1]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[1],stage1_6[2],stage1_5[4],stage1_4[5]}
   );
   gpc207_4 gpc6 (
      {stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7], stage0_5[8]},
      {stage0_7[0], stage0_7[1]},
      {stage1_8[2],stage1_7[2],stage1_6[3],stage1_5[5]}
   );
   gpc606_5 gpc7 (
      {stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14]},
      {stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6], stage0_7[7]},
      {stage1_9[0],stage1_8[3],stage1_7[3],stage1_6[4],stage1_5[6]}
   );
   gpc1343_5 gpc8 (
      {stage0_6[12], stage0_6[13], stage0_6[14]},
      {stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage0_8[0], stage0_8[1], stage0_8[2]},
      {stage0_9[0]},
      {stage1_10[0],stage1_9[1],stage1_8[4],stage1_7[4],stage1_6[5]}
   );
   gpc1343_5 gpc9 (
      {stage0_6[15], 1'b0, 1'b0},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15]},
      {stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage0_9[1]},
      {stage1_10[1],stage1_9[2],stage1_8[5],stage1_7[5],stage1_6[6]}
   );
   gpc117_4 gpc10 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12]},
      {stage0_9[2]},
      {stage0_10[0]},
      {stage1_11[0],stage1_10[2],stage1_9[3],stage1_8[6]}
   );
   gpc207_4 gpc11 (
      {stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9]},
      {stage0_11[0], stage0_11[1]},
      {stage1_12[0],stage1_11[1],stage1_10[3],stage1_9[4]}
   );
   gpc606_5 gpc12 (
      {stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15]},
      {stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6], stage0_11[7]},
      {stage1_13[0],stage1_12[1],stage1_11[2],stage1_10[4],stage1_9[5]}
   );
   gpc117_4 gpc13 (
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7]},
      {stage0_11[8]},
      {stage0_12[0]},
      {stage1_13[1],stage1_12[2],stage1_11[3],stage1_10[5]}
   );
   gpc615_5 gpc14 (
      {stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11], stage0_10[12]},
      {stage0_11[9]},
      {stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5], stage0_12[6]},
      {stage1_14[0],stage1_13[2],stage1_12[3],stage1_11[4],stage1_10[6]}
   );
   gpc135_4 gpc15 (
      {stage0_11[10], stage0_11[11], stage0_11[12], stage0_11[13], stage0_11[14]},
      {stage0_12[7], stage0_12[8], stage0_12[9]},
      {stage0_13[0]},
      {stage1_14[1],stage1_13[3],stage1_12[4],stage1_11[5]}
   );
   gpc606_5 gpc16 (
      {stage0_12[10], stage0_12[11], stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[0],stage1_14[2],stage1_13[4],stage1_12[5]}
   );
   gpc606_5 gpc17 (
      {stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5], stage0_13[6]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[1],stage1_15[1],stage1_14[3],stage1_13[5]}
   );
   gpc606_5 gpc18 (
      {stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11], stage0_13[12]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[2],stage1_15[2],stage1_14[4],stage1_13[6]}
   );
   gpc615_5 gpc19 (
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10]},
      {stage0_15[12]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[2],stage1_16[3],stage1_15[3],stage1_14[5]}
   );
   gpc615_5 gpc20 (
      {stage0_14[11], stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15]},
      {stage0_15[13]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[3],stage1_16[4],stage1_15[4],stage1_14[6]}
   );
   gpc615_5 gpc21 (
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], 1'b0},
      {stage0_17[0]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[0],stage1_18[2],stage1_17[4],stage1_16[5]}
   );
   gpc606_5 gpc22 (
      {stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5], stage0_17[6]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[1],stage1_19[1],stage1_18[3],stage1_17[5]}
   );
   gpc615_5 gpc23 (
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10]},
      {stage0_19[6]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[1],stage1_20[2],stage1_19[2],stage1_18[4]}
   );
   gpc615_5 gpc24 (
      {stage0_18[11], stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15]},
      {stage0_19[7]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[2],stage1_20[3],stage1_19[3],stage1_18[5]}
   );
   gpc1343_5 gpc25 (
      {stage0_21[0], stage0_21[1], stage0_21[2]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3]},
      {stage0_23[0], stage0_23[1], stage0_23[2]},
      {stage0_24[0]},
      {stage1_25[0],stage1_24[0],stage1_23[0],stage1_22[2],stage1_21[3]}
   );
   gpc117_4 gpc26 (
      {stage0_21[3], stage0_21[4], stage0_21[5], stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9]},
      {stage0_22[4]},
      {stage0_23[3]},
      {stage1_24[1],stage1_23[1],stage1_22[3],stage1_21[4]}
   );
   gpc606_5 gpc27 (
      {stage0_21[10], stage0_21[11], stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15]},
      {stage0_23[4], stage0_23[5], stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9]},
      {stage1_25[1],stage1_24[2],stage1_23[2],stage1_22[4],stage1_21[5]}
   );
   gpc606_5 gpc28 (
      {stage0_22[5], stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10]},
      {stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5], stage0_24[6]},
      {stage1_26[0],stage1_25[2],stage1_24[3],stage1_23[3],stage1_22[5]}
   );
   gpc615_5 gpc29 (
      {stage0_22[11], stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15]},
      {stage0_23[10]},
      {stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11], stage0_24[12]},
      {stage1_26[1],stage1_25[3],stage1_24[4],stage1_23[4],stage1_22[6]}
   );
   gpc615_5 gpc30 (
      {stage0_23[11], stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15]},
      {stage0_24[13]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[2],stage1_25[4],stage1_24[5],stage1_23[5]}
   );
   gpc15_3 gpc31 (
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10]},
      {stage0_26[0]},
      {stage1_27[1],stage1_26[3],stage1_25[5]}
   );
   gpc615_5 gpc32 (
      {stage0_25[11], stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15]},
      {stage0_26[1]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[0],stage1_27[2],stage1_26[4],stage1_25[6]}
   );
   gpc606_5 gpc33 (
      {stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5], stage0_26[6], stage0_26[7]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[1],stage1_28[1],stage1_27[3],stage1_26[5]}
   );
   gpc606_5 gpc34 (
      {stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11], stage0_26[12], stage0_26[13]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[2],stage1_28[2],stage1_27[4],stage1_26[6]}
   );
   gpc615_5 gpc35 (
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10]},
      {stage0_28[12]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[2],stage1_29[3],stage1_28[3],stage1_27[5]}
   );
   gpc615_5 gpc36 (
      {stage0_27[11], stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15]},
      {stage0_28[13]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[3],stage1_29[4],stage1_28[4],stage1_27[6]}
   );
   gpc615_5 gpc37 (
      {stage0_28[14], stage0_28[15], 1'b0, 1'b0, 1'b0},
      {stage0_29[12]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[2],stage1_30[4],stage1_29[5],stage1_28[5]}
   );
   gpc1163_5 gpc38 (
      {stage0_29[13], stage0_29[14], stage0_29[15]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage0_31[0]},
      {stage0_32[0]},
      {stage1_33[0],stage1_32[1],stage1_31[3],stage1_30[5],stage1_29[6]}
   );
   gpc117_4 gpc39 (
      {stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5], stage0_31[6], stage0_31[7]},
      {stage0_32[1]},
      {stage0_33[0]},
      {stage1_34[0],stage1_33[1],stage1_32[2],stage1_31[4]}
   );
   gpc606_5 gpc40 (
      {stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11], stage0_31[12], stage0_31[13]},
      {stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5], stage0_33[6]},
      {stage1_35[0],stage1_34[1],stage1_33[2],stage1_32[3],stage1_31[5]}
   );
   gpc1406_5 gpc41 (
      {stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5], stage0_32[6], stage0_32[7]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3]},
      {stage0_35[0]},
      {stage1_36[0],stage1_35[1],stage1_34[2],stage1_33[3],stage1_32[4]}
   );
   gpc615_5 gpc42 (
      {stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11], stage0_32[12]},
      {stage0_33[7]},
      {stage0_34[4], stage0_34[5], stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9]},
      {stage1_36[1],stage1_35[2],stage1_34[3],stage1_33[4],stage1_32[5]}
   );
   gpc615_5 gpc43 (
      {stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11], stage0_33[12]},
      {stage0_34[10]},
      {stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5], stage0_35[6]},
      {stage1_37[0],stage1_36[2],stage1_35[3],stage1_34[4],stage1_33[5]}
   );
   gpc615_5 gpc44 (
      {stage0_34[11], stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15]},
      {stage0_35[7]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[1],stage1_36[3],stage1_35[4],stage1_34[5]}
   );
   gpc606_5 gpc45 (
      {stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11], stage0_35[12], stage0_35[13]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[1],stage1_37[2],stage1_36[4],stage1_35[5]}
   );
   gpc615_5 gpc46 (
      {stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10]},
      {stage0_37[6]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[1],stage1_38[2],stage1_37[3],stage1_36[5]}
   );
   gpc615_5 gpc47 (
      {stage0_36[11], stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15]},
      {stage0_37[7]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[2],stage1_38[3],stage1_37[4],stage1_36[6]}
   );
   gpc615_5 gpc48 (
      {stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11], stage0_37[12]},
      {stage0_38[12]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[2],stage1_39[3],stage1_38[4],stage1_37[5]}
   );
   gpc1163_5 gpc49 (
      {stage0_38[13], stage0_38[14], stage0_38[15]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage0_40[0]},
      {stage0_41[0]},
      {stage1_42[0],stage1_41[1],stage1_40[3],stage1_39[4],stage1_38[5]}
   );
   gpc135_4 gpc50 (
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], 1'b0},
      {stage0_40[1], stage0_40[2], stage0_40[3]},
      {stage0_41[1]},
      {stage1_42[1],stage1_41[2],stage1_40[4],stage1_39[5]}
   );
   gpc606_5 gpc51 (
      {stage0_40[4], stage0_40[5], stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[0],stage1_42[2],stage1_41[3],stage1_40[5]}
   );
   gpc606_5 gpc52 (
      {stage0_40[10], stage0_40[11], stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[1],stage1_42[3],stage1_41[4],stage1_40[6]}
   );
   gpc135_4 gpc53 (
      {stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5], stage0_41[6]},
      {stage0_42[12], stage0_42[13], stage0_42[14]},
      {stage0_43[0]},
      {stage1_44[2],stage1_43[2],stage1_42[4],stage1_41[5]}
   );
   gpc606_5 gpc54 (
      {stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11], stage0_41[12]},
      {stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5], stage0_43[6]},
      {stage1_45[0],stage1_44[3],stage1_43[3],stage1_42[5],stage1_41[6]}
   );
   gpc1406_5 gpc55 (
      {stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11], stage0_43[12]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3]},
      {stage0_46[0]},
      {stage1_47[0],stage1_46[0],stage1_45[1],stage1_44[4],stage1_43[4]}
   );
   gpc1163_5 gpc56 (
      {stage0_43[13], stage0_43[14], stage0_43[15]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage0_45[4]},
      {stage0_46[1]},
      {stage1_47[1],stage1_46[1],stage1_45[2],stage1_44[5],stage1_43[5]}
   );
   gpc615_5 gpc57 (
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10]},
      {stage0_45[5]},
      {stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5], stage0_46[6], stage0_46[7]},
      {stage1_48[0],stage1_47[2],stage1_46[2],stage1_45[3],stage1_44[6]}
   );
   gpc615_5 gpc58 (
      {stage0_44[11], stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15]},
      {stage0_45[6]},
      {stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11], stage0_46[12], stage0_46[13]},
      {stage1_48[1],stage1_47[3],stage1_46[3],stage1_45[4],stage1_44[7]}
   );
   gpc615_5 gpc59 (
      {stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage0_46[14]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[2],stage1_47[4],stage1_46[4],stage1_45[5]}
   );
   gpc615_5 gpc60 (
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], 1'b0},
      {stage0_46[15]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[3],stage1_47[5],stage1_46[5],stage1_45[6]}
   );
   gpc623_5 gpc61 (
      {stage0_47[12], stage0_47[13], stage0_47[14]},
      {stage0_48[0], stage0_48[1]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[0],stage1_49[2],stage1_48[4],stage1_47[6]}
   );
   gpc207_4 gpc62 (
      {stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5], stage0_48[6], stage0_48[7], stage0_48[8]},
      {stage0_50[0], stage0_50[1]},
      {stage1_51[1],stage1_50[1],stage1_49[3],stage1_48[5]}
   );
   gpc606_5 gpc63 (
      {stage0_48[9], stage0_48[10], stage0_48[11], stage0_48[12], stage0_48[13], stage0_48[14]},
      {stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5], stage0_50[6], stage0_50[7]},
      {stage1_52[0],stage1_51[2],stage1_50[2],stage1_49[4],stage1_48[6]}
   );
   gpc615_5 gpc64 (
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10]},
      {stage0_50[8]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[1],stage1_51[3],stage1_50[3],stage1_49[5]}
   );
   gpc615_5 gpc65 (
      {stage0_49[11], stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15]},
      {stage0_50[9]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[2],stage1_51[4],stage1_50[4],stage1_49[6]}
   );
   gpc615_5 gpc66 (
      {stage0_50[10], stage0_50[11], stage0_50[12], stage0_50[13], stage0_50[14]},
      {stage0_51[12]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[2],stage1_52[3],stage1_51[5],stage1_50[5]}
   );
   gpc615_5 gpc67 (
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10]},
      {stage0_53[0]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[0],stage1_54[1],stage1_53[3],stage1_52[4]}
   );
   gpc615_5 gpc68 (
      {stage0_52[11], stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15]},
      {stage0_53[1]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[1],stage1_54[2],stage1_53[4],stage1_52[5]}
   );
   gpc606_5 gpc69 (
      {stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5], stage0_53[6], stage0_53[7]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[2],stage1_55[2],stage1_54[3],stage1_53[5]}
   );
   gpc1343_5 gpc70 (
      {stage0_54[12], stage0_54[13], stage0_54[14]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9]},
      {stage0_56[0], stage0_56[1], stage0_56[2]},
      {stage0_57[0]},
      {stage1_58[0],stage1_57[1],stage1_56[3],stage1_55[3],stage1_54[4]}
   );
   gpc615_5 gpc71 (
      {stage0_55[10], stage0_55[11], stage0_55[12], stage0_55[13], stage0_55[14]},
      {stage0_56[3]},
      {stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5], stage0_57[6]},
      {stage1_59[0],stage1_58[1],stage1_57[2],stage1_56[4],stage1_55[4]}
   );
   gpc606_5 gpc72 (
      {stage0_56[4], stage0_56[5], stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[1],stage1_58[2],stage1_57[3],stage1_56[5]}
   );
   gpc606_5 gpc73 (
      {stage0_56[10], stage0_56[11], stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[2],stage1_58[3],stage1_57[4],stage1_56[6]}
   );
   gpc615_5 gpc74 (
      {stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage0_58[12]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[2],stage1_59[3],stage1_58[4],stage1_57[5]}
   );
   gpc1343_5 gpc75 (
      {stage0_59[6], stage0_59[7], stage0_59[8]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3]},
      {stage0_61[0], stage0_61[1], stage0_61[2]},
      {stage0_62[0]},
      {stage1_63[0],stage1_62[0],stage1_61[1],stage1_60[3],stage1_59[4]}
   );
   gpc615_5 gpc76 (
      {stage0_59[9], stage0_59[10], stage0_59[11], stage0_59[12], stage0_59[13]},
      {stage0_60[4]},
      {stage0_61[3], stage0_61[4], stage0_61[5], stage0_61[6], stage0_61[7], stage0_61[8]},
      {stage1_63[1],stage1_62[1],stage1_61[2],stage1_60[4],stage1_59[5]}
   );
   gpc606_5 gpc77 (
      {stage0_60[5], stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10]},
      {stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5], stage0_62[6]},
      {stage1_64[0],stage1_63[2],stage1_62[2],stage1_61[3],stage1_60[5]}
   );
   gpc615_5 gpc78 (
      {stage0_60[11], stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15]},
      {stage0_61[9]},
      {stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11], stage0_62[12]},
      {stage1_64[1],stage1_63[3],stage1_62[3],stage1_61[4],stage1_60[6]}
   );
   gpc117_4 gpc79 (
      {stage0_61[10], stage0_61[11], stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15], 1'b0},
      {stage0_62[13]},
      {stage0_63[0]},
      {stage1_64[2],stage1_63[4],stage1_62[4],stage1_61[5]}
   );
   gpc7_3 gpc80 (
      {stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5], stage0_63[6], stage0_63[7]},
      {stage1_65[0],stage1_64[3],stage1_63[5]}
   );
   gpc1_1 gpc81 (
      {stage0_0[6]},
      {stage1_0[1]}
   );
   gpc1_1 gpc82 (
      {stage0_0[7]},
      {stage1_0[2]}
   );
   gpc1_1 gpc83 (
      {stage0_0[8]},
      {stage1_0[3]}
   );
   gpc1_1 gpc84 (
      {stage0_0[9]},
      {stage1_0[4]}
   );
   gpc1_1 gpc85 (
      {stage0_0[10]},
      {stage1_0[5]}
   );
   gpc1_1 gpc86 (
      {stage0_0[11]},
      {stage1_0[6]}
   );
   gpc1_1 gpc87 (
      {stage0_0[12]},
      {stage1_0[7]}
   );
   gpc1_1 gpc88 (
      {stage0_0[13]},
      {stage1_0[8]}
   );
   gpc1_1 gpc89 (
      {stage0_0[14]},
      {stage1_0[9]}
   );
   gpc1_1 gpc90 (
      {stage0_0[15]},
      {stage1_0[10]}
   );
   gpc1_1 gpc91 (
      {stage0_1[12]},
      {stage1_1[3]}
   );
   gpc1_1 gpc92 (
      {stage0_1[13]},
      {stage1_1[4]}
   );
   gpc1_1 gpc93 (
      {stage0_1[14]},
      {stage1_1[5]}
   );
   gpc1_1 gpc94 (
      {stage0_1[15]},
      {stage1_1[6]}
   );
   gpc1_1 gpc95 (
      {stage0_2[11]},
      {stage1_2[4]}
   );
   gpc1_1 gpc96 (
      {stage0_2[12]},
      {stage1_2[5]}
   );
   gpc1_1 gpc97 (
      {stage0_2[13]},
      {stage1_2[6]}
   );
   gpc1_1 gpc98 (
      {stage0_2[14]},
      {stage1_2[7]}
   );
   gpc1_1 gpc99 (
      {stage0_2[15]},
      {stage1_2[8]}
   );
   gpc1_1 gpc100 (
      {stage0_3[13]},
      {stage1_3[4]}
   );
   gpc1_1 gpc101 (
      {stage0_3[14]},
      {stage1_3[5]}
   );
   gpc1_1 gpc102 (
      {stage0_3[15]},
      {stage1_3[6]}
   );
   gpc1_1 gpc103 (
      {stage0_5[15]},
      {stage1_5[7]}
   );
   gpc1_1 gpc104 (
      {stage0_8[13]},
      {stage1_8[7]}
   );
   gpc1_1 gpc105 (
      {stage0_8[14]},
      {stage1_8[8]}
   );
   gpc1_1 gpc106 (
      {stage0_8[15]},
      {stage1_8[9]}
   );
   gpc1_1 gpc107 (
      {stage0_10[13]},
      {stage1_10[7]}
   );
   gpc1_1 gpc108 (
      {stage0_10[14]},
      {stage1_10[8]}
   );
   gpc1_1 gpc109 (
      {stage0_10[15]},
      {stage1_10[9]}
   );
   gpc1_1 gpc110 (
      {stage0_11[15]},
      {stage1_11[6]}
   );
   gpc1_1 gpc111 (
      {stage0_13[13]},
      {stage1_13[7]}
   );
   gpc1_1 gpc112 (
      {stage0_13[14]},
      {stage1_13[8]}
   );
   gpc1_1 gpc113 (
      {stage0_13[15]},
      {stage1_13[9]}
   );
   gpc1_1 gpc114 (
      {stage0_15[14]},
      {stage1_15[5]}
   );
   gpc1_1 gpc115 (
      {stage0_15[15]},
      {stage1_15[6]}
   );
   gpc1_1 gpc116 (
      {stage0_17[7]},
      {stage1_17[6]}
   );
   gpc1_1 gpc117 (
      {stage0_17[8]},
      {stage1_17[7]}
   );
   gpc1_1 gpc118 (
      {stage0_17[9]},
      {stage1_17[8]}
   );
   gpc1_1 gpc119 (
      {stage0_17[10]},
      {stage1_17[9]}
   );
   gpc1_1 gpc120 (
      {stage0_17[11]},
      {stage1_17[10]}
   );
   gpc1_1 gpc121 (
      {stage0_17[12]},
      {stage1_17[11]}
   );
   gpc1_1 gpc122 (
      {stage0_17[13]},
      {stage1_17[12]}
   );
   gpc1_1 gpc123 (
      {stage0_17[14]},
      {stage1_17[13]}
   );
   gpc1_1 gpc124 (
      {stage0_17[15]},
      {stage1_17[14]}
   );
   gpc1_1 gpc125 (
      {stage0_19[8]},
      {stage1_19[4]}
   );
   gpc1_1 gpc126 (
      {stage0_19[9]},
      {stage1_19[5]}
   );
   gpc1_1 gpc127 (
      {stage0_19[10]},
      {stage1_19[6]}
   );
   gpc1_1 gpc128 (
      {stage0_19[11]},
      {stage1_19[7]}
   );
   gpc1_1 gpc129 (
      {stage0_19[12]},
      {stage1_19[8]}
   );
   gpc1_1 gpc130 (
      {stage0_19[13]},
      {stage1_19[9]}
   );
   gpc1_1 gpc131 (
      {stage0_19[14]},
      {stage1_19[10]}
   );
   gpc1_1 gpc132 (
      {stage0_19[15]},
      {stage1_19[11]}
   );
   gpc1_1 gpc133 (
      {stage0_20[12]},
      {stage1_20[4]}
   );
   gpc1_1 gpc134 (
      {stage0_20[13]},
      {stage1_20[5]}
   );
   gpc1_1 gpc135 (
      {stage0_20[14]},
      {stage1_20[6]}
   );
   gpc1_1 gpc136 (
      {stage0_20[15]},
      {stage1_20[7]}
   );
   gpc1_1 gpc137 (
      {stage0_24[14]},
      {stage1_24[6]}
   );
   gpc1_1 gpc138 (
      {stage0_24[15]},
      {stage1_24[7]}
   );
   gpc1_1 gpc139 (
      {stage0_26[14]},
      {stage1_26[7]}
   );
   gpc1_1 gpc140 (
      {stage0_26[15]},
      {stage1_26[8]}
   );
   gpc1_1 gpc141 (
      {stage0_30[12]},
      {stage1_30[6]}
   );
   gpc1_1 gpc142 (
      {stage0_30[13]},
      {stage1_30[7]}
   );
   gpc1_1 gpc143 (
      {stage0_30[14]},
      {stage1_30[8]}
   );
   gpc1_1 gpc144 (
      {stage0_30[15]},
      {stage1_30[9]}
   );
   gpc1_1 gpc145 (
      {stage0_31[14]},
      {stage1_31[6]}
   );
   gpc1_1 gpc146 (
      {stage0_31[15]},
      {stage1_31[7]}
   );
   gpc1_1 gpc147 (
      {stage0_32[13]},
      {stage1_32[6]}
   );
   gpc1_1 gpc148 (
      {stage0_32[14]},
      {stage1_32[7]}
   );
   gpc1_1 gpc149 (
      {stage0_32[15]},
      {stage1_32[8]}
   );
   gpc1_1 gpc150 (
      {stage0_33[13]},
      {stage1_33[6]}
   );
   gpc1_1 gpc151 (
      {stage0_33[14]},
      {stage1_33[7]}
   );
   gpc1_1 gpc152 (
      {stage0_33[15]},
      {stage1_33[8]}
   );
   gpc1_1 gpc153 (
      {stage0_35[14]},
      {stage1_35[6]}
   );
   gpc1_1 gpc154 (
      {stage0_35[15]},
      {stage1_35[7]}
   );
   gpc1_1 gpc155 (
      {stage0_37[13]},
      {stage1_37[6]}
   );
   gpc1_1 gpc156 (
      {stage0_37[14]},
      {stage1_37[7]}
   );
   gpc1_1 gpc157 (
      {stage0_37[15]},
      {stage1_37[8]}
   );
   gpc1_1 gpc158 (
      {stage0_41[13]},
      {stage1_41[7]}
   );
   gpc1_1 gpc159 (
      {stage0_41[14]},
      {stage1_41[8]}
   );
   gpc1_1 gpc160 (
      {stage0_41[15]},
      {stage1_41[9]}
   );
   gpc1_1 gpc161 (
      {stage0_42[15]},
      {stage1_42[6]}
   );
   gpc1_1 gpc162 (
      {stage0_47[15]},
      {stage1_47[7]}
   );
   gpc1_1 gpc163 (
      {stage0_48[15]},
      {stage1_48[7]}
   );
   gpc1_1 gpc164 (
      {stage0_50[15]},
      {stage1_50[6]}
   );
   gpc1_1 gpc165 (
      {stage0_51[13]},
      {stage1_51[6]}
   );
   gpc1_1 gpc166 (
      {stage0_51[14]},
      {stage1_51[7]}
   );
   gpc1_1 gpc167 (
      {stage0_51[15]},
      {stage1_51[8]}
   );
   gpc1_1 gpc168 (
      {stage0_53[8]},
      {stage1_53[6]}
   );
   gpc1_1 gpc169 (
      {stage0_53[9]},
      {stage1_53[7]}
   );
   gpc1_1 gpc170 (
      {stage0_53[10]},
      {stage1_53[8]}
   );
   gpc1_1 gpc171 (
      {stage0_53[11]},
      {stage1_53[9]}
   );
   gpc1_1 gpc172 (
      {stage0_53[12]},
      {stage1_53[10]}
   );
   gpc1_1 gpc173 (
      {stage0_53[13]},
      {stage1_53[11]}
   );
   gpc1_1 gpc174 (
      {stage0_53[14]},
      {stage1_53[12]}
   );
   gpc1_1 gpc175 (
      {stage0_53[15]},
      {stage1_53[13]}
   );
   gpc1_1 gpc176 (
      {stage0_54[15]},
      {stage1_54[5]}
   );
   gpc1_1 gpc177 (
      {stage0_55[15]},
      {stage1_55[5]}
   );
   gpc1_1 gpc178 (
      {stage0_57[12]},
      {stage1_57[6]}
   );
   gpc1_1 gpc179 (
      {stage0_57[13]},
      {stage1_57[7]}
   );
   gpc1_1 gpc180 (
      {stage0_57[14]},
      {stage1_57[8]}
   );
   gpc1_1 gpc181 (
      {stage0_57[15]},
      {stage1_57[9]}
   );
   gpc1_1 gpc182 (
      {stage0_58[13]},
      {stage1_58[5]}
   );
   gpc1_1 gpc183 (
      {stage0_58[14]},
      {stage1_58[6]}
   );
   gpc1_1 gpc184 (
      {stage0_58[15]},
      {stage1_58[7]}
   );
   gpc1_1 gpc185 (
      {stage0_59[14]},
      {stage1_59[6]}
   );
   gpc1_1 gpc186 (
      {stage0_59[15]},
      {stage1_59[7]}
   );
   gpc1_1 gpc187 (
      {stage0_62[14]},
      {stage1_62[5]}
   );
   gpc1_1 gpc188 (
      {stage0_62[15]},
      {stage1_62[6]}
   );
   gpc1_1 gpc189 (
      {stage0_63[8]},
      {stage1_63[6]}
   );
   gpc1_1 gpc190 (
      {stage0_63[9]},
      {stage1_63[7]}
   );
   gpc1_1 gpc191 (
      {stage0_63[10]},
      {stage1_63[8]}
   );
   gpc1_1 gpc192 (
      {stage0_63[11]},
      {stage1_63[9]}
   );
   gpc1_1 gpc193 (
      {stage0_63[12]},
      {stage1_63[10]}
   );
   gpc1_1 gpc194 (
      {stage0_63[13]},
      {stage1_63[11]}
   );
   gpc1_1 gpc195 (
      {stage0_63[14]},
      {stage1_63[12]}
   );
   gpc1_1 gpc196 (
      {stage0_63[15]},
      {stage1_63[13]}
   );
   gpc606_5 gpc197 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc198 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1]}
   );
   gpc606_5 gpc199 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[1],stage2_4[2]}
   );
   gpc606_5 gpc200 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[2]}
   );
   gpc7_3 gpc201 (
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5], stage1_8[6]},
      {stage2_10[0],stage2_9[1],stage2_8[2]}
   );
   gpc606_5 gpc202 (
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[0],stage2_10[1],stage2_9[2]}
   );
   gpc615_5 gpc203 (
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4]},
      {stage1_11[6]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[1],stage2_11[1],stage2_10[2]}
   );
   gpc606_5 gpc204 (
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[0],stage2_14[1],stage2_13[2]}
   );
   gpc606_5 gpc205 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[1],stage2_16[1],stage2_15[1],stage2_14[2]}
   );
   gpc606_5 gpc206 (
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[0],stage2_19[0],stage2_18[1],stage2_17[2]}
   );
   gpc606_5 gpc207 (
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[1],stage2_19[1],stage2_18[2],stage2_17[3]}
   );
   gpc615_5 gpc208 (
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4]},
      {1'b0},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[2],stage2_20[2],stage2_19[2],stage2_18[3]}
   );
   gpc615_5 gpc209 (
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4]},
      {stage1_22[0]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[0],stage2_23[0],stage2_22[1],stage2_21[3]}
   );
   gpc1406_5 gpc210 (
      {stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5], stage1_22[6]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3]},
      {stage1_25[0]},
      {stage2_26[0],stage2_25[1],stage2_24[1],stage2_23[1],stage2_22[2]}
   );
   gpc606_5 gpc211 (
      {stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5], stage1_25[6]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[0],stage2_27[0],stage2_26[1],stage2_25[2]}
   );
   gpc615_5 gpc212 (
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4]},
      {stage1_27[6]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[1],stage2_28[1],stage2_27[1],stage2_26[2]}
   );
   gpc7_3 gpc213 (
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5], stage1_29[6]},
      {stage2_31[0],stage2_30[1],stage2_29[2]}
   );
   gpc7_3 gpc214 (
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5], stage1_30[6]},
      {stage2_32[0],stage2_31[1],stage2_30[2]}
   );
   gpc623_5 gpc215 (
      {stage1_30[7], stage1_30[8], stage1_30[9]},
      {stage1_31[0], stage1_31[1]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[0],stage2_32[1],stage2_31[2],stage2_30[3]}
   );
   gpc606_5 gpc216 (
      {stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5], stage1_31[6], stage1_31[7]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[1],stage2_33[1],stage2_32[2],stage2_31[3]}
   );
   gpc1163_5 gpc217 (
      {stage1_33[6], stage1_33[7], stage1_33[8]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage1_35[0]},
      {stage1_36[0]},
      {stage2_37[0],stage2_36[0],stage2_35[1],stage2_34[2],stage2_33[2]}
   );
   gpc606_5 gpc218 (
      {stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5], stage1_35[6]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[0],stage2_37[1],stage2_36[1],stage2_35[2]}
   );
   gpc7_3 gpc219 (
      {stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5], stage1_36[6], 1'b0},
      {stage2_38[1],stage2_37[2],stage2_36[2]}
   );
   gpc1163_5 gpc220 (
      {stage1_38[0], stage1_38[1], stage1_38[2]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage1_40[0]},
      {stage1_41[0]},
      {stage2_42[0],stage2_41[0],stage2_40[0],stage2_39[1],stage2_38[2]}
   );
   gpc606_5 gpc221 (
      {stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5], stage1_40[6]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[0],stage2_42[1],stage2_41[1],stage2_40[1]}
   );
   gpc615_5 gpc222 (
      {stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage1_42[6]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[1],stage2_43[1],stage2_42[2],stage2_41[2]}
   );
   gpc15_3 gpc223 (
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4]},
      {stage1_45[0]},
      {stage2_46[0],stage2_45[1],stage2_44[2]}
   );
   gpc606_5 gpc224 (
      {stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5], stage1_45[6]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[0],stage2_47[0],stage2_46[1],stage2_45[2]}
   );
   gpc1325_5 gpc225 (
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4]},
      {stage1_47[6], stage1_47[7]},
      {stage1_48[0], stage1_48[1], stage1_48[2]},
      {stage1_49[0]},
      {stage2_50[0],stage2_49[1],stage2_48[1],stage2_47[1],stage2_46[2]}
   );
   gpc7_3 gpc226 (
      {stage1_48[3], stage1_48[4], stage1_48[5], stage1_48[6], stage1_48[7], 1'b0, 1'b0},
      {stage2_50[1],stage2_49[2],stage2_48[2]}
   );
   gpc1163_5 gpc227 (
      {stage1_49[1], stage1_49[2], stage1_49[3]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage1_51[0]},
      {stage1_52[0]},
      {stage2_53[0],stage2_52[0],stage2_51[0],stage2_50[2],stage2_49[3]}
   );
   gpc615_5 gpc228 (
      {stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage1_52[1]},
      {stage1_53[0], stage1_53[1], stage1_53[2], stage1_53[3], stage1_53[4], stage1_53[5]},
      {stage2_55[0],stage2_54[0],stage2_53[1],stage2_52[1],stage2_51[1]}
   );
   gpc615_5 gpc229 (
      {stage1_51[6], stage1_51[7], stage1_51[8], 1'b0, 1'b0},
      {stage1_52[2]},
      {stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9], stage1_53[10], stage1_53[11]},
      {stage2_55[1],stage2_54[1],stage2_53[2],stage2_52[2],stage2_51[2]}
   );
   gpc606_5 gpc230 (
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[0],stage2_56[0],stage2_55[2],stage2_54[2]}
   );
   gpc117_4 gpc231 (
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5], 1'b0},
      {stage1_56[6]},
      {stage1_57[0]},
      {stage2_58[1],stage2_57[1],stage2_56[1],stage2_55[3]}
   );
   gpc215_4 gpc232 (
      {stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage1_58[0]},
      {stage1_59[0], stage1_59[1]},
      {stage2_60[0],stage2_59[0],stage2_58[2],stage2_57[2]}
   );
   gpc606_5 gpc233 (
      {stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5], stage1_58[6]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[0],stage2_60[1],stage2_59[1],stage2_58[3]}
   );
   gpc606_5 gpc234 (
      {stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5], stage1_59[6], stage1_59[7]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[1],stage2_61[1],stage2_60[2],stage2_59[2]}
   );
   gpc207_4 gpc235 (
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5], stage1_62[6]},
      {stage1_64[0], stage1_64[1]},
      {stage2_65[0],stage2_64[0],stage2_63[1],stage2_62[2]}
   );
   gpc207_4 gpc236 (
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5], stage1_63[6]},
      {stage1_65[0], 1'b0},
      {stage2_66[0],stage2_65[1],stage2_64[1],stage2_63[2]}
   );
   gpc1_1 gpc237 (
      {stage1_0[6]},
      {stage2_0[1]}
   );
   gpc1_1 gpc238 (
      {stage1_0[7]},
      {stage2_0[2]}
   );
   gpc1_1 gpc239 (
      {stage1_0[8]},
      {stage2_0[3]}
   );
   gpc1_1 gpc240 (
      {stage1_0[9]},
      {stage2_0[4]}
   );
   gpc1_1 gpc241 (
      {stage1_0[10]},
      {stage2_0[5]}
   );
   gpc1_1 gpc242 (
      {stage1_1[6]},
      {stage2_1[2]}
   );
   gpc1_1 gpc243 (
      {stage1_2[6]},
      {stage2_2[2]}
   );
   gpc1_1 gpc244 (
      {stage1_2[7]},
      {stage2_2[3]}
   );
   gpc1_1 gpc245 (
      {stage1_2[8]},
      {stage2_2[4]}
   );
   gpc1_1 gpc246 (
      {stage1_3[6]},
      {stage2_3[2]}
   );
   gpc1_1 gpc247 (
      {stage1_5[6]},
      {stage2_5[3]}
   );
   gpc1_1 gpc248 (
      {stage1_5[7]},
      {stage2_5[4]}
   );
   gpc1_1 gpc249 (
      {stage1_6[6]},
      {stage2_6[2]}
   );
   gpc1_1 gpc250 (
      {stage1_8[7]},
      {stage2_8[3]}
   );
   gpc1_1 gpc251 (
      {stage1_8[8]},
      {stage2_8[4]}
   );
   gpc1_1 gpc252 (
      {stage1_8[9]},
      {stage2_8[5]}
   );
   gpc1_1 gpc253 (
      {stage1_10[5]},
      {stage2_10[3]}
   );
   gpc1_1 gpc254 (
      {stage1_10[6]},
      {stage2_10[4]}
   );
   gpc1_1 gpc255 (
      {stage1_10[7]},
      {stage2_10[5]}
   );
   gpc1_1 gpc256 (
      {stage1_10[8]},
      {stage2_10[6]}
   );
   gpc1_1 gpc257 (
      {stage1_10[9]},
      {stage2_10[7]}
   );
   gpc1_1 gpc258 (
      {stage1_13[6]},
      {stage2_13[3]}
   );
   gpc1_1 gpc259 (
      {stage1_13[7]},
      {stage2_13[4]}
   );
   gpc1_1 gpc260 (
      {stage1_13[8]},
      {stage2_13[5]}
   );
   gpc1_1 gpc261 (
      {stage1_13[9]},
      {stage2_13[6]}
   );
   gpc1_1 gpc262 (
      {stage1_14[6]},
      {stage2_14[3]}
   );
   gpc1_1 gpc263 (
      {stage1_15[6]},
      {stage2_15[2]}
   );
   gpc1_1 gpc264 (
      {stage1_17[12]},
      {stage2_17[4]}
   );
   gpc1_1 gpc265 (
      {stage1_17[13]},
      {stage2_17[5]}
   );
   gpc1_1 gpc266 (
      {stage1_17[14]},
      {stage2_17[6]}
   );
   gpc1_1 gpc267 (
      {stage1_18[5]},
      {stage2_18[4]}
   );
   gpc1_1 gpc268 (
      {stage1_20[6]},
      {stage2_20[3]}
   );
   gpc1_1 gpc269 (
      {stage1_20[7]},
      {stage2_20[4]}
   );
   gpc1_1 gpc270 (
      {stage1_21[5]},
      {stage2_21[4]}
   );
   gpc1_1 gpc271 (
      {stage1_24[4]},
      {stage2_24[2]}
   );
   gpc1_1 gpc272 (
      {stage1_24[5]},
      {stage2_24[3]}
   );
   gpc1_1 gpc273 (
      {stage1_24[6]},
      {stage2_24[4]}
   );
   gpc1_1 gpc274 (
      {stage1_24[7]},
      {stage2_24[5]}
   );
   gpc1_1 gpc275 (
      {stage1_26[5]},
      {stage2_26[3]}
   );
   gpc1_1 gpc276 (
      {stage1_26[6]},
      {stage2_26[4]}
   );
   gpc1_1 gpc277 (
      {stage1_26[7]},
      {stage2_26[5]}
   );
   gpc1_1 gpc278 (
      {stage1_26[8]},
      {stage2_26[6]}
   );
   gpc1_1 gpc279 (
      {stage1_32[6]},
      {stage2_32[3]}
   );
   gpc1_1 gpc280 (
      {stage1_32[7]},
      {stage2_32[4]}
   );
   gpc1_1 gpc281 (
      {stage1_32[8]},
      {stage2_32[5]}
   );
   gpc1_1 gpc282 (
      {stage1_35[7]},
      {stage2_35[3]}
   );
   gpc1_1 gpc283 (
      {stage1_37[6]},
      {stage2_37[3]}
   );
   gpc1_1 gpc284 (
      {stage1_37[7]},
      {stage2_37[4]}
   );
   gpc1_1 gpc285 (
      {stage1_37[8]},
      {stage2_37[5]}
   );
   gpc1_1 gpc286 (
      {stage1_38[3]},
      {stage2_38[3]}
   );
   gpc1_1 gpc287 (
      {stage1_38[4]},
      {stage2_38[4]}
   );
   gpc1_1 gpc288 (
      {stage1_38[5]},
      {stage2_38[5]}
   );
   gpc1_1 gpc289 (
      {stage1_41[6]},
      {stage2_41[3]}
   );
   gpc1_1 gpc290 (
      {stage1_41[7]},
      {stage2_41[4]}
   );
   gpc1_1 gpc291 (
      {stage1_41[8]},
      {stage2_41[5]}
   );
   gpc1_1 gpc292 (
      {stage1_41[9]},
      {stage2_41[6]}
   );
   gpc1_1 gpc293 (
      {stage1_44[5]},
      {stage2_44[3]}
   );
   gpc1_1 gpc294 (
      {stage1_44[6]},
      {stage2_44[4]}
   );
   gpc1_1 gpc295 (
      {stage1_44[7]},
      {stage2_44[5]}
   );
   gpc1_1 gpc296 (
      {stage1_46[5]},
      {stage2_46[3]}
   );
   gpc1_1 gpc297 (
      {stage1_49[4]},
      {stage2_49[4]}
   );
   gpc1_1 gpc298 (
      {stage1_49[5]},
      {stage2_49[5]}
   );
   gpc1_1 gpc299 (
      {stage1_49[6]},
      {stage2_49[6]}
   );
   gpc1_1 gpc300 (
      {stage1_50[6]},
      {stage2_50[3]}
   );
   gpc1_1 gpc301 (
      {stage1_52[3]},
      {stage2_52[3]}
   );
   gpc1_1 gpc302 (
      {stage1_52[4]},
      {stage2_52[4]}
   );
   gpc1_1 gpc303 (
      {stage1_52[5]},
      {stage2_52[5]}
   );
   gpc1_1 gpc304 (
      {stage1_53[12]},
      {stage2_53[3]}
   );
   gpc1_1 gpc305 (
      {stage1_53[13]},
      {stage2_53[4]}
   );
   gpc1_1 gpc306 (
      {stage1_57[6]},
      {stage2_57[3]}
   );
   gpc1_1 gpc307 (
      {stage1_57[7]},
      {stage2_57[4]}
   );
   gpc1_1 gpc308 (
      {stage1_57[8]},
      {stage2_57[5]}
   );
   gpc1_1 gpc309 (
      {stage1_57[9]},
      {stage2_57[6]}
   );
   gpc1_1 gpc310 (
      {stage1_58[7]},
      {stage2_58[4]}
   );
   gpc1_1 gpc311 (
      {stage1_60[6]},
      {stage2_60[3]}
   );
   gpc1_1 gpc312 (
      {stage1_63[7]},
      {stage2_63[3]}
   );
   gpc1_1 gpc313 (
      {stage1_63[8]},
      {stage2_63[4]}
   );
   gpc1_1 gpc314 (
      {stage1_63[9]},
      {stage2_63[5]}
   );
   gpc1_1 gpc315 (
      {stage1_63[10]},
      {stage2_63[6]}
   );
   gpc1_1 gpc316 (
      {stage1_63[11]},
      {stage2_63[7]}
   );
   gpc1_1 gpc317 (
      {stage1_63[12]},
      {stage2_63[8]}
   );
   gpc1_1 gpc318 (
      {stage1_63[13]},
      {stage2_63[9]}
   );
   gpc1_1 gpc319 (
      {stage1_64[2]},
      {stage2_64[2]}
   );
   gpc1_1 gpc320 (
      {stage1_64[3]},
      {stage2_64[3]}
   );
   gpc2135_5 gpc321 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc322 (
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], 1'b0},
      {stage2_3[2]},
      {stage2_4[0], stage2_4[1], stage2_4[2], 1'b0, 1'b0, 1'b0},
      {stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc135_4 gpc323 (
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4]},
      {stage2_6[0], stage2_6[1], stage2_6[2]},
      {stage2_7[0]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[1]}
   );
   gpc606_5 gpc324 (
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[1]}
   );
   gpc2223_5 gpc325 (
      {stage2_9[0], stage2_9[1], stage2_9[2]},
      {stage2_10[6], stage2_10[7]},
      {stage2_11[0], stage2_11[1]},
      {stage2_12[0], stage2_12[1]},
      {stage3_13[0],stage3_12[1],stage3_11[1],stage3_10[1],stage3_9[1]}
   );
   gpc7_3 gpc326 (
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5], stage2_13[6]},
      {stage3_15[0],stage3_14[0],stage3_13[1]}
   );
   gpc135_4 gpc327 (
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], 1'b0},
      {stage2_15[0], stage2_15[1], stage2_15[2]},
      {stage2_16[0]},
      {stage3_17[0],stage3_16[0],stage3_15[1],stage3_14[1]}
   );
   gpc207_4 gpc328 (
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6]},
      {stage2_19[0], stage2_19[1]},
      {stage3_20[0],stage3_19[0],stage3_18[0],stage3_17[1]}
   );
   gpc615_5 gpc329 (
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4]},
      {stage2_19[2]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], 1'b0},
      {stage3_22[0],stage3_21[0],stage3_20[1],stage3_19[1],stage3_18[1]}
   );
   gpc2135_5 gpc330 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4]},
      {stage2_22[0], stage2_22[1], stage2_22[2]},
      {stage2_23[0]},
      {stage2_24[0], stage2_24[1]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[1],stage3_21[1]}
   );
   gpc2135_5 gpc331 (
      {stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5], 1'b0},
      {stage2_25[0], stage2_25[1], stage2_25[2]},
      {stage2_26[0]},
      {stage2_27[0], stage2_27[1]},
      {stage3_28[0],stage3_27[0],stage3_26[0],stage3_25[1],stage3_24[1]}
   );
   gpc207_4 gpc332 (
      {stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5], stage2_26[6], 1'b0},
      {stage2_28[0], stage2_28[1]},
      {stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[1]}
   );
   gpc3_2 gpc333 (
      {stage2_29[0], stage2_29[1], stage2_29[2]},
      {stage3_30[0],stage3_29[1]}
   );
   gpc15_3 gpc334 (
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], 1'b0},
      {stage2_31[0]},
      {stage3_32[0],stage3_31[0],stage3_30[1]}
   );
   gpc1163_5 gpc335 (
      {stage2_31[1], stage2_31[2], stage2_31[3]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage2_33[0]},
      {stage2_34[0]},
      {stage3_35[0],stage3_34[0],stage3_33[0],stage3_32[1],stage3_31[1]}
   );
   gpc623_5 gpc336 (
      {stage2_33[1], stage2_33[2], 1'b0},
      {stage2_34[1], stage2_34[2]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], 1'b0, 1'b0},
      {stage3_37[0],stage3_36[0],stage3_35[1],stage3_34[1],stage3_33[1]}
   );
   gpc1163_5 gpc337 (
      {stage2_36[0], stage2_36[1], stage2_36[2]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage2_38[0]},
      {stage2_39[0]},
      {stage3_40[0],stage3_39[0],stage3_38[0],stage3_37[1],stage3_36[1]}
   );
   gpc215_4 gpc338 (
      {stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage2_39[1]},
      {stage2_40[0], stage2_40[1]},
      {stage3_41[0],stage3_40[1],stage3_39[1],stage3_38[1]}
   );
   gpc207_4 gpc339 (
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5], stage2_41[6]},
      {stage2_43[0], stage2_43[1]},
      {stage3_44[0],stage3_43[0],stage3_42[0],stage3_41[1]}
   );
   gpc3_2 gpc340 (
      {stage2_42[0], stage2_42[1], stage2_42[2]},
      {stage3_43[1],stage3_42[1]}
   );
   gpc207_4 gpc341 (
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5], 1'b0},
      {stage2_46[0], stage2_46[1]},
      {stage3_47[0],stage3_46[0],stage3_45[0],stage3_44[1]}
   );
   gpc2223_5 gpc342 (
      {stage2_45[0], stage2_45[1], stage2_45[2]},
      {stage2_46[2], stage2_46[3]},
      {stage2_47[0], stage2_47[1]},
      {stage2_48[0], stage2_48[1]},
      {stage3_49[0],stage3_48[0],stage3_47[1],stage3_46[1],stage3_45[1]}
   );
   gpc117_4 gpc343 (
      {stage2_49[0], stage2_49[1], stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5], stage2_49[6]},
      {stage2_50[0]},
      {stage2_51[0]},
      {stage3_52[0],stage3_51[0],stage3_50[0],stage3_49[1]}
   );
   gpc623_5 gpc344 (
      {stage2_50[1], stage2_50[2], stage2_50[3]},
      {stage2_51[1], stage2_51[2]},
      {stage2_52[0], stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage3_54[0],stage3_53[0],stage3_52[1],stage3_51[1],stage3_50[1]}
   );
   gpc135_4 gpc345 (
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4]},
      {stage2_54[0], stage2_54[1], stage2_54[2]},
      {stage2_55[0]},
      {stage3_56[0],stage3_55[0],stage3_54[1],stage3_53[1]}
   );
   gpc23_3 gpc346 (
      {stage2_55[1], stage2_55[2], stage2_55[3]},
      {stage2_56[0], stage2_56[1]},
      {stage3_57[0],stage3_56[1],stage3_55[1]}
   );
   gpc207_4 gpc347 (
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5], stage2_57[6]},
      {stage2_59[0], stage2_59[1]},
      {stage3_60[0],stage3_59[0],stage3_58[0],stage3_57[1]}
   );
   gpc1415_5 gpc348 (
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4]},
      {stage2_59[2]},
      {stage2_60[0], stage2_60[1], stage2_60[2], stage2_60[3]},
      {stage2_61[0]},
      {stage3_62[0],stage3_61[0],stage3_60[1],stage3_59[1],stage3_58[1]}
   );
   gpc1163_5 gpc349 (
      {stage2_62[0], stage2_62[1], stage2_62[2]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage2_64[0]},
      {stage2_65[0]},
      {stage3_66[0],stage3_65[0],stage3_64[0],stage3_63[0],stage3_62[1]}
   );
   gpc2135_5 gpc350 (
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], 1'b0},
      {stage2_64[1], stage2_64[2], stage2_64[3]},
      {stage2_65[1]},
      {stage2_66[0], 1'b0},
      {stage3_67[0],stage3_66[1],stage3_65[1],stage3_64[1],stage3_63[1]}
   );
   gpc1_1 gpc351 (
      {stage2_0[5]},
      {stage3_0[1]}
   );
   gpc1_1 gpc352 (
      {stage2_7[1]},
      {stage3_7[1]}
   );
   gpc1_1 gpc353 (
      {stage2_16[1]},
      {stage3_16[1]}
   );
   gpc1_1 gpc354 (
      {stage2_23[1]},
      {stage3_23[1]}
   );
   gpc1_1 gpc355 (
      {stage2_48[2]},
      {stage3_48[1]}
   );
   gpc1_1 gpc356 (
      {stage2_61[1]},
      {stage3_61[1]}
   );
endmodule

module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [15:0] src54;
    reg [15:0] src55;
    reg [15:0] src56;
    reg [15:0] src57;
    reg [15:0] src58;
    reg [15:0] src59;
    reg [15:0] src60;
    reg [15:0] src61;
    reg [15:0] src62;
    reg [15:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [67:0] srcsum;
    wire [67:0] dstsum;
    wire test;
    compressor_CLA16_64 compressor_CLA16_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he234b25f7fb5f4b0c6ccab00e1d9112646b8c0bea1c6ccf7bcd2af4b6cbbc20f57e99d2a86a30b6e92c3a3d152ca55bc9d12f2c8c7f6cfa76cec990b21fd7a9302e0b326edb1d150c2c1dad4d7edfd1738db1280974158f0cce7bd01ac7cfb37f59fa19d39b9c1ed1c31c2984260b832ec9bed24a9f6d98e1b3b7fe1587ef46c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1e02136fb83cdf282f9291bc4b3001552d7b45cf4b92cbe80f4db32cd831e5de37d2e30bd1f7b65bef93b0c6cbe8b6c3d376688b740e7f75e63dcc988a7a2bd44bc7c920b0a4d7a723961c1b7f899a5875d50b3b8d80f4b467097b9e6d0529e33418fcc01985593ab536b0dad6c00578e9ca1bcf061c856775ec62f84c501a8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39f5d4d81ee6a584988f61e72048b71872f72249b8a2484b7088bc271f49aa30b84eba109966738a83debb6f319809a96ef0db8a6038b454cd1d9a0c51801676a1900ea8d308429b1076e3eeda6e6c57e5f3994a4bf6b5a8d3c78a099f4ab99a860460c920428ed286f3cee83f76640bf7e28982b4b1b7c52ac399079b440f8f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb1074dd6ab75eecb3f6ec7520d5ffd2a8d9fffef249e204b9527ae3c74d0f6dc42fef4bb42a8bb47aff2022f55e9ade6a37ebb33fa0ca5d308e89f99f90241f87140520e90b3606c65d7e19f0a06d27d6491a76ce16a0df0847a3a74b4b76cfe71def86f609ab8895b3d3c7213e9adb2012963d571ab8db75b9a84e5064ba03;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a11e97c7f14ead4a6e6d0c3cfe994b92c73d921413896792811afbf11ee03c3807f5c7dbb09fc7f82121fec4f6d20da75c8c0fe76a912fe6b46a1182134cb064b0ac0e93f0e3a6c766bfd6ca6cf179ea64f7d661cce65f907fe341306320be55eefcfb68e0c632fd9cfe09ab197b13abd96acc0bb5d70df4f60a02f831e892c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4840e1624d23a0c4414c0f8b4f18425effc797efbf927e5a8951b93a4988a17199eb1ab534c30716c643acdae3d11075d2b20e48a7e69f8fb9b551e2ea29481a2f1900bbfe00c267d42b24a646159314d73e9d8a66efc90fffdd455cb90814744d0f74993f817f2ebc43946bc3e173d54bef67dbc0f6fceb0cce53f372bb454;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcf6512af0ed12f5ac7fbcd2ed5b1314219500da0c07e5c19ffec24cccf601e28a4b3359e5dd5b643ce0ef28afe73571697c856bd76d79cff37f5d3df55e65dbc3f7cb5a6cd32aa1f63c44406fee2199ef32f11d660818e098095faf42d89ced897bf627a337a7939869a58a4575e4521bbc7a29daf385a6ce9951bbd2c99077;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18b842209b3a3cfae081a2a4fca0537f350412c8a903fb56340d90b92af4c4c899eac0faed78e99f4cdff4f217ee9d7703faa940e59d268b5189fb70fdb7a7fbbe28e59a5ee3ff98420cede88566afce89de267f3f2028b06eae9632618b451e6311f5f492f5fae5d539acc335ca56f46d0b4c0e71e7734481fa2f44266a341f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf67e98acc126c495e26ba5ad899110f0fcc5559655fc23143ddd070c5cba691b600f0e0ed73180bd3e68d66b475b7a14d32c64dfb84354b9c3ec2ce1e408fb46d87de0feb0b51932cd03a9e20b18d27cf1beee7cc0ad3d55b3a07e9133301af31250d879a631cc1da3fbc57e80aa99813f0fbc974f6aebfe26983d25e88e8ad7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf862ebe9fd7908fa94bed331bccb06fc847480af64be6d44af053be70fc237ce32e9c2baf1c8a34c32ad6de5164d76c4bd6be44f1ef7d1c7095602b895d1e9fa409e9511692add0f5faeca755f5db58a9ad4114b613b1b9cbc5bbc2a9562f7e198abedcd51410ae7d1b28f671926b0849d1cc2748e6a80261fe5ab093b7023f3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he34516da39a35ba29afcb25edab137c1b7374c5b7a29569282b91446f8b3b8fabd07e001b3cf93453d9763d09bb0da8a853f1ad3f2564cb99d12bef50a5d9c3ef57fd038d0f5a2f3d54eca3bcc6dc053f8fc42c39825587abf3c005eae4f7b533c6f6f15b7bf22dbb2f773039b0051bccafdbb75a2f51fab4945e55d1c2aced3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd225c08c8c16c581c8f7b8998982279780fc94d0a2e8b431c4f372eb74b32ee35d63ed0164f1c27697ed530b286d6d847c96f6287056c789204e2d9224d114766a8d7b8f2b0966c7d1578047bba55176352a4968b10788f95f39a1f1ba7df9f8bdc1c6d077882a8a5194f5cd18b644450d2a7ce1a13d12cbeea38ca8f609579;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b3e697cb269c24c5c19d6d300d2f7b9459850a48f47457b9f0b35350e6676bf05f54ad1d0d08ed7cef268abe9d9aead035b84c22a0710990313f4c704bd7b9ca6823f6ef70b3d4547d5e68533a88d305463c6e9ef415b8817c27448b6d65631d550b8f6d6e1ac97a4ca53fb2842ef9dc0baa96ce0c9e3ab1f7175a2201c624;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b13c0d2dbb967f9484ae7a4323de9c08dd0a0ecbcdee3e2c0c285aab2906bc8227d15d35deede9756b3cada1feee283a555fb75cb992ecd37878c0c7a19708ea752f0459746e4003ce59a6ce6cb938ba1f56a6e1745b787a7340223dc13a7dbe01fce2499e8ef045179812287835da14d03a2fdcf17294a5ec4867647cd9be3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5485147a490b7b840843630753646fa3244e792ab3b135c279fe28d6ecfc83b9ba7a25fc84ee4c6c404ded936dde30d851706ccd76e2046f14269ebf5a591ae7b309831ca7535fca04e69b041ff86106fc28092e5f211865049d950174d2233899dc6aa984bd5d2f939052a4673bd866c8ba702a95cb4a0c12ca3483cce11784;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2206bd4706a704ca1e7736b3018889aedef8fe3fc5b6372186620fdb9b97c1a3081cfcf179ea083edacf557c93eefbfb5e3444c707dc7ac5135c498f5876bc3f67cd5c63c3b215b4ce3c712561c19384d7066ae5ada2297fadc7cc82ccb933005882b0537b3939e7eff221e5d6b0c9bbd32372f3cab43eb9450314dbd1125ae9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d29e32c2e168e653834eb218abc15c73ead856361b8f23d0ba56e26b9f68ceaced7699320682a2587eba7c09fc80a235dfe5b839e2b187384b2868ab30ffb05b9e52bb350b9599184ead446e8c45ce10343c6f7d0352b82ea04ed7c9b4a1dbb020aece85706ef2ec8c6b46a30576ff6190d085a4015987cd4d7cf8b1333efd8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60b65c7d81dd64ebc0e048fe2095df3103c72debe0acf08fec26ff139118d584e87b21b85b8011ef423c0541d075f5a8ff4a014aec987fca93d29766ddebf3e09c4c5c0f3891d2602b6a29e62b593f835b3ddcf8d6f027676e0f033f0a0ebb6221f26db3ba2a205b221266ed56a30e20b959198357eab17ebdeb8952b86678e3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cfeb78933f99ed389fa44a1bfd0d2a9f2e0f539a1b90c228f5617cde39e28bda4bdf3b02223323caed37aeeb0ee4d44df6a057fa9e1cf838eaed1fc49d57af78f6f171dad8b2c54691645a9f00b7094c59edc91b65865b3bf53ef79aab6ffd0a3af754b06afe7766b8cae992e662ff886e1d177bdfbde90ece57a88738f9387;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37a03500c86cfecdd91388f1886a54122300717ef41c361da83f03e366b1ebda58ba4428230d5fd95561ddc987784af2e8407901c4952e6ee3d213ad7d859a5b25719b36a0946d3a1a864ba107657f3342b6a722c60261fe9d7e113e7052df4dfb2980412c8c3509eca68ac7dd4f57d887335673d9b68e69bfad887ea587147e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1d5f2633271f31273c5284a124aeb38c262059f0e9605322c082941c3bcb940074e18f9b9b06c454ce4d8a6cfc5fc02281f1a8b29a52e9fef1d35ea49736d80581bab9d9e639bc0672aac6838b687838218c7960037bd552e1e98076419c7de18aeb909b8231e76eb5ab22a0d4fe964a5993ca7b1a8bf3e3abf7e0e71281a53;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf125b4c3de095abe01ea7c67bdbe5a11cb2123cd56e9f40fc005a6cc1a6b9395ab76b4acc4afe30066f119087fd89555372bc594bc443778f5343e34b3bef8d63c36a0a64bd8a6419ce1937352522ca5877db20a11072ffb45207778d6344d45644452eed29e21f692baef7893b819c93e175840f67ab5f3e9c117725123d204;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7d897c9a12f0eae132e239ed1e2cd2b726ac85d2413083b99de6e23b8c7e280d22971f076ff35549d8be93b2d04bc950792654336352d21e26e3b54c8713b5e063db2e3318fce595047622d4b6beee3c013b64831ffbd5a82778eb2b87de88f8c755672cfbbb160481ad7c7971ead6ba792f512734e0db1a63dc4a38477c80f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62376d68dbc3a96062aa5c56ecf3b90347586a19327b4a7b6e5d17366025efeea88b8da96c4395ef417beda7016169c2daf45f54f9f03b6453bdb6464134a088f1230019c2e3f0887688a82f252cb718a4f1ac20360a635c22ee9f6c70e659718aa2d8183860cc63f35121801c3f9de0e8dcf49c65e470bd22e81507e675b807;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf12e2f0391c00b290ebb7433d5af07642c3a914563c9b8b55ab736ab26d01eaa4d8596f9c1cca508bc728abe9de20f72aea546501125c3afe42d175a02a3cbea55be3400fb25e1001f8eb08956df92e8b37a9b4ea91f7a7b5301d135a324864c9b81baab8923a6d29b50ab8b2bf0d98053346b6ee8207a5ab00f1dfc9dd6ca15;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he972bcc05af8f0568e26a0f8336818d7c2bb573ed302510e82930e58a1f87c14025ff86cd3f08331a1d143dbc1d4b89bc48e7d278f5a34c82807b7212cec3016734c58058f13cf89abdb93e73dd6e53de2927a74564ac60c7a06a3312c5b1aa70f75d9591a52710e7c3e3f9e55cc8d07c0a846f459caf05ea4c60206aac35a5f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7c3abd39ef0bfeddb7700b6d92b2f747bb85753a15a9e1f26b66a90aa740234676b91f5c34bce7a37a7d95f2fb924278518d6135f2c2becfd51040c5ff92063ce78b2ccc9e421919a56195158413a9e898b5b71f1ecb6943d12487e567b1b974fec1f9c96017857cd3bc8e6f6fd973a541bcb77298e0ed2e9879ecfbdd4eeb1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc812739bdc6fdd7e75d10b8319643582d69774f03b5eff50dab3961d594026113bb2a3031af18972af56907ccf5e16977cdae8e39d03ba2c2fdc02cb6f146c2b3ab6ca1fd4321042f3cd8335f038af2c0ef78e3d278098dd89eb4aefbdcb313121e5359c51675345094dea2173255d0a1355c662d078b81e80050c3250132e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1175a0cd8f2b3a8b3beb218045460a63763d89b504309a88cd3e1c03dba108de861b19521517ec32febed78de8845584a77bfe6518377572a957182e7caf4816b2e067fb60b1bb15bb6c9d39dc35b7f7ee4d989439ede3385f8551f9a49abdfa91ded7e5d69a03c57c1f27389fbc41a86c2e1310281238f70022cc636f11f725;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9099723a1128dbdf3821721d99605341640b2569f97f63fb808134d092211d88eceb0775aea848a335a8db66c178fbc0ec5ab271cd4d3fa04a489128e3f52fceb1c7bc1c939dadb36025a53198f73f7e2b38f5849da41edb5385b4ef75d1e68c7e44c1f921f5ba42b5daa6ad2731b3ad298e4cc99312ee606cd01fd245db3624;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a9838c3caf5ab352a5178e5d414337fcc664f0b5f3dbaaadee37b37405f9cb707206383eb3c8717bf5c16b349fa18bb29bd6d749cbd9c8742e8229cc03ecd44696cdf47b670dc380c4b0653fdcc106d29af5ab6f2aa942b522fc5f25cadf57a5463711721ad3faead0cde4ef93f0b7b1350c4a4490dc406c5ae3af0ddfedd1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he38e78dadb0de56273ab7df6a82a47f1d08a5d95c92fff22484f2a5e8d696897a5617d75cceb467cb10c9abc451869903c84527fbcba54cd5d8811a7f65e51c26344553a8f44106fedfafdd23765deef51c5afae773aa6a1037856a2871cb099c8f0cd1f729c30022a85a04aca04821fd9805f8234229dda596d7a8d2ff8685;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75fb95078e65d6cbab0e468be7505545ed014025ca75e67443b5cfa287a8abd3e8221bbf4977fd2d073bbe473a8180ad1d2d817ac774fed4c05fb628d0b630fead9c4ef6b0aa030e442379b284bb5408e568cfee359ee22a42bc78597d37393e36bd9060eb8cf847cc12acfd476ca8bd7af19d4df6b97a346378493d071d4871;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h867e08b4ceb4360bc81e6ab5a4c31dbc4fa81517093bcf9ad50a78be95394cfb7ccdbb6d2ffb9004c764869dac59f0aaaae5379760637c34d61931de0c0e8c21b5627c26c5d4d7d27c0226e6d87d385e678736df577930c7c686f5eeb4532b1e441784e8376300b991a6f0058d09a1545ed1ac754a597550ed7722512139b444;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70b504405afa4a98de7ae7bb8ad55f9337ddf4f1d01b0d8b014f14f652b9fe70a4baac064b52493aed131c5c2a2ac4b1ef66e3cb304017e3556443126b717fa2afd516965b1a3592e806fbae1cc69337a03f7e156b3b9f2f79cdd8317fd74a64b39147a6b1a0d801b74bcf98eac6f43209f995c0b07b72814a7e639b3827e6d3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h483b6edfea14d4c91bda9db100f044d59b23fc53d5fe2b30ad746e0801ab5b70e8357d9f91cda1e28fe99d91f723d52301cdaef55f5615da2ed9a1a6b4e1e202dd8388a320c9ff16a2a1a57531c5838c2216537edea257181e097b8774b608402b3d791e97a8e014d9a694a9ac7918674cecd0af4f9ed2cdfece5cad99b78115;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d5f2544f477d77b2be9927beab35a1bb258caaa768d63e8abf6efe2a9c4987c261b82dc3605777623a84d09341503096291e7abd69c36ea3d66ebe0ae147dc5f6713d5c74dbe40afe46b0784ab2ec4fc29669cb839631e6aa215ac4cdb454c1b76593790d115ca75ef6147beafff4902e0f15d21c1f68848b02770be43cf7f4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8047a8dce1517676449d5739d653672803bc540203f03ab1f5d99f208babd361b690a9297e9dec620239bcd1bc4b3ad98a26d2cfd7a7a3f75d7b2a45a9f23ec5d6794f7a5e2dad368144df6258be6c32e11d69dd3ad8bd705fee22e9860f012419604e59c4147fffb4ea71da7a62a6e1b3d304162fbd6eb2ec6102e7f34f8d71;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bd43973e3d81ce1a20e28e94eda4d55aefb135650fa246883b41d7d9e1e21e3e9a8a1afa1f79f349b7529178a5d30ab53db020f889415d202bd2bcb5401e45d61d4a50eca93c9785d8bb0a748b2f00017903185791e5a6fe2edaae9cfd37977097b839951397f57551686da21efe29c884faddec8bc34a2a71d5322f9e67278;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18551acff6a4845fb0a4e557101bd3278eae2dee31e050041ba0bc81c3bcdb4c4a11edd49f89d12ee09a26fbff1b1e483070d71b3e55f8ac755ebffcd0d6d713da56a419d55c9153b5af67a0292dad22332a96cf24e3a2b18419df9f13e30cfb5ee6aebad71c95109189e7a183ea8223a1f590543fce5594e83d95e6d0597d3c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc92f8fc9446adf8cf9fc2ac4f9c31e50740dc433d4fcc98452609e2861f21124592b8fd397841cfab81322b4715de7977ec1fcca5fa596441b94b74aac4ccd0002759e43cceb056bcd7d3331fc02257c0866df03f1ca05f6e1f745bc4487b841e17a1995ccae1e003dd20f8518b2d998ad3b07c6e341bf088290d33b7cfc9b2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b7ac4ad82776769387a41aff7ffe9f3fb436583910e5f709c5d3fe65a858e78c5298d8f493325f31cd98ee0f6610a5c0324b264bc112f72eea0ae06642d2d96febed6017408b7ebb2b47335d428be4e16302dc63d5d0ec491bc7ff2beb51ef0a81d7a9d2dda6dd883d8a1050fc18731c718bbb8e905c9721ff3c639dbd1ae6a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d8a0869b0fbb7fc95c1a191e24b11b52868e6cfb7dcd5ee578c7e0d04bf162aa3fcd570db4d88f0fb4193826652307a05da13a1286a213e7404ec154ae96233aa29b21beb38e8bd0cd0133ddaa08bbcb8d66f1b83a352429870eb4e4a945a1eeaacd293288e4e454862f506ef557be08773889f3ca55856921ae97c9be65bb8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d0b372aa50ca73cdbb05d119f5e4aa3ed1c92eb9802b86559389e62b92a0e78f9338d0a9fd173476639f5bcaea700e57deceabfbc5c58e5b997e73438e0646b4735a2430d1ba54691a49d27bea4f6f94379b16a1c54e7bba3754b014a382b2d35e938f2adfe1a46cd18eb3727233a0a48e39b53e07b0ff47743eaff2253cdcc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3367dda2b58a9682980e1069ebbf24d0d1aeb0d2cae8093c851639246a4bd7edf490dc7330f424587c915065ce830f712c7bb0872a0516d104982b51c4c9c772c3c6114c1a80567dcbf3b8ee14c2484ce3bb3b6bfc04e7bfad1f91a66a25a59000ecf99ee2765e14b810de9ae81dd62ea8b5619902c43c550409952436a3d1af;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3142e95dd916bad7116760ba8cb510d6180155bafabf95e8ec8cb8924a537b0397cdd5f7fb02ca16ab43356e9056c48a0055f8b4aad968fb617debb813ff607488070eeb47d1b42d12183a7d683715b049be4ba162da03c1261d49abce340a31343f853ba1d194efd3bdc65448d1acf6452a63c978b75afb4552e0c4c1caaf2d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd49ff6129004f3d0962defc7f9565d6d69bd8783fc8cac8f5854e51b61af7e3b8a95de0e05e73a573af5f8dd5e3a6cef6355ccdad6a2955d7f0fb2a9736f233586138279fbe24e508199982babfc48caf9075ab9de08a2fe025823e1ade076854611cfdedddc086682231486dbd72b49e5f6f3dc153f7b14056b0e8f8ea625e5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he996f5e4bc094f04bf09b2b3322a187aa10adaffe509dd3c33b8623f94f3a433c710a069335d411dc72c5cdd7a03cf5df02d1e079e747cb5c565aa9f1cc6e9ae9f3234a81fa054c4f9a807f75ac96d73e0ef79dc13305e192c509ce074faa03e6eb38d445f9a57a1176f95290f933bda267ad262e76fc375379e5534d117fdd8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6856b8398e69f9bf0bc77aa6a6dd27f940e056031a27104d92c6a637e129541f5bf8f5346ec832888b0d250fc29e0c4b8dc3f9ab20c6c3705bfc9f1240e46d61a1fe66696118d74f5c5110fb26ed681289111cb3660c630d176537f6625c00d5bc82d83dcaa40cee254d729c26b46ebe5b5ade3727b4e77e81d2b0010e6eb0a8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b8038a3d05e610e24d46563c3b30e26079a866ad31900e7b9a4ed414756c7b7605e151fff4d0f9c0f59847086faccec04546015fcf1934c8a8387770e2b14a63584790ae2462815ffb3cb8e76759dfd6a347d9172a3bdabcaf09c82e8c74caa293268b349968ef135a61d58448648c7ace71bbb5df358e7efe45d65a4f23037;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7de2cd970b88625c11412cca12899c7701efb6d0837875e0dd895d8fd1a18acabfd8edf8e40d1cf6adfde6496fdca00d5b176e19bfa8870ff086cdfa9b1f79f35c8c22d122f52e03863b31a376154ace3ca045bbef0967731f06281cba3964ec96919fc67c7022b46242c7f9826c3ce73ff20c7270038da34b64dae9b12a7d3e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha22c2e2f6fd0705d922955d97053fe06d65595b0b1046d3ca0b3592bb6186fefacceefecf3eeebbbfe5a3433e3e851ad29b9e522070f5326d75997a744e8e4e9b5e1d67eab7ae62a899d357de5c33ab57480660290b0f14b961a7cf750f811423cc12295a9cbe5235ad5af04924ee81bc5ad4e8b61511db875fb3cadb5758506;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he88a35a9e61b3bf137da287bd6c2e435ce9198640bc884e3a2770de64e530c5b761e71b500c77299db2065923383e5bf3d282945874a6b60be3061ac401ba634e160ce5807702359f3e9895316a6338172c9725b335b306488c1da5c79f3f18f7f738eca409c596505cdf1b22b80c720f9241f5ab2055d2f3efac5b600007267;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97339608785c8b4b57643fa93ac63f89d1fd93d540b818b82f3e2c2c64e8a9f500ccd5b2a927f272d72c135188f0a3151375f9d42d4e0c3ee73b76d1049902e2e9808b5ed616c1f233b9c0bf9dcc150a200120b37192ba6a93431cb948f58bb5b88dd8ee1da71f44bc4032e4a09a9f90c66626aeb1ee2a60171139ebf0c3ad16;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdc3b0e53e97063e4cbaae8a99135c40a2bc777672210dde6559d5f21d6b8ef259c88b8130b63b22b293c5fc204956e2b6b6615114e5a1a92caf2f5eefaf43532646ed3fac4d3e8f753c2fd6a149092112b592a5a35737219cb3e858fc30d1287b21d83040d39c84f185a1fe341989228b05f5a007a0ba65617ff1960db0f3cc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcfb3f70dbab4eb24957c94f67c9a7f599bd5bd030f4c2454391d287fe2c24beab0c2c9ecb950014f6c6e0a10ef0e6a3a44a4ad397439979d586292a27bfba8c0819b9fe520d10de77f2b791158d89e6dd6b14b7b43050f6a81fe545fb0506182b1b58206ce164ee8b25bc48361d74c4a811e84c31380abef6e1f63c0c2a4233d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4560db31c49c4f67fa6f7debfdccff56f6b3c7c96f8ba011e7b1f03b2985caa04d2262e6736433590e1d09d1dcb4c6a3152aa2ada48bd6f8766d799de5ec42baf166df2a7e5c69a16b8d8c1d766b7de60e3e9c6cd0cf561d11e88147593b81bbaa2c1ed040f23df7c4d8278e51f02429fdde95d42f50611a3e04e9e530b278b8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5baf4e6bcca0ccaf538c5d4f8dd85c02a2814366993b84d1cecca4af05657fa4adf18a880c66270dd4cdb01245336d9710bdd7f19b8927ea70cab0b4322144e5f9b9d8b0cd10847d3057b2d205a8da76371d365d9e82245063e8039806c4380612cfd44c399330b9dac969193c8c5540d4e345b04e276eafe171224f3e37a3a5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e05167dfd4dc24e93a20bbba64c585ce1599c2270345b5a1c8f992c6e38ce6f287fa249ab225c870fbbe6de0da72c395e6dccec5f49893a516e575082ca5c6b6313f1f1ffb351445b23b596cb3388e2165b36841ad73a6bda15e6adbfcc03f99db2c7ea486168e421ac9d806e389f6e2e4de1d4f087dbdb9255481b7eb1cefb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he23bbe1bf26b3e61623007821b651ae58591da9544547a703724b1b35fea3ac36b387f8cf6622f874e2924bf5854c471e4780d7a42114f96ba18f165b974fa080a9cb53e0b711e1fd0952a6adb8165c50fb808f777f9a13a75f6aec49046d37bbffba872d913af31fd63054052bfa506b513d3a4f0ccf189f3bf3f318854f11e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a525189aaddec66058ded26554fbac7d6040573cfc5667a0c43f14307af5ea048e65c4c77fd940a2f70c099079ed7fdba40b412e9f064c2649c7199d55cf02b3d41955d9b514e0b66055244177e283986a18bcc5a222cb2e57284c87f22985c2538b9288f50269ed0c589b1a0519f0e343e470790177ea4f235bc311395ebf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1d3494cfcbe403854e96ca8de5df1bf77614e505f8e03e470fe77ddaecc3f940de6bb26a21984eef1d1a8f63d63116cbcc05e624b911b2417cd98e3b14ca9f9ce359475b94a45770fe26e5872dbdb5114e9d43637c3e13a77c7f4c931fa78def71d7c1366794b453d5e1f39ac747e33e25be3cd48761fd1281a940d6f100fc1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7a978b8993bd62012327b5cb27b15cde39ff22b8fefb5cedd5ff834aabfa91070dbd210c8e3f7ef2f2372a90ca7a3f3b6b7638990ad916b4401e90cea15c731ffef0bab715dc1cfc25f66481ec09844fda677fe78166c779c34de178273e8941e4b933cf4465971a7bbd7ba4fe381762304807cdd18a8f333a86e2804464d92;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99eccf4aa21559f7c7f55560d0af780bbade3654c32042f64c1a8b2edc3b5272d0d3e19e9e91d6eab6b27e5389aa7296e19e20bef240534da5815e9cc76d1617c7e92906da3f42c164f5faf917c771c5de4be9ace16961cb5ecfacb3345c1d382e7cb1d1d9f6453a66aeba8ddc1180f321b24c5565521b73999b9d63606892c8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27451564ce48fdf40cdd913c78f52dcc45fb5be1020e0f57ed4d547307573f26cdb38a01b27b769ee420061340e1363e930701cc7502734e9b041c5a8582fbbbe8f87796be7484f71a9b33641b7c7ad6813de0563137a3c2d401152e2f7f1b4913ff221b60b7944593acdabfd55bf4333125f992302ce74dc699f85dbcedb00c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he925b7434996991319a3eeddf30e77670b0d4fb018e48abef90379da7b6a308f195db295997750f27881df1ee562e95148048681462013bb79e7441ac4c91eb3bb17780aeb81103d2565bffd72335052976833d315dba4431c9c8a51fc9e54773481bfd68a37179fccd8c4c8d0234ed3bbc622186a05181ff63c6c020235d750;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf3af7cdab3f1060db57a7c9b959527178f74e408b76b73bd1b3afbe638a9ab61ca3723ab08d686dbf3bb29a31a7134c86dea0cd5fad36bef42fe122e3c2f79560b956ff92907687223f3eb5d02fe884005cdd7fb0a201bf3cf6788f24b969455f9f5ece6206cbe622eed495116a1fc208e8857b91df7c81156b10989f47f2fd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ca3a6da946cca3aeebeceaf2f007eec7b2036336e8471f2cd2f7d0b77d8b295b39ed18a4ad3db98a9c65b88fa7c5325cc449977ae0c28e560b9f9494afe4abaea3c50a3caffcd373c98e805cb35273b87d7dddac951b6bf6b586a7a102b2f945f930decf240f7e93abe8864ae4ef4687d1654a4fd11528e8a4c6cbbf259a2aa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9932e5fffef895db1bdc3743b7591b114ae8a9d8a079faf4c81388092164e9bc3eb5a0539db736124fdd438804953afe9b37ef05d08257f3e9c42b55139cd081e25cf9f24168b1da2de49da83492f346387f700771cec28b3c36fe7fd44d0f43ad1e1c32926144b669cc043057ab4be085e35a23e2ce1b2589aed83cb9cd3b22;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54923541e4922f906e5b891e920558ffcd724fa64f596c7f3389882a5a0c9b484067a4cfaac4a3c1ecfd82d990698f4261bee458a60dd16ce00b11882fb7c6491a965d5f738a5a35ef85d593dfc6f942e84d9f6c9581bf727419ed796fb4f09bc9ec117482a86bf9f5d8485275daa83a4a8e76c248a1b0efefe2af92c9280666;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20a6465c9d40114b78ace4404e391fe6126355943d65981b81e726a8ab1bb2ed7943f5395f8a24c98bebbe1eef2c52bc8cc983ded4421a9f77635ddf23f0b3a989c4e394fdb1ad06cfbd914ae76fff2854d4ae42edd6a65738c3219a8e1658c583990356185ee6c345fc0e53d87970a32dc8eb441588a31700d9eadfc2891422;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bd7bea1778ad9a91f0c71ae0c4e7081c3eeeeccfeca48f360fa75ccefae324805ff6fe39b5253fb6c27b839e5a1b137212255c278fa9f1d2e3590d0a87849fa585d42f2e100b0dd0f57939ce728e01f064e81d41ea132a7e4f296610e4bd6918489fd643fcb5b521615b4f94a36db053deb44b97f0b9010f493d129bec40c84;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d1e7294d05f815bef6206b103aff7021f434315936d03c52335308fc436d9fa4f96d44a7b48800b935f10f6474d9c7c1a1e1b35a573b8550daa6810181823015379acdf3f9bbbbb69282ec6efa54ac069b6abb4023395dd46f354d29342590653ee17256ba2b0e77a7b9e74e163362d9cef338d308d70d725abacdde9d56531;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69e949fdc3c0583801f147381d47e7026fccaca39bf7fe9fff154a7fe0a60381fd7dac58d8cd068ae3f88fa1e6009e18252cf28fe365d30518fa0a20806a6ace0a942921dac64ca2a280ca12640cbee5e274e83a2e89c1cb205dc0bd7746f534bc1fa2639fe84c529ca28e6abd2ed569330ccdd4a8e4690961573166638955f8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde6a859a21a4497cb3463941154c59a89081e7f7fffed2eea74cb42573fbe3ec18039a254ae125072b689c287d388dccf54247ddfe151c8ed87cb2fa581707cb5911b5f73ada021b66c1067b325aff8dc8bea112c4568f4138431b55be399a2e610cb1f60e64969635241894dfd0f2b8ec50fce6bae454e60cb51ecda99cf3d0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14f5511a04d518406e20e06caedbdacee79d093359c5c3c4a7c2c9804a906ddafc6e230c156c8a7d295fc6b5f218d1315b876574748515aaa96724ea0d2aa385e20ca9a8d3d2a82bf99ccc13185c9d4cbc77408391221cba13541d53b5cb23d24e3f384b6ee1e9627f82ed118acc5ae056837f6de3185d33dad2b217d02ad432;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd56c3e9824628844f2936e6e084a052fe151881636095cf7ac3a742085f5adcd0cce5347e9a829eb7905b75e59be1126523f51750371372227f349e2f4a270b00fe0d32f6e6ce83cc6d04979dd9ff086c22decbd06551e6fae539ffa1144172b426443df01b17db5513ecca11b355acc11b34b152490eb48e0cda0cab926a607;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5701b096ce5430caffbfccc100a3a16b322f9392f17cc471d79d55ad701e1f16429fd641f08200c4cdf652cd6ecf185ab2061adb9478329744cb123ff08bb2c4d553db3d34a84b08a30038fecea851d70116ba04347e317207a094428776603edf1f1ff65fa02f89d1a4051586111d0c6c890124b292d5756707e6b49e489812;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2f66de2b4bb58e33ccde0747d2faf76c6b299b01ab6eccb589d0487ce11b40a695dfd37045b23371b81c1bde64b85805d80e49cfc28a89447edad23ca025e9bb7b70da39e4f1fe66790e3127c723001c0a1f07ee2e292cc64b7d5a9e761c91afa24fe6824132d3646aa189a4cf1e0eed0906fa792fb870dd5e06152bf1f897b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6335b5d73abfb3208190efcd51d1f616e848c18e24cace2bed9e1fecdcb48dbf5bb3e5ad268bf3c9da5633888e033aba22c70956350472bc42947b6b355280626622fa30e1c55b323581ddff134b29b411ae926840fdc209ae0385551d714978590bd670ba0acb1651b1171163c6cb732a51750dafda329e00fa4c82ec4b4935;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb376ddb4ace53c2b45cd569d99f841738f835c51768c95eb13ae67d4338f299cce22e53595d7d89b996af134aad9c67deecbae68a9d9d543e94178974cc0a4bc3310ac19ec12cf5f62f868a994f68f8a6c3d4c50755c437b7b2150aa8ddada31b2f988f99c05825316d1f122b4352b5204bf688bec86f31de9bf0696d0b177c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c8ca4e038904160fb6917bcd5cb12873635d2d25386c5134c4b85a44a47925c9ee5a8693eae04aef4541114d5336c124550eb6d69df72ffa076de92defe05fbbef69ee6a750b22ba534bf1a9ca11c7e97fd82eb870f2590af2d4fefab8e790558be1acdf1d9b3be550ad646374eedde2f395959288b5f3057d259135705ab4b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67fb3d6edc292ebf3a4fddc60854c590a1c0d108cdfd77a2d6a27078ba8ff15e8ce15f909f6b9c0cfb2f71bad9f711cc8b54d7b28bed30b12e5534788cbc4842b85c69546f26a55453a7ffeb52a130b20a519c937e5a12d22e0c6d99c50670d8a486a5649d4d7ee871ad61d5812a234e22e05d4fff2771151f32cad4e924801e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5a4a0ec9874dd15d3a5f742cbd3c268a1e97eb584ae4bf28880fb95120ebf280db804b035db50759c5ad4dbdb9f0b016ecd02b2beec9d53292f82a650950d6b7ae9f97f21e589ce7172bf7af0ddf205eec5c750c7816bf73f0c9d9c2f1e989bd4bcc49d04845b108865cad6379cea7371b507ea3d35676492c3ca931e37560c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef0238261c01f2c498c65f99f92cc786ea8e5b5387b36ad731fbddff7c6b1ba8ba50f2c67f6ad98e0fc61c5dfb70cf90447ee884fd9501bf5fcd1e9b5624cad26cb5d336bc314ee42db6559fd16b0e64c82b5371400307f997c09b03875d22beeed8937605ef879d54186d2dd1c09fab2831f6d1df4fb8c9b55068dbcf8ac505;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ddf99b79582501689187b8ff4432379a7ee6b036f6d475e82fcfc37da77ba54d77d001da3591f290da28cea4ead087474ed88b771fe41ef2544c325716a1602410ff1fe8c43fa627213b284ad8a236cc3a687e41cd6bda9549847170d4446a35530ed53a74a1b58c5a61d1d235b7d939d468a965931cb7ad3393ae1685f607f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haac3824316f6cba0cba466ead38718207dde805887620feb14ef9b38a62e2e00d44daa4bf11f743983cb26757e368be826f71b29588f244719f890ddb1e4561c76ef5943b7c5bb7f0803c6aaf138138ee422b5a292e5f615aed64154399d59e167b67d68bc9c03728d178376f28e568948fa2f596a2df0e18bb650ee4bbededd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7649306bae00169f31af9bc11dc03bc71dd8afc063c5eae2bcddaf48c0e1d7aab6a15097acc2d617534b251bd6499d61e3e03aa945d613f3b7552103713ce177bc0e0bd37c33f640b02a2cc2777b647e6746df350e01c92e2720a231689099b9f47c56b39e8c62dd9cd4866d64fe9047128cf0d68780e6c28fe1c397d71ebbaa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf228e7249915bdddf7665bedc98b5b834746684b67b54f62ba05ccf2d8ba0fa99c193555d978d2c69e15cd26757d10d4d28074788efdc13b96e77c5a255139c0d64a38b7acf0875addfeb3001c78b5c9044044dac6845caa50aa02a29a589c79bc1711bb0cb499fa53c243001f96d33870f3ed454dc01d7425ac321d7177eac0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fb5bf86fd6b1d6447d02aa0b9347bf7874c3cb5e3ac5f41bdac9379d6c5ce7444f80c944dccb882a8369a472947013059e880d941956277b29250005b7bade430f3c64532e1bd349962513fb6b87d1cfd7d2aea3e907fd684e7b9cab9539a0a992dcac95ab57d696826ff32b9fcf57e61214107883676c9a68255835c3a931f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb97b34d716ec733527bfce52787e50d7c26844aacf0b0acfbfd4b299dba34ada4f03bd599fb5ca0a6e9746d0b7fdd3e46ddb2480c3a9fcf37a2c59e46d765f4c23e06f957b89d071f495ae80e4fce774ff9b40e0204d17a509bdccceee87decd23559a9cffef408512957242047f53ec5efa377a889438f1ad9a86e3c47331d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73e49e327decdf17dae849f3924c2719e6d00ccc1031f6be2e9d695caed25530cf068c786a5e4412cffe3ccbba410b5df3bf7d861cd29a2999b5e52be2fe9b9dd73ae116d1dd6a1c1a4e8013e4f4a7d1b7b09155df6a32cc8f596ca4603fadc9d7fe217ab5bba29c12751cbd7958ecf0e85a5f6d0d1604f3a5bb1b6ec71bfb4c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc02f9aae53ab2a8e8d7d6cf8009dc12499723529eb76e4210eea64e15f3c7ab2a5879c8e32db9c712e51773c54b0b196016d07ecbb61968099dcaeff3e3e49fd57994a90da33fa366ef0c0dca2dfe291018f726565ff1b86301e342d6b6e7747e1ccc07226120ebd0cf5d043f8f7b9f1d118212a85e68ee996dbece941ff6a0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4df10c83b7162dca8ff2bac472b495a8d1cc02764c5d95c7422b12ef007a5ebe13b33d5c4727643fd442d3facc3afac2185c60fc3c84ca9401f9e807d6b0676f3b9ab885837b987e41235e14f284c8442026a207d6a367ea20bb1cc4b5485e467fc6843f5228ee7a73f24bb8393f059a01c23224e30556c033d24c72e122f761;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50ddb4ff790ee1d0f9dcdb82a44a6930a0a4998cd00313840dab77306350e5a1e78271ea8d094ab1cbe0f53cf6af961ba166658e27b56393d35398d77cf07918e0937da3c8d4e7025ba8724e61b5f752ee28d0fe10a072818b2dd95024c6ae0815cafa61080b72d3f5e17f1eda292d23bac985086e4251d5e2fe54142972f1a6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7c8c0cd6b21aa8d0a54c3c0c0c02b0a2729f3a8c82d780e27b30307c517d3d3efd885476449f23631495613e8a40f11148deba666edde6c34542f4bf4e869b1cfd958293823f81840651d09a9b8cc0b480774f092816ab139a9515552aee2feefb7f887a721dbd42bddc12d57e1d749ac338cac8b2d7a24496c6cc0b4bde541;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7076efd5d2383c87031b240585ca59f1c0973a8faf8c76da5dc689933a279b3a0461db4205b7167887aac2757e3cfe39a022941aed93808ed6957bef191c672090c254e0b7dfddcf1c07e1cc58f200336f0e2a499f68383e50ef1fd05b12e719059cd47e53ab598152f22a6bd69b87fa281530f849b6d1a5a9b7c8af90fcec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb4586515920c6c3725c45dfd6066b6d567cd1066f382550225f59b7b1b080beb0b6facb45a0457cd0c98f4cfdba13009f89612435ff095f6505883f2d1a006d60df1f573e25c70d4b7ac0b5077c4c7b4bb250e725603b2fa1345692a7e790b920f39b4dca0187f1584a5231a8a21600a94349ec04d104c125fced97993a4913;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9cc709404a3827c47bd4db75bd79f6f0bb8be2cf6772a0d7cf07ca3dfe6c4c90a779f2831def4faaef4fbc59434e1cd31c179cac554b732c2859599d8b7ec832d78deb85ee0738a3ac709f78e47360206beff650728e8592e7bf7ee707da447967d8401b443b085be570c398024fd7495d268219e084668994e207d57c40b99;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfaa99eb65244bc166e305382ccb52c7d402e4d6bb43198fd00fe7c96640560dc637212fe90ecede2e59116de57e321a41880737926b2b12a51311a7e62cba6d55d5f27656c132435552bc660e605af87d03daf38e74d60b581619f4844f5c65d6080d6652dd3578a30b991663355fe99fd0c959e557fc4f3ebc83a884a8f6359;
        #1
        $finish();
    end
endmodule
