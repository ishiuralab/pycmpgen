module testbench();
    reg [21:0] src0;
    reg [21:0] src1;
    reg [21:0] src2;
    reg [21:0] src3;
    reg [21:0] src4;
    reg [21:0] src5;
    reg [21:0] src6;
    reg [21:0] src7;
    reg [21:0] src8;
    reg [21:0] src9;
    reg [21:0] src10;
    reg [21:0] src11;
    reg [21:0] src12;
    reg [21:0] src13;
    reg [21:0] src14;
    reg [21:0] src15;
    reg [21:0] src16;
    reg [21:0] src17;
    reg [21:0] src18;
    reg [21:0] src19;
    reg [21:0] src20;
    reg [21:0] src21;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [26:0] srcsum;
    wire [26:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h244a329b57a9debe4670c705fabac77298ae79e31396485fd5f3dd292660eead4f46b2224daaaf7c9f1763fa9efcf66c6ab419e2cde86ae3daaa259;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd9cc11af9a204af8def37591577442a0bf6a0c6b047618de02c330de8915424c9ff59065bfc87976099aefc56122f1fb4247c851cbb75463f195083f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e32368a9517e41a5f62e0c6404e6027b9d980f81f8e39ea337f34ec695985f57d2305f74b8d8822c8ad1a104f5dff5f0bd56c330add0fee4ca45ee42;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab2b2191de8d737594d6af7c4d480ee2e5ff2f6f3273b46c239976b73fa47ce9ddb17d710e2be7b574eb5eba1730b3f84474a247783835d9ba8f64aea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbddf3469c60f33cd26815a0040334e1911ee14e9a1afa3b863b9759fecd8a2294563845daec8cd0bc22c8e8a97afcd6333de0ab6d9e3350466346f82b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4513c97055d1a0ec4716ce9624edf309b7def257c6e54f4c471b17992f23e14d4ec3c6b730e0b49476cbb4f6c74db8ca19fe58103e3bf1da03b692f4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f0815d59c87263c9790a65800d4163653694a679b86174e5f5811edda181dd570a4600353c59a2ce5a0f42c44198ec0be9a57a5c3201767281735fd4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8098f64e1a4b45812cb5c03e2b692a113477ec8e8e585e4a9215717b9ffbcc60d92f28cfe6e8e57d89e85c324cb630c8a3d4616c9e69e3c55754704a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98e92280ee6eeb8aaa53cac77a410b29a7455b880e67f8d5992fe0a5bedef6019705ad10b80cee4afa8b116892b9ea255c54398051caba5bc0d1fef34;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a9c10e507e971bf87f210fd923309551a1403ffe0682ee896072aedf756d0257cb0b55e791fc9f3832156707e9567087380e1db5280e26bbc80945b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a310948a307bc122c9986c4d0811012e85f158df5e008a217fe9316b6540572d81dfd7e4f53b93a5c77cda9e8fc5ed0449c6ea21386ceebb64c6226a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4a0fcbdd2173eb5b6f5e9298e22567764f771afd9e05f643005956c9fe97da140cc69a1d5704468ba126bc6e5ccf70ef9693cc1b6b72eaf8dcce157c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f7cedd3f79decc4afcb4206e083ef5693ff4284ceb881adbe1b7688764803df1da80032bf586915194d82431fc6904d45f6abc00edc6e6a04f80c846;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h249a8e9670acb88daf53a886c0d57f0df157ddb3af01e94de90da423a1c665678906017e977234ee591a16653b58b08906316f49afb9fdbc64618cd34;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c08e1e3903215716a740b69fc089c599b0e69bc825f5bc754de0c12b718c1b3a36fa97a0f02471e8e397d42dd6f73d2c22da13319262db2df571c52d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e64bf4ace394b0ceb8b8ced1f8a03f38eadcbe61c0765c6864f13315cef8d68a8f7e8f772df744f799f916ffac4ffe0dfb9178f770df52beb9dc24fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1c16bd346dc952751541427aca3e6a126b6f0d5acb07846f5b5861b18138c5af273070277c580c25e71f81b795c71c55720b36d4658657f4579312e4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b0279b997f7b5e684433dea961435ae3d7755619d9398bb06c44fb5b20cb93f65347413bdafe7e766a6a307f74cf88e43da6a91d0bbe1b2d2032700e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f515961d60af0598d85e5a28871176ff36acc8a128515d41806c9e6acc24cfdcbac2da0f81b3269d17fee9a00e32db5e1e5e6a5e2bb2d446d79cc17c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2f1728ce133f176566e07d12158d5eee70637f40ea5115d95d2aa1b55e46cbd2c6ec1022828771d8056c957f37743c28140e9a80daabec56c1a31f8d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d0ebb01d0b8bf9ea182c7144e2e05a61fd1e9172c963af9fbeed96664cbec8d46e6035b3ceb1b72c27724415215e3c77d3b7418c46baad926e1e492e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee8b930b11b32f8ab31637285926ec2dcff105ec32ed4d255007c9dcf8985d624d42735031ea8b51cf6bb90388cef7f61cffd5f4e4855776ce3287c8d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a8330f1243eaa9f06cd9f710625ad04ba53581be393ca91989861c075e6872500f352a632a3393197aa584c915649d32ea5a72787b4e85d330c05962;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0e142f39ae0e8e343b80f5a014b02203ee7ed9358334c7768a86cc6dc9debdb00c30c8c18e6e32757846ab87e30644706d4c2915637ddcc83439c2ab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69f071e5afa6c75df8e0168cd2ac6e8008ec56ca7e0e3179ef3546858c49ae49eab0d6324dfa880495869acdea32051dbf4822d1f263f5213913f9a2d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb315cfbaacc9a723f44e77821a42009a0a79c3548e12050e4e7c9190e00094f79d8c2235bfc1db0fb80e2e618916d0b147096595cb3f8a0802d4d13fe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44d9d7a4580bdcc33f2234ab16884137d5428c227ef13be2023823f1c963491fd88074c2670ab9f78acd2855f24d1692680946159b3afc15918bf5a29;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91e145d5abd05de18afadc2721f09a2da922c29c7e9381c6830f6a8f6c331bf356eafe2321bdee07d014e7ee65f5266edcb63a43bef700eff4f9c2717;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a2cb8d176ac98a2bc4b9fc4694ed715f4321ad7c87627e36a37df1ab6000b509dcaaba38162bb39d0af49afe626b91e256b689df3057770d8959b005;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34d06c3d8591f050ae05527fd4cfccbeeb451ca0762d0d5d4095f388bf2b37f7b5c3b02874d64238be0d8057ccc8360ad34a3cde329fa9abb06e0bda0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4cacdb84ea83425385c57e158cffe39399c64f0ede8ef6287680d88f13cb266157b5d7593660cc9a0d457b16573ae19e9d7d73d91691df879a74e51;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc083dd67db33db4add3ef5c3a14f5560bffd316d50869bd82632846da465806bab1c5734b0e1c6231101d0ef2d622975e53b83eac87fafcf587fd3e79;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28719c7e29086e1873bff8d6179342eb7f83f738aa085434c58d56443cdfe5224c9495f08c84fac7aabacf6a5832c37c29d7afa9170a75c2f0eafe679;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1635f69d8ae8a4fb5faad4d8514f337a27498fbca348c9a85c804b05b63878a6115de42fb532027563388e4c124ecc97eecf59793b5a5f65fb522dc0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fe2695c9fdd526fc3fe3d5f9585e0dc021e897cc1776d9f8502879d79da3890c0f2806261749897d708330736bacf75889063aa85fe62f9178d1f53b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc529047a8d08fae806cf5f6d34b3ffaf33a8740bca7b649296105fede0614820cc24972f473181a582d407713a57c26cf2fbd8c2dafe88501f370f72d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e4123cd89fde86859ea5a573b300e7a59c63135466a09781413d333d339f73ebc5d0e8fcc2353c0e04d86fb12a5ac05130ca5925dbaf225e1bcbe9e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8cc5d191f6747380674b2db6a5e1bc6747ba3eb22995be12e5b2169d7ce4c5330e6cec89bfd39b70a45452a6db2a956d66e8a6845164dec35186fa418;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb626388cadc4d9220a25d1b2e02703b4c2475ffafe530894196b306828343cf2fbba934036e7b4a3b5649927da7ea398a0f92442eee6e91fe78a82888;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98945f9396d34b3535045c2678ecf899b3715aa21aa1a7d1a8399871ee12a93a60322f022e7415180e3367e04c5d2d817b9ff1792e2d2c7e0df55a2bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfff1fe5948f268ee07661e8a2be391c50a2ab28b781ffbd3a94bc25aafaef6bb486a766aaac623fd06ec76ef3313d37c1e3216f8b1f3d244f6a9593d0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6bb94bffc4e0d9fdbd58f82a6343b6b35997fda809546bdd715376581f4a7f98e27c910e6cda0e6bfd0d242d50c0476bf6c416a7cd9416272912166fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c1d7f379c603944e245e011ea3cd51421ec7745d327934a2fc6aa6a75531e0a1946acefefc48524c2637907f587bab4b1c9e2db47c7bb7a2232eefb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h662c8075f86cf40393adac66c8d3baa127d4922bd388e53a197cae8c85067953fc72ee527de11e2163631b8ab1d415b0c6b4a72876b50f3c050a94075;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f350af640f91e53cf0338d5cf0e5846359de86f12f71d835d7a5585ee8232dfc49dc6d8216333eb0d98a052624018576c339adb12064be85ebd1ceab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6506d47e6b38d846c46f0abd3977de6b47ed6547c08782cd1e7440083efbccd6eef3ace62cb28e9f8614ff5f392dba7be80974dadb04d4776e4a37c5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e0c06176620e966ba2f3fa60f10c97ab2dcf255c11d2f0870c0d6b2ad8985c9dbeca3d3ca93f6f3c0733f64cead70c00a89e87211fcc70c28d5942c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he857f6af7e887c1d7f61df928e9b0cda4752b5ae41a94fe470f667966074d78735eb4d448ccf85c8ebff296886f18144f776bb3898385faea49299900;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3244bcf22773ffc669f8718576706fd60f0ba51caa093d610a65a581fb89d42ff99a9a5b6aec8f3eaeed6435f91945e740fb7e6495483344a1dd852da;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce60e23fcfce45213e0bb37abcd1c7a4ff3f2495fa9001b6e95464b8660c3afbee0ed0b3319a23fa1386df707c47feecbf9b7bfcbd08e518b1f5a8300;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e279af8cd858b8b8d1925892a35ecb0dee82097ccec896238ff36ab9d3b49bc5ff1ecf9a28fba6cb1a0ec6085c7891a7e108ebe90136acda621b5fdd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bd0329e6f37813c6141730fad85ffd124d5d66a30e53558bd61c460c896a3658555a11de28ecb6bd9b727e7f8d3c681920172d408be61cc9c339cc6e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfccfac79765d8d7de02d69cb2339550195e3164790d0127600af2d9dd703220306d8ca88f29d1ab6eee3c5bb4c48d7127fc44ecbce0f0f2717b415476;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8ef615e8a2f528db70be7a3d7ac4e2147b46fc0d3f274717b9f041cc3c21f60875082e3a4d28acf5065f83e1d8771c79d2727e7876abb83051ba8db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h188387153387c0e643fd27c4a27f47fb08bf8f957f31921d3e807f37961ecaae26a75da49784f47031b88658f088e769606a860d98372d30559112c91;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bd1de8aa199b90b5a78d9b6454e3d4f5ba5f6f88abf7ef3e90a6540615f302298089e1a995031c0d2735681a7543cdfd7d0d87fd8c62506e93fedee1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h970bd56115a0e39bdfab94558da6abbacbe287b7e85dd5aa459fc92ca149311dda6f8981050614066fb58fd916fadbbdf01e71298bd99997565905b93;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4dbc2964462e473948681114e7a5b9966ac394466bca30c7acc2e33a4e1dbcee95bbc6152e7a0b57a3855c05ff8f5d34abf9afa6afeb2c2e3180a3a39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5797b35b2bf6c24af7b0eafc7ee410bd0e15bbd7dd3def48fd179d41d602f11d582514f4f5bfc581bba2c942bc4ae24c51f31a7ff50eccdbb17b1cd56;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf51677e78f97935bc3bb5384e44b5fadb2a12d58c7c9a7ce7a5e91b9f0ad7ef0c560ec0935c0ece169911df322cde12d3f94b6b57d2fd4bb605887a75;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0c2fe89c65e37dbf51a4c38f4c1bef8138e7c1c1edb7932585347cfd5a0759040170f34269d4e071d36b427b9bba9452af86551145d3f15620537621;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf068f5a08d00aaa8f522f3ae5858aa6af07411cf818c01ea234fb75328161ea77cffc58d334c457bc40b3411db2cfe0ba284ac9c1098dbd4e986b7e47;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfab939eef327bf8bb336336391fe69e1d8fec02fd20f1119a8dd91265d09dbb1fa7e78855537e3da2d2d3f9c06b8f84b4640403cc6f4f2f3eb9d82d95;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8e8e3b1f3d8238a2400eebfb566c4641cf5adce0d5b1d58c278ddf5403ba0457e954c9fd6661a8f0fe93cb9bb72891e6b24501e33274ec7d6f02a82c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8fbc32505309e5a22b3f69116a0edf32dd2059c69ed7bb318951ea6670900c192fde3e8904e66f141754970fe16078aa554f3c942a81ccbc726bc20e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e3e08b78da963752b2f7a307ce8dfbbfccd656f444a5b5a8ab710b98392bec009e0125b5ba8cef74d6c5aa0a88145dc1684fc4635bfbdc7c4120f24d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a13bb34befe0fb7fb2216126adc6b574862ce8386b2da677cde96715dca4b9d8da16ce2c997cba8f08ce872003a86bebb9648d7cd235a5e816b6c8aa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed89194f9d49036d03fee827a55814d4bdc2b433b674b00fd5a032485a6fbd22a4bb555ece5756feafd77090f3747c9a73b71fdfcd10034e75fe4d2cd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65f998d6769767b9a92ae116c28ffe2d1c57f1a44c57a475fd35ef32ae77e1a8b186e1b8d181c7e6518e1349bd491eeabb3c03fc1084fd2ed4b5131e7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h953c76482b6606175e08ff536c616feb9f04f5fe0fd9d964076d0e33b7751f61ddf82747adade67a331ca3ff42f0e888f31fd0a278ae8f4b858066911;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he559188ce174b393a050db60b5817bd100b46d46a4c01b41775692b9ec9c2895a0a6115b75a2a94c5bde1384cb2d1f6ef58ffe4aaa44da3b240c1e04b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0c6665ca5942be15834dd3f8699da668ead31ed34b6053a2c77aee373274a0b8e167c887d150c1525207bb0d9866d0cb8c165e33b24001e27fcbf4e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9c4aee0b9d483f45bcf204ebb74acced27f1e0adf3a7fcefca1c1a7903a90502ddf9de86546afa3dc20998f612e5f6df1f010f18bc787ad83d26d4a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2d36f4f447cb779a9c108d818251f0856cf172486d0213db9e3f1cba491d548ec766e15062c7a3dfa379ca993a2cf8ef16c8753fc78559e31e0db2f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fdaf57036437181a42be687fe005b5ac4422f7fba5dbfaa50df6f68a1098f57ac0580b629ca55070cd27eaff67d821b41dcad98408ea216a526aa3ba;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h967b3abbd67e60b5da0c3068b4378cea1fcc1410d193bb18d81d0f1633235fecfdd711dbc8096d039430d0b068c55757612dbfb3ce5e2b2353273d6e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3121e480a69f30aeab808d62d9c13f5cbcf95449053d82b2e30af70cfd18b4a75b3ac929a77c9bc2c56b20d9ac294331642dda1c5a59f3d8326749656;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4539580d11a606c9183a524b11403d425ecf01378af230f11df97ee9bc108589e489de58d48f56d1fbde0077f370ce8dd2fc904e07137a6baf1b32a10;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h23ea7ed6be9bdb4fa029a12afbecea69c299f2947048127284afeb91ae3e9a3293a18db853a504e50883f293605c82b90192647ab80f4beef01c51141;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe916a3dec1dcfba46b2a4c441d46883620e1fd43c3b420286cd27d208b0b357d9e029d4dae09c4ae749e405762274fe009764c0a048bf7cad85007a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9524aadae70c9ef29e323d1f17d43d8c9b42c0fda6050bef0b175cf95a235d0a94ebf05fd87580180a7930d403e750a145745007a1916daf9d8c6fddc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f5095b9c23dc17210420377b8db04a5a9076f1f5b046aa0233137fe79b98a69ad6bfa2d68c4591cfe9a47de56079c52aeda1b32df86e07702be16ac8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa677609473e4d11661edeb4abad074a93ab9996a2c8d5e943b2b968803e3d2be8e0ac7b424caf218fd6840a1706c412957215fe8f8f72d2c98a95c90;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac1ebba936773a0666c5d6b6486972988bb362f5254c65a490896a7953e2399d4db6e43b3664aadd9c3cdd53b1e7c9f2dc402427b3023916ccbc7ac4b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc2940564b29450455275645c4324bd64b525d0f7040c24d3f8d4d1d13c0c758747a2d10c9ff90021be3ef346057275298b2e1147dc5e65062e1170fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5feb6af35d35c6dd1eaaef685854a20f83e00883a4066919e63aa606c97654470d68f4da79477ce5fb4e489736ecd6a280683868060df6cb3a6383eb8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2722bba0a7eb5c445488269cb2dc78164075e364164b5eac4d05e67d5afef985a0b34acdf86bf0e45f364d29592b8605876240a887f729968e7c16116;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha78fb09f61b911673ccf7f4e42db9936b74a6067116d9564be390cddd7aec5951be141322f4e6e16f9843b5d4da002169d6d79973c30923f322ab1063;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h871ff8f311e2c61b49f35a175011bbac57572a8171ce3c4fccd37498289e1c1d80402dbf58493f2b0f7936829823b4c5308e8ee985fd146e3d81dba00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6981baa1fb09f2795712583a2ae012b807e52201334e01f7515b297aefb87275ad4a9d9ebcf418797490dee7d47487b0763dbfcb423e01752d1d955a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c9a643c7e7b5b6f73ce4545160f2671850dc41e4bb8ad56524ebbdba0a54b0621c8be06201ded062bfedc90a56cdc8337d5faf3de2c95bc5b5359abf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8aee922ab810aae51f9662c770e062f1e98f265135568fe586bd9c9fece2684da72b69755894396a625217ad5e95dd7f33653350882d5c2438ad5cc7c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9cb2299f40a6493778dfdec6914f6d71d095857e79b6195c8094c011f2185c1e63e836d153574519a0929fca0ed5d6f805c861905928025c9938be846;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ffe400e9922f44491a4b3f6081db4414c3350f24271791ecfc64daef3a6d863993b95ffc0c3cd09acd0236ea9fe8d2c8b9c062ab6fbd1fb69cab0268;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb603b5e21d111b122d1c5443fc8761467d6085c09ea227790b4ff242726f692f2d1c6096772b8ffd1444634b6fbdbd80f83976e979c122c688877513a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2e98a658d5422756f4e7ac06b77e8abbe33c7bf6aae065d337ae16753f37e67addf0be66ba7e965d54a9825fc013e1f56cda6f3540ed4362772c6340;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b5f13ad459ea1fde56385b24e44cea10a9b80b90f84d435e93c186e5f8dd416709a88f27e2ae1ad08193363ed620285fb254987b51edb0a200ef0e60;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h802a8b43a80eef75a3306b0e7b98dc71d65279f22c8c0ec2f4c4bbaf2a43d368ab2ec426565acf78873c4931f351d2f49978642774eb8f2e835d3217;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2d8a2538547b51ec952eff601ccd4ecc59cded9971d2f444123768901c7e2aae809fe09387a02bd181dfcad33db68e2b025531cb5b85b772d32edc42;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9251c8e557b3d6b0567e79a1f4ba63726c47f2e11c90ecd4d334b3a25c28f8c4dd6fc934e821b0d5c9fc3a4bc01346c7cc1f45052c09ebf4b529c986;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h481b8684213f9f2835422e4ae6ccd66345bf04238e703daad50dec2f046e1fb84120f99939058dbe77b77c43df5a1bf06f6289f72a4490a307c792242;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf45ff050d588a3aee74389e1c6abd118b9c1bb45e5c461a1d63da2c5106980d3e162c7cf289a56cf7d2492f5e93df6908e2deaca4c35cbe74cb642c2b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9a680834bf7fa557d2bf238e7b566fe9c108ed0ea562be45421e1addad1ce0626f5a9c91eb62b36097ea4e1a3a04a25ea148e60f5b54ee01c3fc3b46;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8287f7b352fd5d1609a73e6347257a3560ee3d2f9af02a748dc3cbdecc900b88192fc09ba78f8270d950c18ee1559c8895626960a30e50dc0d96e22a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a009a4d249b4273b660b738c29835478a8d6ad7bf0ef68e66deeaa040c6f09d30c9287da25a7628f50eca180e366df5e617806554dd0a795d229bbc5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd41980f4c156842c95dba6e3e5101628d274ae5ec89c25536aecfdbed57228ce2470f429967d8312069dde0c4f6d952588a91dc75a179336d3b9cf845;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b7e50a2c2ed8df1076de846ce964ff5c464ecd55dee52b4ec9d634d4691f4dd6073a19fbd7cc6ab063a0b1745a68e145fffb6e5babddf144cc152324;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5dcc6a67f143d87da9eef15807e00beffa560f8c709fe14adbe9e862238a91c0ee6485987ff2ed4433bcbb54445a66ca64804a4ef04d1efff0a59201d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c2717941ac3bb1cac977feca8229258581c09c11bc10f0fa2e71982aa618806ea62b2f5685d5e138d7fb2cb6b661631fa5260b5c99d1a55516dc8277;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9626da69c9e3b4fc55c225cd8e002e65668e3b107976beaf7e9e726ae379c1a06400d2d406da7fcb398393ee96eef92e4c67a345742cc732e28f8ddb1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52cf5fd3117f1f2b47d5a062ae618031977cba230baae7de56ab2822b44c375fc97b9ace8a7452c92c640df1c61e76aa192ba25620e0c845f190ff3dd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee8bd6f361257ceb59f23b883c8f7b9572bbf08ef05d3afef5357efd1cb1bfe93dd964932d2798fe6918bc9008659557f05aa94661c40e60e349bd614;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47f74a7d2004cf2f1d97761192fc79342032d877624ffccfcd349a056f36d1286162605fcf2270d5012f64b5cf0a812920c88bc0f983e6afdaec0bfd2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc9f24edfc41b70281a9f44b03267c43ee2c25f06a7cbeb38519d58b260b4c1091dfa6ea705c6d56914b39bd57213fb8d133ed4a70acdbe2dbbaa173f1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45f2bb5ff77f9555932ebc450cfd364e073d4ed9181d18c82542d5faeb3476143abe7e589b5fdc421ea3d95520d2f31630eca03db8023d1f7ffa4cfd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h674fbe72a10e325d1e0a17e19cc4e6146627635ee0d08e3c928db6a2169ed6527fcd72091596d5490e5b81dfefd4a0e054aef262283bc4659e10a6d91;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5b2f119360d38f2a7eef1d8f26ff3f5636997bb5db2ea88240705a6d7fdb6ef1bbb20c39b9b80c763eab3523ee2adff907ab96862df96799270dd457;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58be3cdf5dc4f2d01592f72ab7a822b0d83c3722af39d4289845b15a7f8f72ddcdc5ddf86c5ae217fdd8d24cc719e77d65f692bc251640a1a5022f544;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79db153556d7d64bde82e39b62b065a5f53d730a2a1ff33688c904f421ddfe77c9beff05d19bee683250c66097566890286037977fe2ad2a686a4e7d1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67cc8a9e61dd56d630fb3091c277d8bf26f66fa7115580f5d9f69c8d8bebd569a16faefd41c353ef0c08937dc11740992820ca98bb1980002547d481f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a301bf430107209ee728306449dccee6045076bc828c2341faec34557283e0ea3e59e5bf0a1a536085262e3fc9613c6c484bf10ba6f3e1efddafdd26;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a79a77e5e7d25777f7fefa1272a379b6c22f560c197e845782c525fc2023ea42ee302897b0ff585ac001d4791a827adc75c65fa1a361ec329293c3bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1cbfedde5d93073081dcbb951a4ea7a582cf099aba0093d63287d7e3cf57e4002db1c18d62dd70121fc017bafefd4ce079d7c791bfe3ebd8c370b061b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4b2608d777f203f287b4a0e10854387dfc90d9558b517140eb35ca68925ab2c4f149e8bce2cc4d9b5ec8c8f906565a9f41d04ecff2d7781b0fdcf7fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46add792b099db108b9db4129e32b92061dd8bf254da5efa742867f4c3c005d54fd269b0ed74e08b92bb923556683e54b07303857219debd42f3e2ee8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf65a44a0f7d30bbc81a31c0dd53ce906da88b3e2e19395a85a5b7f6f52c9196caa4c81ebb6b2f0671348938fe94e0d49e00b2aa8fe84461097fd44c0c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63e1d31742bcebcf8e5a8903def44ea56326e46b6c6b59c9445194ec00e01542c84826427df50920e76260407ea1c0d66a68866796a8cb60c465b38b7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5781c222a3912efaecd175e989294fb8300787c5234f8a1288508d79c214020404c8f061d119d0cc85f22eb6275b690b600cb3e71fd29d3d75de9aa5a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86abb083d37ff6ec6af87c2e29e11b02ceda4703af459a03e5d980f4dcd6cd3af08c2db362d43363334f55e586474ce605a3f732695cc49dfd2b55e8a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3de322d26f0059d76cc76b816e7517e1aebc39b0ccd692cc6f6fb5ef4d30047b39b309ce3b43fa17b521dec616bf712fbbca60e9b3682b793610bc66c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b5eeacd2ef17875197cb58b579fbac21dbfb4de8ed9e3bacc4dd6663cc7d955f54db03f59810a91c3f74accfc08544af39ffc62fd0d9b4e3c96474a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd116d742443aca2cc93f394385bd2136367ab522cbff0d5cb928cf1fc2e8e87e6f9fde330c2c74cf1e6d5f1f6122cceab75d6ecb374e80519491c7d51;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h158723a115e569815b3bc798fdb25f9ba84a3b0ff81f8fcafd44f834989674b595dbd07769e1d45ba108681b18780a2e80d4942c85b594d0622e49b40;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hffacf7cb7bba4e88e008bbccb95bfd68541cfc796f25d05abb3b35594b8625989952c59c70a166576dac625f757e18f29f732298cf0d8ac1b144068ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1709eed732c5e0f7dfec54dfda80cec8043ccc3f0877c307463efd8a3938490a3a857e6acaeb92718f425e30c689234361ef5b3cdd1f007abe81c435;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a8c5e130e5a47d6e51ebd9cc2b75307d2c02704ad3135b08e24fd09e5fa62c4cd7cd1e761d0d4e81ab1eb19642a7648ae101764f54a981eba5ef4f1a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96e703d34dd086f4e8e292a24d3e549bcb35b45e0fbdd20237152450e0612c348d62bb85947c0677a00162e359f62a6d12f693f18eeec342b75d41922;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb885b47be0884010aee7d779db106421f1f64942e3629cca62f8fa3f726a1a111d1f49286f2c79e5b68bdcc37016560f2dea8ca287fb5cb0d8763e45a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb843499dab24a48fab754e3baf2652436f7d04d04622aa67cda2e61952fd6cfbc2c790ee12095ba789764c7a81173ffd2e81105a500c431930267a86a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c80eb8484f2b7d8e0f1c75e3aa134fff71fe062b55bf436b4d6bb97aeb079999eccc68f1c36b959bd2b4baa93c3001f9b05b581335bf7f14a4aa7870;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8aadc33035452355be81ce39c025e614995917f32bdc4843e1f2f5fef544fe3c65cc80b67a2e26433c1777fb39b29b7bd064c12f2a39d8b770cc573;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h977a39a45c8b07ecf983540eb580cbf558cdb339d465731b8f9dc777ae22c22d7fa312fb52e8a4bb7c4c330d31a91c70019028c66350801141c1dd404;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71d8ada9959c6523e6ea4c72915ef6cf38e223573a59cc98eabf618ffc2f49dd6e19b85c5147b8eb8644bda8fdba06e61a5e4456a9d6d4a6ec14faf2f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hafcc492fec7ee161ac9fe8f6fefd3fc41fe73d62a42fff0ffc26e42531e68bcd26bcda84fc3881b8f4c876980ee7dbc887abf57483c3f635314a8dc11;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0517d6b9990d61774076c654948a0371643992d83380e06ec8b2b536c3c8fdad2699a8643e979df63767fa9bd9892c867edd3d57dd0c18873cb69ec2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69db7a7fdfd05a0eac587c2ffc60b72c05a9c27bd30f28b9d2d6b2b899f0063e221c471e65f5929fdd24ee8c8e53d69bdcf2e69dc988f699832ad9594;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7141d21fd8372e8b113d35c3633298a7eec49a531ea840a8c129401f1d4aea8f172961f59ed4b07c1b710bf3021f9f9f185a10a1577c2a840e40dacf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d0a4ddb7fe937d48d9b87c5e301057bc2ad2cc6e853c0f5fb97ae93bc3c9f181ec2d951412f96eddcc956b8c352f98bcb357cbbbb3eb9c36d45f3dc5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5fcb63de8264426d5723ad557dbeed613bc8631e0d77ce1fe4f74f005f97894368c89ec41f27c319c810ef464cc5f7ee7450a2e50d3ed5a54fbc47d8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81ad40f9c764465d7149b339a99737184734be7ea6463e8714b8abee8378c42b289ac6496ddae3a136ee132eb3f50ba971e7e05a898dd6db500e8c733;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcda06130151420500699ffa2b9828c472eebd483aa361205095cb4afb9ea7d15f66b7871a3d9b7e7577dbce4165b4bfe5c07a2503e562861881d8516c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff8165cf931b7cf3d91b40e31e4f12dff5f838af17f69b5052cba522bd35e74125245b2b834228879c6f7fcc3e1ce6a8db5c7f661f2f58224da88c8ab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7494b31c8b51b22829713df50a18524a46f251639033c173b3d81ab0885e04de0ec73a7891900a16772d09e3b9d7a1ad83b60d605bb1d3c8c94d9c127;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6fe42013110d9b5ba382a67e38009db5a36f5268edbb491553f02ec724c82f96d442ed03587c57654a072bf5d97120027dea0a13902d75b7bc49694a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf8b491ea24c31e5f733c96b1bd198520d04a61a83d2e8bbd69b49f4f7e24e708df98c491b9219302a96a91e7ed95fc598c1bb9146e5288c09e12e646;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4be2e80f6a5bbd6e49253c4d165fca3aa747494545f7843c204f0c4ad209a56c71a9300ddb8f6fb13690869cb899fbbccc082616d0d94493cb3548739;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae0e98604ef90da945552d38439d85253d3e4512c1bcf4d50428ca334303a7cb75123940037bc3b5f4feb82c3cef97b9a15e26706362647d0bdd7dfcf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96f1d2f736280d753b5e5b66f1f742cad8cd61e9274fcb4f1ae4c6d97793cd93ce4ffb151dacf1d2c60cadb119aa294d6958050806c766de8af7e397a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9c594727b076c4e9b5f0f4c8f42d561cc90469b03435b30ecb641daa79e00e16b2e9fbe8bac1acc165f00505896e4f199bda62950aa2bc6a61c65995;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h646274c38166a3557a42fab22d2c4bd20242d74aec5eac6736be7dcbdad460cdf730b4bdbe0954f061a564a08990cbcd8e025e4b409468edd4d7796f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a2bcf860de4f49830b67458dc0df2d57cd32069f2bbc32ea0f4c7f8b2777cdf3adb65f35ca033248c0566e40edaa57a7a129ec1c1abf11e1f32dbb59;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9aa80cd2dc167bffe4cd11a21381a4a90db4725eb21898b2c5c3137ee315a36c12ae8ecc031b09cb2d50d7ede04940b746c284f2226ff6315ba0812dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5d2cf9b8515407ba5aac928b6534066e411021b5a023279432621e22f4a5bdb0cee091a00f89335dbd2c5093f127b354c20d94482f0272718f5bdeff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0d788d8feadc50470162ec077ffd798a2035e94235eb86253ea7530149365fd490be63fc774f20bb81cbfc2c7998d0260173dd8dcd47394501f20f98;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66633bb676c4be78dcf319e28b360a179b19dbf73d936db976cb407b2608cee913a59850d277a70ff96a7028f88887b17a411ccddb2fd47bbfe943354;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c0402cf8a71ebb9d450ea0a7693a87303c5fa605b5dda5a5a5165880f00995d35fab68957e2acc0e40290e44c68ac762239d790dd187061e17713ab1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7d8dc5993f4d76a37ba5b4f6a89036d93be76c407efa33f9a5df28221a6d37e39e8d12c9c4b6ec288dbdeb712b86692168a11e8e5f4ab1881b8e8a52;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h933587b1da7b905c3b613e2c0c5a28d33f61bb50be28a36c74515848c3902d6e583a88eee675ab09756fb0f296f1259e7ef4a65a64815ee20b8785479;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc25cd45d08a956618df991ca2ab3659b3dd0209e53a924dd3ffba070f8ece944e8b32f733935a646b1082d05fa9dde4a2895b283c4d216fe4de19a808;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76ceda09aa9dfe62bd740ed42f678dba87ac6e46f31fd9d2acd2583936336256824058a03ed833c47f0b1b77c96214f0a39925679c6dd8571fc6bde42;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8e1950f92d7b1e04684f1093483b2eb97668d4b70410db1c656e7100de89a95a8dc039fcfa571b22f844908f5e7f16648073641051f8adddde1f362c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94787faef1ebd3a129483d92a566d80f79902d5776901d4521c2e782e6df4dbcb480116743fe116320c8c1098caa0ef07797d5882239d9e83273524de;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h434af19b00243bce41a7f148ce9405e5753b7b077fcd5fb191d7c551bbb90f136b45354a6b97cbd5163974da2baae4ba660ffcee9acc2e37ffa18b8e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5b6702de720a3a2f7420522f2d741add7192be3cb6c4d731b194e21bc867df739203d12b46cb287b88eef25dadd88ae2a77703b299a38af9d0c83efa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a952fb25b50cf9beebc8fd26dd7535fec640874b42d6b4cde51fe104c23f4db1660f2417bccd756d6456ebae86194649942897f01e8fa6dea1719dad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h579976a7c969adfb10e3a2343cf43f6133d266d4ec40ce8800a660acbc14528390ce3bfb48902d956b760b139eb44d9b4bbc2a7a103155e4826c96573;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h208e6cd038a396a5f336cf6ca5340c50681c797c429faf1b77cd116b4bff34cb3cc561113268f9ded3fdc8f8014770b3f3200ad4e38f25049dc3af22f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb170beba5da408caa8011909d4763d70a7fc1f7d270d540aa4dcda5638d7adc0faf1726989c8641d5fbf05c290c065df989287807e988384cfe0341;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c8e1f44a7f73acb21ca2150b93f01002a6ae0014fb6912f8d2011bf0b2cbd24912f5855dd00e3c81533b01ebb4724f124389235d521326b7db4a6aa8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ca4d9a8d283e66919724e9e6b688a76e7569ff9a7bd8ccbb4a1e77f820a244f0107aedc5b9ea1635e7677526febe0d3bb0ca1114e0f2702bdf46a8d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc77701fa6643f6ed27a4441f74d18310d0c49fabbdb6468ed1cf9c047e681b2e33629c87d86b0e5e54b513ee867af53ac26dd5e8216e59186cd49ec53;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8891a3ab589efda188bf87bcc87a947d98e0e093812c36f300fb5ba7d7fdf459c6630de7799851352626049e041f2e80b0c2055a8b14be487e455f361;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1369ec2be998c9fcfc9f9bee2bc3c33e6919a20ddef9cc12e7998add0949c9e41c5d4ef04fb1d550382ce678ca16354da12ab8e58570b7c58d18c78f4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43ba29b17b47004664eb1164112d14c67b92e12f8b556af1d3275141f8fc1646684624ba67f8ebe9ac4344bdaaf52d3f0ca51b46462809e64fdbab95e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h531480d3d690d25e1317af22661ec4a86efc18d5843d2649635877bfcd67b611f72b5832d263abb25da47b114e97e6955cbc056748bf429ada41b9a82;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3791aca903e5b3e4b7ef5ef9fcbbceb5e5d61babed41c81455b1e303fa7565c51309a2ad1bd8bccb3d3e261e85a4be4b8a3600325349e3a5563ac2fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6f6b43d2827fc095139bd34b02828022c871c277a91e272d9f5b2d39ca91f947f3e7dc67bee39d0ad4bb8684bbd8a89fb1b7a22a4a03910292b7b9d5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h409fdcf92b1db6967fadec63e1f283926e0effa80a3ce1667f3b9aeca6f4412bc9c7e89d7a01665a86f0cf2c96b3414d3198dfa4ec1d0e33aeffaf926;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h691ede24d6612a32abacc8c0fc70b42cee2c85c344aa17023e5131f239aca7b3e2425cccc7ad7786ba9e4de2a838e26d17382017b718fffbe294f574c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc12ad29736cdd2f0af4411f6f84fa0647946fb9735dde36d754bcf96ecd377e499187f40805f5cb1d70b123815319230c670c2a2c55420e82bd81976;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65514ae08603ed8e076ac85c8adbd3aef003942555998660eeb76b8cb32ba6ac87cf34b0afe1622492317b95b27338734ff6da2e148e14fd3183defb9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bfd4c33700afe1767af018b2d7594f308df4ae4c52672c9856421b67dd5d5159cc824635cbf345b4a05aa1c65f552d2bcc3fce3a4ca6c42b4453b618;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d2fc0c87ee73d1975c2fb6bafbf8b550e62377c769b5fc2cbc1b778790dc3d0ff700209b6cda03bd23c73662d9da6543008530022ea0cdd6d3326858;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cdab044b6883c36fbf7e0b1f6f6744fcc49d0af77931dc1f0ddcd6fa38d0426697f923d2d875dda3f762a4b06ee4c328df986b3ab1a954ecfda8e19;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a945a1d94db9c38aa8bbc0a92217e5dd757f74c020d18531317b1f61443d938ae1f0975b461a2954ab67ed0f756c8da5793c38df793d3d3bfeca15a1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43dd856ece076da4670b7d9555d2983613858916603305b23a0883ba3a2b12eff9c71294ff6670653eae1e6bf265ce4b9dd135b54653d5c2ff2150450;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d783a95ec0f0541e11536c37064334c1c7b445834ef8ea9e168045076ee7297efcd27e8053e3e4b0e13e53f88b00b07782ef5ffed82860ef06c30304;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c2de5d2b62d30ba1036804e5e6e871a433ea7a619bcca476b48b48e33949551589a6fc60a0c241b599abfad79a8e469e4795be7957e4030a5fac0f9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c1b1c54b9f3ff134ee5e844de657c3f3807f6eabb30cb891796b20c35758d0a790d75eee2f95417303020b293579aabbd04ebeaf74cc95179e917d4b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac18f67bed59f70a282c5f61ec733490842168227b0b4edac60564d47050a176e816fafc47d765d53e8496a3dfdf4036f05142eb13fe74bccf37fa35a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd6698679a29eb842b80cd2fd8a1319c8738fc4d5c34dfb14cc320f1aaa99b14b21a46fd4906a565416b98d8458125bad23f4b9796588d84af07019f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42b418587d43049f464026d3c2dc8691faf961776bd29d57e0ae3d6e2a2012908c311e5e084d9e8b591fa08bbd14961eebf643578bfc65d804ed2131d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17b5fa1619bdf51f702978a536c2d2022efce4f7c0ad769800c4703626cfe8e562afe8eda8fc37052ea2a8dfd500b208510dfc9cfc1b71d5c0829b0ec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ddb168b90a8dc11d89b9d37eaf6ad490e6e757ec82ef597a9db7bcafde16d1e5acfc005b5340a0d4ebf9fc6009b72b716be2d4535b2867c9af1abea8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h718dca6acb18df5b9b8cdb4ff0b41de67e8805458bd88f46dedd99017552f8c9dd2b801fde4b4b8b583797545f044321ad9133ec603dac9f1b42aed7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h645ddd59b30285b05f66a28f772534c5df16d96f2a6296c4915ed7dca68606343aada8367e1783d35061d6c266e1c8d4381af4734afc1f1ab2e1b39e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf29b19fa0a0f8d2b208bcf7f84433fadb3cc1571339142049dcf8ad9bdf6e308d35a8c60cb5fd6b3265e28ee59ceed4259f18331b3de503734e263b1c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65bd47dde803db5ce8c82f84d57da87566da1ccceb7ed07b1b8c772bc2605cc468ce81bfc95899b85bd68375ce65f282ebb23e5021efbbf97d20dfd98;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf9b43467568fa9bb4ede92587d54c2d9f4de8168ecce5fed03fa813d349d5d6f8b4a285a64b410e301d383c6d6962a75ebac8bdea1dcae6cd1ad82f1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b56531c3d94740c411ab3420aff5b00ae68af687e608382f3ee044522d07a040cb95c766b1cd9947b96346a8f2c3e77750def861ed2a7f626d2647e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdba79f6ada311c0f9b05db7eb3c908650672b76c5cdc8aa288850d9e89e4c04d7f328ac85d3ccd50c152f27d4e6b059d8f95889c7b4df37163ee7d31a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe11bb4426f6ee56dab26b61940c57f2205b6d7e6117f3425257283233149b7c15f8186106fc49be9f87b3f3e2fe40f5684c7654104771a6ebfa16b8d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb22867325d2c3186424457020ae69c0b61d1b75927a97d4f9c28256329ae60c0acd02a48ec73b8810c2e4934ba855e28a7dbb58b54fd710e920ac73f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97f6baf90c3bc0d01c95725ee093b591b2e9ddee3ea80800bdc05b59c5be3111f29404b10c909ccc1ae3dbcd14617c6da8c546468d054387f0bbb6d9f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha262ecb58c9c86df2fc79b4183606d5fa83289e6a38c1270fa8fa176008eaa81b9893641ea160d4b77502a6363552169ced0007861c8c8c62ee65d6da;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11d2fdba34f18ddb97cc43adb5618c3bce1c7f2f49e76511d15773f9cd9d16e9ecc873e45e173a8a32a9f2b21d50d54fc022ccb012161b09cc8864cc9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15d9ef4e84502ab4496389f039d95c2a055faec8680f681c0297dd5ca1326031387f25f5a2d338ac78e3a2ed59b7ac08b0fc6fabdf282db1ed34c348f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ca44a0ad3f39891d31ab4cc55d1b06640744b09a981b0eff837920474e3ff0df9a67ac4dd998f4e971742a9c2b60819815efffaa2803c23d94f1ebc0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h819e4e820ba91878f5a0cb5f1df7c40e9d1dcbeb3eaa26a6dad6b11870d460f5ab5ff05b1c1d2e6ec4d802bdb7e232fcce807037458c2c2615bde244f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f2636df0495307a2d2a9fc8a2b165b49490b3087fcb06722fe0fa30ef0f6b42bb6f2d0aea802ce493ee9a8a7abfa560e98fa3430026b3505fa251423;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bb9e8c687b3881cae282813e089bd7ff063bd72e85196e822d5bad8b0d302b68e077870ae2f4464c3c13c9eca7a5c7026f80c6fb050ebbfe6a9a4cb9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b61123bd21d89719ccc6bb47875d81b5b2b06a78cfbc3ada17d423ad12818211f70434ae5d725b25019df8c43b4b8a097db065a6fc0fada94ceda30c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h844ddae6123a1931d1061ade11d1f88407b0432eba57aadb2bbfed48f0410372176793706563b93e50ebcb56a7a7b370ddce2315ffe0c8cfe205b4b61;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h649ada4b4e3c5706a65af8bfa56f973eec106e7b37dd54a09acffee036fb81dce29376724e8089bc5ed234816988f954d7ee1948422b7121a61885cb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h795adbd32d8f9e8738b4aaac2577bc259f908b0a898cdc177ebd678365e7de5d18c1357195fc14c0b1c1f5645f4bb228694f61e88d86a2926afbd37c8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9fbf852e180b366c8998782154497dfb17a5243b792b0e2f72210442cd14e6c87b30f0678f415988abd389ed7766718cee678088143ca6fac057c583;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h961118c5ab22ba4a8cacb8b0455431f70ee48df346ad0bac6fc67261169b91f7b700a722eb91ddbc95ef5a7255391f443aa518a1c68bf611315c18d46;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64065bbe63b87a88cda5e82702831b7239d9a317b8d568f513cb1600f629e84833df936ea13850c444e61157c2c72614031da49cf9720420f315d2df4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h885ad4bbf78b6e525651be30e2b055f6f12f416accfdc0e9a53f907d850555b5e089c95e9dd3c6dc86ec46a32f11e39d967069f5456a042bd236772dd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde4b1cb74c44e699acb34df0483f8ad0a8ca0be6691c0e13c0f4ab64686f462af8e5976b4c94f5cfae405d1eba287533c8fe481c105902fc638c0bf3a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb981efc838b5748ecf3094d18e29284c44be319274fd95d9d056619ac991ee0572c6fa7cfeb9dbb8ba653812bf9538acd1da7f4772eefc7aa2c5b2d7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb9a0b731df96d3765bd9616a8b5660f12c62ceb18b5a46e21c05a9f2374ee15978e971ae648b24383e2f8b2ec6e1122066a97a5d8bf9f0d4b0427022;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fef8b82e6abd0ec70d4d2cf6fca9a1248123601a8ed47724185048a75cbd909632a827e427cae1170a3dc2d98fe2ffff4cede3387d96afe93014fd7b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf99ba2e4951a8ac0eba91f8f57ad4022c56beac2cc6b506a2e57ee9b64bcf60eb120cfdbd89966dc3bdf5fd2ed5e790364119d2f67ab76b8cf9056569;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5ebbc7fd4d5018a55bf3dd8fc0694d6d198c42add386b6d74418997ff66eff71d1f5515bf7f5ddad84696c15cc268c85a96b5b220b3ec82f014b96c5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h393309644c3f74b7a0858fc5daaea18e14b01a9a121ae418879c5776cc7e09b396468816fa9315ac5643253284968e533fcf5844259e8d7b1bfb9573;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a39ee6176fd7dbeb50cf3ad19bd5095b1c1d89b686600e931f7db65c61ccadcd49d0fb8cbfee388d96c8cfe26fa25449e1cc0d9a98eb5597e25b557d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6613e85fe40a80090e748387f39ded2b7a6425653562a26f220d034d598c49a30b26599f4715f94fc91bf44ab4906fa4aa03715b3dc71d08b3df8fd38;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha49504157efd0607027b1656ba9ae3a1669de7c8febed341b94a75fcefd948ce121597da5b2dfca88b8663047b2ceb89bd92112d725c179019b380b03;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7651d9d811a81de8bb0a6d8caf233b43e0222045621cff0b0191cdda5c1ceb8289421a7752c6b1fa7f8230a36aa56f468efd4a7d0b0e5691b85c981c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3016a85fad3b67bdc303237590a0a4d5ce7afbdebed4c80cdd33cc9257bfc3d3ab79a4acb0d943bd046d2b690b0edb18b9d86fa525d15cd5be8c7b497;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h890505ddfc8e8fc54bf8661289ebe2878cd7e215df2b50c747b294ced6989a2361515bce1d060a791bb518e70e181da9b2a0cf45b05810bad5a7f45bb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4dfb7d87713befe15945e1beac68ddf3f6255953dab338c7197407f5f07c372a2c8e6b7d393e8ed4c2ac10032c1736c1ca6dbb87343ea33b0c99a0edb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3e306883e3aabf4588ea1a6d74d361dd7d3fdc0416bbcf36e097c765073b85e2dcdee2d2c52c46f209ef14d1ca2738ee43e6553c874abfb8f765bf59;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3deba621d200b9cd9ef062dff656e77e2139795ace0b01bd0fbe9ab2027e63eb57092ed671505f13c042ce768b6132c3f0047de3d024c539fdbb236e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6a664fcd33cfc7a287a7c0f22f31b43c3ced0a703f4cd67d37f080b17592e5de4008fc7cb1d55b0f7ebd148322af5451955442c3d568afbdb0b08ba9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda461d3e9309a590506accfdf5d1c10ba470747764ce9fc1095d126a929abf93ad43166cceb2d7d60e24f4c276b39bb6b299b1b61b4d31227b1689652;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc88946ead92557f71b927f9c0b904d4cc9576adbc73182e5c930f7c5e1a0410b3a008176ee908c92838a2b7d67f31baefe69b2d398e2a88bf1dedde5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fe0f139f4ef83dd3aa9bfba921a6bdaba9114a3536d7302bec14084d6229c99b753c004dc7c7f0ee805211f07b64de6aae6bbd328e9620042fa5c5cf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he402af27fb801cbbed60b65b47e6fa09907f71737f44e0a44040844744a5c1b70b4c4e6248532e2c06cb22e15f98631b57da9a6a63f0bbe30c83c85be;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4c567d1d94b794b5392d61f8a80a702d481fbdeb2b4b99404d24db192da709d9289cc1e2807b4e5294b0914c7731b494f868b052e71fbfe8056be228;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2858d84b9cc296c1d4767a74b6f515439964fc0f168098f6c43031bf08a7d2e5748c6ea61d4a70a74f28232d22b80a2e6e277ffe021d06cd57ad28895;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba75655e3f646ae8b751da4fb50fcae0d15d18b8c072fec66d4cf02838f70174bf4e8de77d989ac2833b68293960774c27517f40070e4d59ae2f02a91;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h407212360812a70aa7bab778a33407103b07e13fadc4ad2033f2f6cdd3581df914498d85e662da27318c92ffda97105704feedd4427663dbb48b2aa34;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e3534ebda0eea894c54bf866cba16ee54e8a3f6a41d6c8b0926d7882835ef82eb6623e6c41aa5597709661f41daa8b0324df5ca89f299ef5e1cbd92;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36bad9ee21e212cd336c23a07dd0e2b9000d7a90a79e6c47ef427409925f4c3066314029bab34bb3a6bcaca493927b8f1717ad17b1b13a317a5aa3781;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha65d8a0b8d73f50da65b2baacf49f4d20114832db8dad655f6f2e34ccbd6df85bd6662efb2a3131d9db996e4d9266c0b6d77387b48ef4c5e6916ddd32;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1fd15b0db8adfdecebf437da9bf0b095162bed3e7824e1002204ea7b87bda51e276e216d9b3b4df9f71113ef78ff273c7801f2b964ee2119c45ced23b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8376d667f31f4a855de7a91ebad497408a69a4f5e049f206abae759f5796a96513647c939a9cc4ca9529e195705afdc9d56b0f186b9a089eb894b4083;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4e259cfe8d0f45d524f9ed94bc22fc9b45dfcd9be9013c6808045f6cd9c30e765eddd9bf7ae0faedf3f249b076b59cd02e8716a50116b6d0736fe52b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f6f329be5c32ccbd623078573bf717b00ee471a5f05f72f7037f46e70f884bd73b9f87f3b613c5a370b27989b3ed3411b4bf40acaed48425920c40fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha968a1590e9b56d2c72b323732dc88e2c637fe2a5edd293adcded56d3b1550fb9dd6fa4707b1850cafefcd913c8363fdb94e9456b8bc1fcb238c25842;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d292396a79883859a59f7b04264574566daeb3ea4a4d9fa4ed91ced22fa5117205e23bd2efcaa643219670ecd75549e994545e56e89c799f467fb6d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e573b00aca312a0989f154ceeaf5fc1924a84aeb67643add23b9faabf350f84ab88aff6f2b60b64895452326b93f70012d850ea2172e88aecfc8c965;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h169e6b63b64fde36ecb4e550ff6969134d8f649f1cf4c700cc9fbc130c4f6a47348f4c39b091943415dd53abdbeb1c6f9519e4db63b15d8d524fba940;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbcd7e42ee75461de92684300ead93e74079d76d67b5bab15f9a14d93ee82e616f843f7ab14b1ba06cea533b0c20f45f4f4fb604c8516a6088f5a1a55;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78a345ad2ce35c49cc0f5af467df633529a0e3fcf72500761653d9de5184cfc0273aadfb75fc858c8a8f459d942b5bf2a14bc2dbe574fea4ba0805269;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1aeacb5780e86c47770c08b0a0f6d01ee7a9e6d011b09e8e0f765ce6cf3160ed032182857363fbace9742edee76ce24a26c5410bd5b3900b861203d47;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he33ddc408bac93d63ffeeb91d3f23c57fe820c56ff660aa8c4b984529fb9fe724ee6d27f6b37398f8fd1d48ab8efc46e6f06d8e58158bdcdc68d82d50;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h457631008ee0bc0a8cb088c70266ecce65b63e5fd80fb0ad681419531b0aa5b1ba0bd79a93b65277bee3d0c25c26f96e9457bc0792acdbf0c1cf2d5e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hccd6f6b5292abbb11194bb49310139b0990cffc8e1018fcc0fc438a40bc43abd9da72241c1ca2db9a47ca6389196df712fd620b18af1580eeaf0d22cb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h265102bc5dd89fe09202454b381f45900ad7baa4a0a3d2f1ee1a3c73b19b1d256342d8f0eedcb7e6103c11f74ccd0e4767ca4e19bf324d96ffc7056ca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25c512b3327087740d2ffbf2a56be69643072a88bf197557b8066ba3d7d7a68fc727ed73c3a72c5104772aa35c78040ab418f0972dc1b10dcadc51a9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he727c1064afeb6d986ff4491aa48ab2d85867e5c8d7bcca138495fb0f5ebda1ec141d0e3baeb7099da1b68956f7fa0fb4eed531fa006abe1eca670609;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69f666007904ab65b56a0325cd4c8763c16883f9b5c8c4a585990cb0570b9a7e58d876caa3bc9b9d37dba4601b9a81aaa51406716ee055ac1c104b71e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83219537b486280e6a96a09bca9ea8f7bd6110c84b3d81ae9dc58713acada65c8d57f5d753cb14cc1f368c8ec3eca6342ceda6ee2d7dcc27e40a6b1a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf64eba5d27ec6854fe917ee410c68a86fc409220d6c5795b198f5b96fbc2a7b48e2cb51997d3f25a3a607f9766facd532f6ebcc629344ad9eca670e63;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2051af6b215926b5912f3804b69c8905e4bad1bc14dd25e2e1c33ef45621ea4d5e92e0dd09dbffc34f6a01eb4dad5c0ef47f430e1b5b9864f5d687c6d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h834cf440323626956b506499cba87dc7b87d7ff4e7f5e3a02038aaf3816101db4770278e935e5fd854c1f2100fed37ebf2d8fbc887b9c02488ccf07dd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h466656e6e16d5e35c4e8caf97314598fe372ab96223b3173c5df4f4c5cb2f31c9462920f8706c64f8a18249fba09044f5337b5a27b83f2dcfa3bd2173;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd3f04af50cd5f4a59bfc429e8af0de30b9d5850e41585253d165c06483eaa1ae89174cced8be179e7cfb2abdb473645ec6594f21c48a08278ab2bf59;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9de091dc37d870e139c8191cfff36da03442950fefeff758af57879a3b323a387d0c706d3f749ca96af4cb5b90a428038c549f4cee4dbdfac02e409e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ed2ed0e48de696b880bd0bb5417eec65ef55117bb7eb733e716e6780c4e5c654197140768046434ac99596f23c85e2cf7be3bdf57ce03f738565e806;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b94581e087091d9bc93e40d8f11779fac76c81fb41de15eed492a82aedeb7a874689b715da40b059b21bc89b389908237141f5e961c622d047dfbbb5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e063396dc67944467431e15c51a21963c686bf1d7eb8f2a94c713739fb4f46150c1e518f720d620975faf7e49c0d5a0e4503272406562c6a9814fecc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6578751b98596cc779b58b794fec0e4eda533bae4b41c02ee69a2e3330cd0cd280d3c842dcc3aa91ff2f3573211573ce3b06d8c5ceb5770b7db705c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30b75b7bfc63305d66dcdeedc3d351a4e3afda3eed48c2db3e151cf7b975a4dc559000a0b338b7e6be76174c4c9b589be6dceaefd4742a60b08ef0ad9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8935035e3f2277ec9d0d34bb861268828b2b530518339816e0e340353151ac62d3adee0f738db44c5f168168210442b914ea546aa7093d44760d63bed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d2670a0158ea9725b9417e867c2bb1982250a8d7a583168dfcd3ab812fc3517f0f00e977afeca2a9b86c6e3bdc6a7c044da7ec9f23ec252b609121ae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc232bc9c62b15098e90d7b46f896c57494df29b6311ac8ae39cd496e990dc6c638d8b0893206829d6fcdea37865eed7c7d87eac15bb94882d2b67b9e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2728d502b2d516e4459c99c07d7109e1d356ed654fb8ed1eacc067b0a1170dcc0febf638ce1fb6e1cd6d91c80c52b1a0382901c42ea72e8b015f1521c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hffe182c15ace5a51eeaac291a9676931ba9f28249dbb205b8465a657d77bf9304352d83fe4172d9febb979aaf272da50e227b9baeb0d877e9b554fb0f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc5bc08fd76317daea5985118e27e11d81ea11706e95bef9e014461a473c85dd6c169c5e7628c156397804ad5179c7f6a525d5d1843f89a571233377b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9676449dc5f55ce3dd5c1cbda47f34ba7ae35c0bb6a8624dca7ca1fdfcc228e5b36ecb708bc08ad22bed7e27eec8e814ec60ce785238607e32c5e6a98;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92f843c0a8efbb6e077e3a083536577ab63505cf52a8b1dfbcb5da413fd2213ecb9d52963141c2554bd3f949f416055086a1d6ee1897ae40263c69ac1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67f8b6d0d186c949052c1abceede8cc8de9c6589093e2309a2ad5349b3a0a711dcac2b60f9c6fa1130f59ef0c6010a4a44c6acf6c13bdb740415c4191;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6390a0d348d445420a5da83e60d5f47135f9eb7fd2b505c9a06ee2baaebb7348f748ddf2c6c1ffaa33ef1052cc5ee3d124a247c03e7738bf8030abd1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7417c2f8777172821374a3c3ab9141d6864dba072c8e36757d0f09f3d133466af0afd5bbf0e3caf299ab506f86d07b155daa0cf27cd45862ff877be11;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91b6301ed8316040cbae95d05dbf52685dc738e6ad204c63a5039262053a52c7427927edfeda06774053415b6b09efbc3f44f9d38a496ff7948455f62;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28aab207890e5fc7d8d6b235ab2349cf36a5eb11a4c760eb354676cd1e829ea1dead941da055c136849c239c3d763205af49a0fc17c032d1d27303de7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4165d08e2024927dc2427fd0c6a02e1c68fd60b8704ba1e476bd4a9e220e40c6766ae799f767c275778a8e1504e964e46b84672dddd3fd5d1148ba108;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc70866a1561b92e1d20b7917612671523f5d978b54d94a8f5b331e20e45f89800f4d38a57d757eaed177202732bfd99bcc3406392766cf8b17d2ec617;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52e1d9c6d4c1d98b8080ec98857fdda9c534319d2488cff0264a6d40a8018a5f1624326c63915acefb55adb943edb89fb721354ffefc4bcdca1d39dcf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31a5b629333037fade032533e162b23a4fd02de6b367f4e9cbde1466fca6d8df1e41b63ad50bc2005668363610e1339b7a50ecb389b5ab6f305e71720;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59325baaacf35c1bb20bd04187496110f6652142f61b944efd7652f9abc15434e2dc8c00ee133de5bcdbfc36b3fb10d6a25ed371ace6600a89e981bb8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd8127968163eeb8170d16022e2196cf614f002a9f4453d8b95d0512018f580910c6a117e56958b6bf4eb526299e28885655034bd4ad0a3eec87bda59;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d1e752972f0e86c6a9e304e315e68806d5bcd01b43e7d6cd9a849ee3f50260938bb4d0bf2f300c9e4d3d52a3b12a408e39f42f69092325613cccf3f1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6f07b0a40f6b9999d254a5e719bedfc74cfd9f202e86b3f7d28f1934c9b90262f944491e2638136a4bf70297e3340494ba54a97dd95207f928e95f36;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45234fe60474b46005128c187ebe843aa8aecc3dac8823c25c022e4198f8ebc25aab3643786bd94680291a0f5691eebb2ef464962ba2e9e92460a2f62;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8eebc1c54fa897ec6d7500f1f14e531e1800930550f8a939bbc5acf2d63b2924a26903a3f0253f15a4fa6298d0fbd01be1762a9372a1a8597f228707f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cdd73a22773088a24b5ec7e9cd31fa7fcb1309a18708ffb4d34090abb2073a82959b1ee9f7699645904de060b8bd696a21a3a9ae1ae060909a487d95;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd71b8a51f57a9c073de55634b9d48dacb16043de68355051204e1930777b900dd284065588b7a981f17ee0b8bcdc8dceec124504a73d0202361a96673;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8f050af9fb4a578f95d8206f34e9570656f26e02b54021f2da753df16d1a02eaa54869016bed143f442957ff3053526b3915dcfc9a7ad777fddb3240;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39aebb5f5605ead70e4b9fe6e104be4961077a8b70bdd71c3f535b90dd824dd5d9d22f0f464a616942c9ffe57766c26ba7116086b43bc48af0006e8cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9087fb5e6285b8759c57bd3994c31a5104a63c21fc0685b424ec90ec3ee574dfc43b5e357584293250265b44956b27419e4364f6018d36afac901599;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h254e33d50887c7cc633af313b5b429928c208917d79304715b3e26b19eb8be7d47cff74fdab80b9bd625682a6d7bbd05bbb85e2d3a52edffdb53ed1c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f612415a2524df224d279ccc22142a96f88a634ede1d84b65bf483870f11b942d25aec88e3aef3212921317bb50967c38ecded3ee125fd2e0de7c2e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3eb89a047fd1e91b5bf2f89098047a0de69be3556615ea66ecbe31041a073f2f1d5771ebdb20e6cecf15fcc9502f83c684a1a9ae0c5b5fd310ff2c8e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf26314f3068b1c07c82437c54063540a74c0b38993dd656ad8130db338d986fa8094f1b017e78d03a9512e54e3f6481030b9a1d22ba66b8985c0c1b5b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he241c47e29acac9e275b64fb61d983efffd5a7dc6faef779394fff30f2a497b2578ae87e6697a707f43d03416b75f84a09e3977000561bc98f8ea4df9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d18e04d0ce8373ef3a7b5592b94dbf739eb4a040e6fa05d7cb82ef06f34c5f5f60c78a88adbb9e4054712d88ed6bb2171934428f4f2834ebc7a57bc5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6709d5fd5c5c56f2aa88352b119ab64198eb274a7f42b9443571eb1d6175705f4f381cc47e5c2d3d8cb9d22ac6bcc2f0badc2fc6391eeca70b68943d4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha451603970d02b52bd300e5de80e021c20b219fa9628100f15bd1e236b2a4ade42b98af5bd8dd6fcbfa57ae9faf995ed895573bfc4a6df7e1f7240344;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d23b2d6f382cd08c85ab3762c9f1559320afe3ada3dccbf498f070e31ebd454a71eca57ad519b4bd97ae7dc1f2739ea6e9ba617f2847dc2bcc78af24;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3aa5fee8887de1745851a3332a315b8fd23909c2d25a880a489eca033044891e09ff6945a22a8062daf8ec348c4e0adeb3cb0badbf7d309f32d147473;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34a03836ea7f94ba178efec9c607b7f336d401d369504e2630c2ba23ba38f798f2d4dc1aad916b503fe21c9ee1a7810e7fd72d4fad125aab9224c966d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9da2df244cbd9821e03e0ee7a0e38fce62707b7e7ab544b7b77001d2ef72a06442dd982f17633d811dded3e30cd7a55a0f4ebabc0d2e9cf942f35108a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb94eded715b82ed1910f385dd3bcf6b92bc0a2bf77a1fd8a68cf9557464a20f2186198d78b329b1bed9c9ec0b352d26c1837403195105a53b72c510a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97b7ec9d57893d4e1da12ca32573958d063bb116f42e83f00244e6df50adaefe6fe3807cd4934bb6a6b3ef2e97396810e9620db939e89239a324c9c11;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c7dd75947f07cee942a1770ef426f65cc78e39628a79c2f7dbac305f19a304acbb6347a08a28fe8704edfaef7217bf21464dc71b7082f36fc2e19ef3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8bfd74a1cbe310bc47f5c5e8b3e67f9ef479e42bed5f155cb9720ae8c2fda8243e3c677e35cbef9a86d62f4ae50e79443f8f524cc986825fd4a903bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9941cb6dec55a2a8d764b232cec40fa53b1af8b986e1c9c82354e15b8ec2a6eeffa32529acffde7ddcdb4e0363334dc2526b18ebe84bb00fd4be357ed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87fca7ce4fa68563a2dfdeb5d3798682a1c60cc1555f3264293a126921f8cb2c4a0cdd3a9bafde72540c5fd9a355722a654ee8d55a745e602196c9df;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd51c8db839cbd42fe54ce8352d666a0cf0bd5e74bc6c477d3f8f10ebde5a4f9c9746264e612a8c81164375388b1bb6fa05d74f72663ceef697a4f66f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc12f61bfd74ee5780e4b56bef2ddfff87d1cb9aefab0f2ce3477bae5daaa6cc9caa7895204c7cafd2521b97635108ba9f198fe3ba1e15db39ed3686f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca2e9e568e63aa787742b28053bfa743a10791cd3dcfcbf0b96bbcf2121dde73ba865fd1483c4cfa3cc292884dc78ee8a5f8f4bd491a4e8f0f87dc950;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h747460557362cbede002af04028b48cb86108b5c2285d4b3ea4afb08100529ed4c56456ad73627ce8744a88e05d0eed82e0ebc2d6e4345cda6dff3c48;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6b60a09e64cdaf8cae88a2478826f7ed0a9da4f6f74b6ad34e816786e47c88baea48df5f7198b15757e4fca6c37133040e636b10948e66fe405dd845;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h472feac019a3271f9d4b04f5d2bdeec6b6923e8d615d1984e1a1a56cb57c819a5a629bc31050d5ab68786ead95b15847d6c799fe574fcfc2291a2349;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h318aeed517f886296783f4c73e5cd9601d6f019cdcfe274df1ee2f8a535863ea30f21f617822351b386fce49bbd20d8bb4a50424845b32de87ffcaf19;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76a057f5e68342af6b8cbc65a2ca5111e1eeb1e4d36d2564ea8feea691edea9f7a14bf3a0e6cbf5c586b683c3ff5cedf33f0976ab502916f00b8ded8d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45aaa19505893fcb9702c170c4e909f2a4c8d7aac4d00fb1550a9bfec0f9116734ea3719001faa52f228f9dc67c5157348979e659c1a16ae6533085a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0e2153df4bee93e9f5e348b29ebc72c124ce3ed9a39f3ab30150713b9159042a3734906679e6a30105a855defdc57bc345c7b1224eaa46aa024847f5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haaa4afc548bc4dd36cdc232699f01408eb6c6decc0acf396681a9a286ea51f509d3996c8e502139e62fd02b01b18a1c0b13e45f5e5ac252e9b337b110;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf61f944ac2c44a34d9d863e762aaedff28cc8c7efad023bfa351369f355d3def05fda577e33ee6a8e44bc6342b70e42a70d9f177d38a58da840aeeae8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8df66ce66657aa4137bde5db7099fa73407ea6d065bd9ad4409f0ec66043ef6ad0b72c3ec7b06e5720842fbe8f9d9a9b8fba719c30e7ef4271231b0a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf956ebf1384e1746a9a3f2b846ab0a175b648d935e905252b05073718f0e60eeeeaf465ca960b1dfb65b69a2684a1ab819aa6cfdc278cc9412f5b5310;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h846c10c35fa2a6bc271d90c9fa7a8267bd08328c82a874a3410a2d979e26191033090631732f1906248904cd079f99a71df1bba3824ec5086a22f230;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4260bc8cfbdfbe1cdb6e0f51729aaa09891bd81b81320b25fb19b36b2ba374e050e5c4c85493bcc1bc6abd218246e66f8783c24bc5451b5d251e3bb13;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf75cc325b2fe7dfd3fe1d09545d169eac7b589b4e6982d11dd653ab570e0133cfe24abaa017120e4ef487ffc48b9f6e749475dc113ab89fcb922a1181;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed00c19a68bd32fcb1d619e2850edd674798a11c6173768b837d621fcbadc3ed6ff6eda0b29e9b05963c1efa6bcd6ef1394da2773566e0e879b9cba4f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36d6d9e57d649af82f4fd1f9226792dcffca12181c3cec547979873bd3d50fbc742a2dba5dcbd6e6873d1db9385f511300ed3d662dec3b573622252cb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he02c36520ed5c656a0f0bafdf9dbcc3d6aa4da760313b545ca944eb99f1f97a930c757ce2da98fa0e0f6198c59c36af8138983ff0954c548c34a6226d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac5808daa6ff350f151afa1b3764148a9044194896e3d23243bbfc7e7139ce5ace599d0093b48f29fa3cb54e70cf2812758681f91b6e5669e649675e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a05ad0274ead0ed60148e187db213dc2cd299db4dd8776a6ef9295d1182eac18310081f1b1fbc4d54331b4f8f7df00d09a095cfef25b098802a41e0d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7560babc42cb9fe6d63002c4ca5d58fe749c838c57f738d5a97a90686b3126e5200551d313b3f05b1339adea6cfa80d5e979f1de5c4fbafc63aa31550;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h615953dde2da4b7dc2935203ee38be68a43cb0842d5c4f9523cd50d594cc7462db49a01b7e2fc57202b8c7e21aaade61455d59956530df4a6c8adf964;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1b27eb805dd033139583b1b6a2336c20f98b680934f0de2c19c77486824c739049fa787183456c6ed9dcc43acd6d998a6c55cc63e9ad047c7a88ada3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7483b35c09a7a7494477ae7bc07409f706e5d29bfbc4fd63f0390926388c856c6e655cd0332712fa54d39ab559428bb6f44b5a50fc42fa9df384a0909;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb114aeb9c69e9dadd28d3fdbf0f986586d11e5a41d7379ad94c5635ecf7681290bd9aea223c452ece27a4803e8ca5334ecbb79b5622fb5d8e3d708b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20645749758fb2a67101f955a31a97803945ce01bdc8b4079545fecc9833e16b3ada050c648a08f11530828e056c565e94a0e1cc1b92f985cb8449abb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36760da22d57af473e2af79d223315062f1b965434ea8420dd284d53663755c9b676391d1d34b07659f2c766dfa999eb150808cfb8d7100e39fbd280a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81280ed351a564f44bbf96b84774d5fd2882b28c2d79a696c2eeb6725a4242ddf2e1271838df51d31704e27bf871677d6c2193b9945d6f64d2f087fc6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9e7919fee346ff207c7c6aa9e5de4ebbb6cc58ec6e7891d5fcbbd4afa84a2790493c339ea8881d48b2295bea36780f019032dd4de714636abf74b01e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he23f794f3733b3137672bf12ea507f97cf1f8cdbf490e063bd817013d25443cb56b108a0e0183248674de615ca415aac16bc6c304231215af6eeb441b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h432e7c021cacd2688e0805a0f0f5301b28aa9610e7914be46083e3874767e32db85d02b10aae8e17857bc4f420753ebe5c37970384426c9f9a547804b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h286c351029c26acd845e21d954af26c6718ece79aa010acb90411a686fc466582acd08206ebf4e887771730f69e2f82220ace8f4437a2225bd49f7636;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41b71eff3303d672a00021075f879208d767b32a9fda214ba371dce9bd63b8b0f584ffb67524f65c77f817ca50a7c8f3581486a84fbab77b9c5fa7e30;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62d1f7b4ee7cb81633b1f2420f62fb64c39b613e8f67eec027dd39b081dccfbb2728e8e6f57f3704bc66cd6140e0c904e98c249b84c7f4510ab773211;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h536d7aacd187ef99be5d98d2bc92549704e55cef0c04a7f11d79cc9778ac7b6dcf4060fee5e09e82b56056fb6d476d1bc6968c87fe235c05b46d308f0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73047a75a22104dd62516e8ad3758c9ba9acccc93d48fe579bb86ef5107ecfa1470be3310ba67488ab1c47ff049dce67e274df3663a8747833771d757;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h177edc9e8d160a87c486b72f82dc7b69bd111f7a3b4ef2034a6678b33c759c1f59f7672f67302c79c40761d082d4f0a653a857ce8de79d89016721809;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha42119c67c278da17e221b8ef9216438b165fc2288046493901044dac216e8dd9a800aa592872479908741ab0ee15db24a57c5bc2b2f4b2cb8dafb86b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16a3c197fbb4d6707d0093cc38bfd23b685966109b590b9d37d93e7904e7375b330a13fc0354b11d6a3b130b836546f6f74b84540ad96319b8475ae15;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48c368dcd156faf7d37e3d5d479332df3a176869068841daa557d952841ff0960ca9dcec4d651a0937b84ab27684f8a4750b165129df1e8c8975bf265;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefee33e412830f006d2f7659df1f8086701b945a29ac8524eec06277ea7083a0ae5a56a26876361bb7b8038fc799d6ca5cd3de7ef3502740e03db775b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h437de2bb70032bad72acf908249e5a1fbec45700f5b9c9a8a7174d92583c1c92bcc9dbbe4f1dc007419bc4d7ed574b4087fa8acaddfad41d635b1cd9d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2db49908cfad1e6cfcbc879a400680c186009dc1a2a03c2bbb8c39ba56017031afefc122aa2dc5a7b2e78348e875d2622887a97761ac0d4736d478a1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h282a8b85f30eb2ce88c518608958f340964c163cd8238725b35a3ba23a18f371950ab2b5e837cf602ec8a601539b99e277b2b25f2097cee70eaa925d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7973fa3b10b0d1f78ec8d498bdc7e6c6a87569ffc6a435c786770b5bf9e69a4fb138f256b31d72160eb0eee23afea4206fd639b835c7e8fc2e4850e24;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37a8aa0730b625fc9fe84a2c08cd7d2741f80e418ba76d8a33066718ee5a614367028181aed24522ad2412f3c12151f97dfdc50b7c8883325973ac611;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda5380f493dbe45611f1970e599428d53bd51b70b50325d0b3d7e949d30060a48dbb7441b9c734ae1880063927a5868ba6234af036f6ff8644f85b0e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ff9842a616211c623eaef294a8da3c8894491b400ad3ca872a62b84e6145fd4d20ab0a6365fbf5a75b63129a161664fdbc6a22f3a466b8d08d168fd4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h630f2f70a5ba214f9a26f426d064c7f869863526dd842edbb14cfc08dfdb3c61a3c6e8d40e37584e240b0dbdf6726e338bc0bf8d136d4979ad9d83708;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4596a2dbd5a226500695dba4cc93abbca785c40b2cfe54a68c341036476060572c6abfff05323b453d453d0518d7fa2e05016dd02022b91354c3bd54e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h879d2098f4457b38ef07fe109cefb1508ed3d6b973d3d519598f789286a9c6d720ca9bcea2168df83c7210293804f4043e3af4980f06b7fc60b16cf17;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd41214849fa30aa9c0e01bf61aea2ffa451cfee177bdc0bb20d604b46b6c2b28def4e8088c9148d133c83372eaabe768a8020840b6151a876d27ff3b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0e541813252bc45c2a4de3271bb5d843f4a9bf96c8df9b348e4968904046ee3069256e891157df8c7259b98655f4b741696e740e40f69b8d4319a1ec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa8a6693dcc37b651c669a6dd8fe1c19ec25ce5f8a8a4303f19258a9ac6d66d836ee017e472b48a3b5eeb25a07d58732d3445adc88e669ab3551167fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdab84beeb45537fdded7368fb9e39c08f8fd840c05d8aac394eb514ff8ff2ce68a5ca0db85bfd6e0b4f6ecf3c6e58723d499bdcdc2682bcb15cce5c99;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf22924b28061af0de2f89bd5fd9cbdfeedff2964c57fc4d88fe00ac5d4486b077717100c96c31a3df223cb1092b15449cdce5cd2aefa7216db08b67e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc928c95690dd1b18607cbfb6038fb59a9d97685d5401d796bf947050dd43d1740a93c5cfa056671837b7cbf3fc4a68c41341b98ab6e6c71b6b4e42b4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52517f7c608e9f42e54f3680e0af870638de0cb6f9ef9d0d25ba6f1e9ad150f7ae58f220bc3e9cd4027aae25eae7ba1bd790c436b0b4b0bd93070d2c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49d8e6418bbbc19576f69999303bd4aec69e8b9b0dd99ce80e54aad8e36e2c3182df0572ad48382ba2d3ae3d13f123c3cb1be2083ca67fc619f4a0bc9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0106bd39f35e3733081f5d873ea642dae71512904192b4feaa01a0a448c66677b29d8d7130f68e44dbea4c7502fcb33541929d4af5d694cc2bf48c3b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d6b27795146bf2fb3b8597d3ce35bad6b458570b76c4f19e63bb3c870b4032ce5e78d2f7f4f498a616ae304c7868199a2c07fbf65ff29614a7ec4868;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h874b597f2905157230d6cca9718def1a707c8dcd5b4560e8e6bbeb091f781ddc5415e52b689c7ef3ff460c90c894e59f1577786e62e9a851867d73bea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9186293a26d1cfc02c10b2ff0c92f77de2ffd365e0195849154dc51e98cd881fde9c655ae7ad6c7fc43be0e995f4c1c22d7a22925072a460b7f7d101d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb65e166bddbc4119805148f908d6d3c54cdebfe8b1d4efa82eb855c28766b1663f77e691c11c6b670b93479e83f4cfb92cf906ce3f414225ac57a030;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h873aba2f2680bf36e8d450364944b4edc6476cb4d543d58267ce7ece9ceb51fbc0929ec59e3153db86e08b3360ede8cc6406a2ea54754e7bef399667e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedb1b1f414f1acb0e815a5afce2404e8eed7ecf679599e84d501e594a73172ca59842b04fa5be9b8027f8f7636fb3af3ee2f1dbe315443572c37f6109;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde3b53a14381d8bdc762cd3c71c5bd10e3312b931287f8abeb12bcfb50b94a83a24375757aca4be1b0e5fa9f185f171c8b8a29d0f72e74314712c5764;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ed70f16e492f1b7b914277173f30168f29c1daa3097b2d76455e31e2f97881b91c199a5c3b5522e0950461d10ab213a8783c74c6e425258416473f9d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b18fc0cf5db9e0d2cd8b9a3440538332349005bbe462d4e0c44fb7b8e3e595a1cac0102dfbd146bd909bd52b71f79561112e5070f5108659de8866dd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d52aac7332c46fa2b8cdc4926f2097228ca2e39edc7cecc1f3fc9693eaee558b49555cb57d9cde5c62b9df8904c10c078db60afa006435ef24d7cb9c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0eb9d16c89058f7bc9c86edc5b620766dc22d988409db778f8b9bea3ce1d0266bbd19d9d184628b1a660b89ad9495d9d0a62525facf33b964023ca7f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdae43c7a186822b6a5cbb2766d45e85533b5d8a2d49df47781d0407627e58ac5c79d7db73f3b6431e47cbb3f31fb0f56ee4b2c568e0a3d4ebeb6f8e6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h969a49cf423324ad69e717d603c98bcd76c4ef0c259ee9db473e24ddcdc851105f71e7258403366d23256e3bbe3e41e35a35067f1cb733333084de0a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe2550a2e6826f95fa611a4971446263a945773995ba596c3fa0ebc925b42cb38a28d46e053f2db11a65cc02e1f72bbb09e2630c41250efd5594d73db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf60eb6bd013e49988fda979a25caaf6a2316ca5ee21b4058c9697f6e8f6b65b7d7d9c83b6841d113d82621a5d8a58f63262f6e426cf77d574a984d8ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc608e0829033b0877a05e21ca31ed45bdc4110ed3fa10f9e723a8b6a2ce5853750e2bdd59b3880865e3a7ef04659663e505f6d57787233fe3df6392cf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ccdc151c6c9478e54e7c2cd02364d4175e6dcad183f814828961711eb52dba6c97e7e37bd90521d668e00d0ca6ba80b57fa0c22adbace0fdd042d8e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa840277ccb32c9cba694bc6f4938abd4db2cad757a765095d3929814e08cc8d6abfa7701beaebce6181d3c3816528ed0fbfd4be7fc348138c7f9e527;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b042cdaf9e65d8078fcefc1c50d55f748fe17a1f056865ec6527d37e9983edea82d3a62a9371246eef35de96a13416ce8f3c1f203604051d5e60a23e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6324e33c24ad31489af0bfe933810ea2b7fb43a4cfd87e97648d354beadce9e803ac305582faf16ac24949c45870b5780f6c99d3c58e669bf0b4ed821;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0064f019b479ccd6277335a2ce2ea53780c765ba4e525d14c49b913f17c2f49857280a27fb5d65fc21f20878ef573646278daca7582350d27a32dd4d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14cdfcfa58416ab65859bc0beb5bb3e1071bf6874a98bb71eefe0fe98947f118d1e77edcbbffe5e532f28a538237653f754afb2c2660f85672c2f838a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h552824b9377512654003e5e0d121215334f6978ddaae0481c4856cb024cc0e901ee9b3cbd25d0c0de5c903d5a6779a99703bd7021841ff9fae10b0d8b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd44394622f7d5a60155790732f74a51bee66622aa2f6ef57144080c1acf995e3f6e5910e22a21017fb822d08a0e1aad51dd2df09d99600eef73150889;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c79780520c7a4f268101eb862ab314451d0cced188e000301390c637f30961f1d8f4464cac34c4e763cc09667c7f16ec3a90ce543f25679328515c01;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56dc960267d2c54337ad42176e7c40f738c9dcbeb8b10c0de83a03cafc5092ba40e55cc3514c8ee3b039d18e8f2fd67547d2a17a4d08ad8e7d86408ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1e33919be06492425302357d6254826e4ee02dba187770c20df498417ffe3defb2c96797f140c4b050ebeda44d0046333d5d75af34b22f309bedc83e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5684f515b1e0c6adbae88c317cb00732e756f176b40aed5c2f0e8bf3e1424399b1597dfe1df30fe509fc9a11817ed343fdf102a544bbfc1fb9bb96f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1cb62f7cfae2945225f4c9968318219ecbefe832b449675233eb3db32f80f9ff2fcedf3553870ccbc7f7f9ffbab1f48187b339ed024bb600899a3374;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2883593aae71553aafe5720b2b105f512bc49d0bd7bf3c5a76aa60a8aab7e51bba31c712c6f2261387e2c4733882a7b0f8ef7c5e4752dc8d8309091b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h742493c5543cf1176248550dfc3cf7afc9f5d9cf41a96a639d49cb06e8b2da6d9b06428f903ffa9d90bdc1700ade6f7268728197f42bcd9fffe22c335;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf52fd3b10069fcc878cf608db6a450214152f4dee1159571415fee1c63a559ad0b632c09e9922e447de379c3dec453399b508227111b327e3c1370f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a066f2d494ecdcb0b1c8355f41b6fa3447d7b42d29761e6268b74ed88661407f55d33476d3f2e883667794f441ed2160bd1b8d8dcf49511328571dff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64cd80d160f317d1a1b9154107d8a26178f0d78866e4bdaf15efa27cb96c76c2e66bc8f617a59e38f67d0055e77ddcbae371d7b82f2d4e84e2fb1903d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17ae692f0d3b4f941178111053e534d3a7eb40040534ba117d8ce8c8ea81dbdf31c19c3ae134a7ea2cdf1f37a0339845b31fa9d8f696d13fe3d8bcf0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd022c9ad90dbc5c3cb0367a1c9be8f79062217aee0ba063a66123fc030dfde0b4395d8ffaedaea34ffa10275de32413cfcc9a82e6ec10647c36a340a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h639d636a9a2929735926abe303c056276ea1eafbf76ffe609206a2b358b6bfe82c6e4fba53860e9f6278991729807a888f2bf47aeef75267d7a02a44e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h763417c013010027fa79e88b2d6d7d813deb76014eb91812144de302e6656051086b3115f51d7b99cfc22698c96b74cf3333a7b13c9486d599882d8d4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97ede521bb670dbbd538e8ffbe175d6cb2295dc73b37afde1e4844eac5087ac13747eaf41ff6ce1c965fb1ebf93da83ebb27a01e9d73b650ed07c1312;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ffebda604881bc3dc089357d45389da821726f4ec678622659ced0e9e7e555e45b7eb83569bb347757db08a657bf6901b0ce5bbebe1cd2ae1878bac3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde526b7c7b24a2403404284cb2dc1dc3a0f7cd12fdfdf21b9dfe6398f7719b1aad52bf1acd23315b8af3a5913d2b0f70d9711c9d0bfbd52a28d6cfa32;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79a65edf3a0e5b630adb242a22808c21eea88a74107379c2ab4c86a9484ef216efa8cd267f94e4d0b42cf6c9a4dc272debd9dae91485d4c22af06ebed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcaf76445d3091da455cf2c403ce30ea6b348794623084c7373731f27099da62e44bd6186d9eb96eab3140c8ec2e926c9c79bce3e01a2d7ccb20f40b32;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd36070f0cbba87c144f3cf4a4ff4779b1d6034eb3dc18b93233527b8c6bff8ee6fd2454f3b11a1a31fa85593cf5992e3980f1a34c0924bda634dbed9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb608f5fc802b687525cbd7c5b4049b50fea0b256cfc7bfa221f205f536a8f209583cbb49efb4839329c405049e0a0b29ec34488600b65564385d0c6b4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8810ec78bc40cae40ef2c326844b9e91dcd27cb5451451b551e5e29bf7e1d19227548f8866d193e86cf8e2d5f0410fe9ebbe4a1f216bd4a48f1b91358;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34870afcaf489b29a7d67e01406ce88089f7f7003de3b5c02b74f76479d5805e5ae40e38d7b7933ca20c5359518e5172377c7e38880384b469b329125;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ad3a78af397df3acda8d4069e199b289edde2794daba5edc1662c31e6419997691f8801aca86209aa2e106994b4f802f1683671c0afcb3101955bc46;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e374d3c8365818668cd8defb986be5708467fd8a9ff5a7a8feb6395a52ec248a8bd12efe921165a6800afe3b709389bfff50f0823ff84bdcabb1b8a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h969cbf2fb42493ddac2630817f5a2dcabe6b1031f1ae217c8744861eb35511da5e980592f571d4b6ca8b303bacfbc3829f7ef2139d50194482fe6d114;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6dfb54930367481915d9baae4d51984de276056c9e0866478243367d89d6219177837e1681084fb37f7c95f13e512e1a3ac12883efb76bfb9491b4053;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16b2623f421f12ea882434d91c6c166bc66d625a794a7db4ab19b3aef35cda3b38b72cfe1cb798fe374f61e096d05dd4b5d4dc7d5af4b8903d1ede522;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfed2b2d0dff2f8bdb0110906cde10c98eda0cae4c6091268716580af62141bd84cbab55560b0504863d86e98c3551292c40629f324b52b90713663759;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6448e03ef0691a9cd79be2d0cfdeb5ba0095900a088f5a8850e771eb212001e12a1f47968b47c2d2cc88c7008f23dd4f75901ff5f4843347d8b0fc9e9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h541975bd421ccb288d653ecb0382f26dd2cc18c7267af0bd9b03d761fa24c232013d4a3cc7684df649f532e01eaba2e3616cee4f375918e76bf10f90c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5fda2ac6975e9384e27272858748872a2d4afedf8ac1e94c279c366b775d23ed058d7ec9f5df7d6a5fea26a95057431dadca36678b36347140d1a331;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9bf63787ec515f17082f7101f44e3b72d5f80725b1ad9ed17b656d5ba5d126c27e60e05a57900aec8843289aa113f3d5e950db22fda689587db6b894f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h478b32d965ec1e48ef41d6a930f2ab909412475381108da9404f0d406927d55d2752fa74c05617b0f46b73dcfbd2804d80a40774c150e52d05f88ab3a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h576e2d1dc928ff435b5de78bca3d0108ae1199fe4f4b73328c949026de59fd38e5f1bbff8d9f3c434796e010c6ff724379aa0fa4401d3b5b7b2114f8f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8552b0b0d83c87886770776949a09b7b9d324f3a3996e9a4f2b35533ba59b90e7878ff8d94106f99f88be9360a76e47ccb6b16c2dcbd4d42196f58aa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19c760db145497a4ba150f4b65608f84aae52c134a8ea3c89b34bcce49f34b172c78007481e0333b420f77ea33b79dfce67f7ef9a2b944e9289c81212;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6734e87f22b90b5a12639a23c7dd479faaac78aea2d7a82a7b570eb0203f246deafe101c9333ec5daeba1bfda9710adba1276d748f76a84529f0b8506;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d03d3fbe2f1ea6f672bf6856ce6c466f29559eb5d8a074891adf3e746cd0c4438b1780601916d26c882690fc1dff560642266fd9d3de5ee5f14e16cf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83b027a34b0e63bc460aa37168bc9cef661f7b7b11f4d2bd69d834f64fcee409b1f8274aa1e7f83029e529689d1a778c264e95a8b4d34ac411286eb8c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb56b4bef7884d911326e250629f0d7ab47ea3ed7006f45c150a2473b85c22ad4588e19a18875bee7dabeb0369e00243713698dcb35627e9dad3d8865c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha912e63980e06e4b3642ef493bbc2d280a9ceb16a16bf85e82da24ea235ad37134d362c950dc76018a23f4e50d6cec5785c9cb9de68fb13ddfc9767e3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ced729d89113be68e5bb01a6e97e1ddecc49bca5ab64108e2b567f7af73afb56a4d59647af577d94effdc21f33cf701e141497a47fbbfb9387bba1a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a30b8beffdae63fc89293270eb973729f88e630410e55a70bae4a6260c17e1962ce071207a73c40f144fcb2059353aaa808543f4d71f56654f1f6e34;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf86bd769541aaaeb1b3e2f458cbd8c231856b661b034c380eccb1bf332e26c389e45155e7c1c21382a29665616b1f6668c00007bce4f50755cb35c921;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33fc9984792019ec91bcb9a4a9d486452319f187b04ea393c8a1e9dc9340c75b61c9446315e2e378f18a6e3264a3ac9737828ca27f2efd322d2ab6223;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ceeba0273185dccad5545e568a94f4e057e103ddd3a3d92337ba931f0bec318cb7529ad1ac59ee55839e70a903cd93a767d1096dfdcf9a246cc83c98;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3044be239ebbad4f8343e12bfe28f97f8b34fcf055cb11cca0d32072482ce9f288cd85dda5ba713ad091a7e5e4ebdaba493edba8b50215a48f7ff434;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8cf30f841e21a7d6be9e391983102f9856f3b7df0e08bd67634d029ef617921ea1dd2680ce7f1997406bf5b6569eaa4fad186506b6be02d037331ed23;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba810fa5dcc9ad33b1b57e28a2af63f063cdf63636e072c1df8ea2aa399d38024477ac2d9a0fbb1084dff90a81fe1ed84669d74bcc3f5783b4861f403;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ee7fd6fa4b7e424df7a737a807d723163f4e7954ad51124357ba75c996989016acac5e6a1cca70c6f858f2e969ba5ee1a47961264ab8ac0bb1904175;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0066787719b174828b5b97b47812a645f0de056d7dd819b08ff5e1b687463792ee8df2e5b854d38be8f7768669de10290537251ea981483c88ad156b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd719a3a99752538f5cb7274931a705f51453fbb807be1ceb31a2a5c9de9d78842765b8310da78b7905dda401c1febcf1322deebeaf8e7bda6489fe2c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h925d61527936af8c8fd6dcd73d3f66540fdb74588c4a83533c72bcc5f4c54502bb9ad39aef843be0fb0aedbbfeeaf1b2e9edaa35e6f27d9fc7d12e1c0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heab058e9a59ee21efea47d17bc2331589d7e3f505504b36a0f4fd9ab7a83a81f2fef9c48062be1dfe5c6be7b79000e29a203c6acb75d7c76ed053bd74;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hddf84ae244d9c54b66a7ca025d5618dd31e42534dc4d506705567b74b1d6c1d01b9f24074671de94c1dea1740049a7b6984716a04ea4c3bb82184ec04;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b017c0ed4103478c31d4fb22da57285462d70148bc0bbc88deaab4826f86656d13da15ba6f799e945d48d5eeb9c97117bf4e4ae1acf46d4a9ae9fabb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf240f45f287c0a4bbde3204958b97b5c4d4d59581f14e674d0efd48596038b30bc2369c6ee6f2b2ba8671fe4080f758e9073aec57bd2a26349402aa5f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he62a139299be94cac146006d7aa59ec8d0483f36a75169a7436aa534eb5dd6d298e22a0357e7b8fb4ac0402b9e60610aa561431cd9b7b68dfa790f986;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82bc311fc5a28ff5f63deae09f7e39df8021b0c32e6b9992c8ce981abbe5c1e79c6c8b3ef912feaa334b12482e2228c1e492a0034dfdd62b168bcabc6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53b42b2f4cd37540db321656d7a1ad8773aa5611abfe4889ee5797fc69a3b8ef245a203794d2f05d7c015114d5e2e7b1b4e7e64533de1acdefc21b2dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a1250230533a63bd1adb91ab2fe401baff3513c2a236a3ed106a959598c8b23e3810c9c8248b9e53e44129752bfdce1bff69be8129c6a4cf2474b489;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb30e7027bcb149c440731491c16237539fb9daea23def009b308c1fa1b02f5a0ec60d7d608388701a9c504a3445013fcd010190d56133a77ebd1db820;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6edbf3e6b7c46da256f8210050215f5c3ea8f97f4cf66224861f705842ea9024ec5882e05a1578679cc663c7fe350d7d9bcee708419f6391e32f3f2fe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f87f84233f212c3c3a2206d40efeb361833b58aca43cbb825d2cc36a9844b107e5d5174f975c05234e2fdb54746e5fd1564659f4dc4eeed14c04b4ca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc12355a833c0e4c48774be7edf2220c331f7a6089a7dc708efce9ae7df20ae00b801d510bc3ad6f57b0c65bac725cf4970f774731b13e93d7cb17ba2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hadcc0109bc15a459ebaac455eac1d3a80fc3c2428c7f15462571ff1dadc8da1375b56b64ada718d05d58a09bdbd6aab69ae0b4cd37311f9a5422dd0a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8db8ae03862065d98685595f61dd299974994a475f63b532ca6b9f50b0e6b7e17cf8f49e5ca2752b0e4c56942fa1b5583a39eccb1429a17b791a03509;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h194e30da0175e2850632e0123a71d5d4a9ba05136573548f44c4712e2c1c4aab418c71dc9dcd1c2fcaa23f98864b37eced23447e5c234d6b58026abfa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h782b3f955eac64416f87ebaec6dba33b52d6281d453f2000089521eb943533a0bf2abe3cdbff749a9018684f02be294317814b51bc8c9a21e875c50a1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31d44a55749a78ab40db4cd085eb12ea8c3f34d77bc3e2ee90d70e0d56562fecc2ece63c1103590dea74b98fd49ea3f144156dffd85fb794608bb9f84;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fa36c8a649c57f66b4a41f34468d5fb181d47de696b2af4a5919cb6cd8e5a9b4a5b78fd46b61fce84d42f1ad2b25afd0e2b3865841c8244c8eab782e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdfe1779d3698d676bc8af79c27b42ebda7a50bb63327c9c707b29243f64c145d6e50ffc2791a7de17e3a73016a6e3adb66eacfcaa1413097e509d70ae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fcadfd229c96bef41d37981053b0edc42c3fb44cf0f2ef5b1ae3429aaf62e365e5a7ef1767fcc1ae3d4f430bf7827d31c75d199eb7abd8588f2e1872;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a1fca25781e0dc2ddaaf95ff9b619c075754528930cdc29e434c9e21ac8ccaa9ffa24beb60c65b2624780c23a9e6bb6647088973d6b9c1c6d26816;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc808e6b958384b022b19c260a4ecbd8b5f149ab7c47b15fdca6f322d200e98aecc98f608b249976fd5d877782dc550a8c0118196a045e3942acf8650c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9928d8194a3b8fbf2d7b82f086ffdb76afe4610316e295f9d69fa057457276012493270cd9d2441e8b6a14e0e5fa520e26d138fb0604a2c0b9e68a9bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb22b94a737ddd6db7b822b102b1b63591ce35b796cdbe8488697b418b68533a063ed92bde59e7592049a1adda9e5830070fa44b32f34b1226ee55b778;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h679b9619fbbf54653bdb29f2120b87398c5f4c015668f05947ea06b93dd642516fd86e523a9f233881e3e313811f8a37cde9d79ebed6a3b33725383b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9eea2b7d64a8bbfa9f49d9c6a14be63c8712a3c13bf77ae0ab19d4225b7b58ab065c654f9f3c2ffc657b9580a278fec95239f6b08edb9e0b3de661b37;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d409be291879c559c29731cc151668fa221ae0d77216e5694072d6d7aec94fd26b363c61062de7c03bb5dcd2e132b7ea8581c523dd81636b185e68b4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h623cb2870c1de3af6c5b95828d92dd3ba6b7cfa6a2a0c826ac3eafcb9aeda4e075a08afecfe61796d4f755ce48aa1b9886fb9e703dfa10f0c9d15c91c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2cf221f967ae12ceef5632ffeb3978678216ce0a56f67f296597dc6987406a9f69de2ec7dff4fb32a226cc5d4f5a7277001314fcd41808e59b2c87d1a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hecd0926a1fd69439b95f30cc86c16d6dc5d1174daf4174810df7c764f661a87629de59a5acaca6c8878ab358e17de607d084bb66a119f202eef3bf4fe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h246c8a0edeea0bc08fcd862d646448b28fe826b0d3fa6825b49daa280476e19d533fef27a66c9f56c382ec58246651f359ae5289ed3dc7450de07ece;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbabe19eba1ec254477bbec3d0bc54ddffac69bdc6a90251d5a01e9c1bed2f0f9469b521e2dfe5a135ee717ebdada342acfa11047e54f2b962d98b86be;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h681fdc66116cd85b3f25977b45aae23c80fca89fbb338191b5107e0c625a0eb1cd6e0bba0dfc919e86ff36ed8e4e3abbc283d32b9cd79decdb1bf8756;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b8cf7c2963249533cda904e47da35dd24255d5d6383219063fddca3e2b5520831e7d8ffff7cad3841eff4af0983e60f76ad1ae9273410de48f16d569;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92745fd0116b379f145c2430b62e40f58e81a817354da480a28c871806ff554a98af66f8becd29ff46eef82012a655468a42da5c0ddee77e3b37cd301;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h312f9b1c1ce770474d16af50b55a6fdd104aafb7949cce772b5a01211083e27fa90fe6375d6cdaec2f9c0e5ba68d306533c5fbd503ad53c9634e15800;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf896bc2c223490e49d15b1640d1590132bdad0a89cfcf15f69656b9734dfb31aaf93707e51101948dccff9d92cc925594b80a94725220596203cf4db9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he62b91ec0ce0c7875e01a26bf311d13bcaa7e09a9f90ef821a9198ae5c65543bd1dfd1ed3269a783c62a2dbf24594fa662230089df6516bd0e222bbeb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50452f449c300e593d201813f77facc4748be76bb1136623617dac85c30197128414d4a2c0fd36022e7b7dfc9f4252ce3a3ce7b22b495cdfe9b7374bd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e703da1fed9ffad8993964d11d1aa7c711ba476f1e337e8cbe16a2b35e3a3843ad057d367a0f65de503758af4cca3f888ea2941abfa0a3ed2d0b3e9d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b5241ee0cccf84ae0d7e1d9e53aefd45ccc2b72e9bfd4c5b66aa91384d000b6fb711b5bcf143947e6853487d1c11644c377b199dbe8f45148f02aeb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf504e06d2c1fbacae66afca463a6e6807a83e840bf6fbd21b088e1638c46ea4246c1154c8b5f449e5341cd40536038b1e2b8618699e213aac257c16a1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7139da4f48903378745089fbe4aee0e377b663caaa1a0c4395502c701bc292fc4f177efb97896b6dc7780ef17f4d8a8cea456998899ff8a41ce04bd42;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7eee8da0b321f9892a10c6da054483b92deeba5b2d9d3853cdecbe86ae0e11c16f4088a505d9af27e228afd497cc444b8283f24bafe884e8126bade32;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a9a645f41a236119090f56d42b1674e21957f8b494b26ec92963e11462d3a4f5ae54229ea36ee723e0e7f43051dd7c26032dcfd0b227a8d3fd9fd618;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1480144bdcf241c23aa6c00f7f729f31c410f88a8697a15803d467a2372d544f4c11e79719df24fcfa07702e9bb626cd909208e21f67c04d21febe70;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdc2945408c399f18864887173d51a39849c147ddadc9eccf9fc0321b747cfa7a745664f9765b0d4188d584555ed3d42b746399f375372aab7c0c65f0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4036a70e7adfe4681227b9a8c71535cacc3b03aa42a6046b0cb65683e9da130e05036b62900f491390d4757b9c931fba58e5e8d36e3eac5d6e4539dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46143edadba5bf45b394a6c8cdfc564669d961713761ada899f80e4be4fc5f4123a606345a2b0be578ad4abf99d9535f48f6c169713661abf609081c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1707e9850406b607861b571721f9b41fd86759db6640e96f86be09930a188a7be43c23e6c4a16360453c1b82e79b9cab675899274e0faa8bc19b7d6d8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h297ef316fbf0dce25e4725c8c52d181bd8f18c4fc48de040a7c8a19bd80a965a57441478472ec05a0d9e3cdfdcbe281bc7402ff229d23c5158844b248;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec53a6babfe3397d08f91ce1ec027227c3e1151abc67519da7bb5a559931d2e81eb3f15fa3e9f4117ed5c172f87ec328dbcec937277c992f9f66f1716;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2dd5beff327487a97b39b8e76bac8381881bef252ac8c0aa9560c113b99a2d1cd3720627e5e98d8970d1e3a2e03931ec4b63cf038a12808eddbe45df1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d6f4f55441c5cc715f973345604a085fddc99b42efc909ce1e717764b6e5d8256ceac0a0d0d76368df50715cf80f880a8680eed5e2ddcadc912ebcc5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48aca702102cf73e71b31e8dfb0061503491d7194684403305deb3f4bc32af04e6451eef81e610e3cf69d5543e2cbb4ce4ae303332a02bedb6311cd69;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16422ced6da64472adf5087cf0d76a2fa8c2aebab1a7c88070b47016894b7c337ef117ea4e933b3c2b3a1fc0048acb40ca5bef7770e2942a40a1ca6c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37eea7f1c51da54446bfdf702a7415867882cddfee6a58acb510954fc5e9b291fe68b8b1e394ba8c4654d6f1159f90d0b11ce3923170d8bbdbf300fe7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2974e9cf73050893d6e88369e5bbc77b99ff2f92c196e3c4d8b973aa77636490ca2e305bd1274267dc36107377a00300dd5991896092c14765451afd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef5928a32b450ea386f0e3b53fefdd50c65b20df255bc788d5b7d84bfc13b249d5194733e2fd68280407d40036d3638acb330ed38791d3c11d3bc9c62;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd9a4bf9a5c469d71daf3e6b3b2e8a63e16e978dbb2f8572826c1753c280ea235b522761bdf48015a6b81244f596a62b8fd862d0110e3bc43a2b24d68;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39b71de2255ad78f6e7e0b19f50d7595fde105de16d5a5b7172f5480d510682c2731977234fe2336972b1194ece7bec056a182e6d537861ae7af1eb22;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacd0714bcef3ccbd60b03f35107ccbd251a2bbedbf93ec9532d99478bcc0b02c1f133743072db10074d74f245d47d007728dcf007ab4cf2f1ab916c6d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2b73d2e1ac5cb7f7d382801659e0eb6773ba4fc1e6217dafd5d5f49a314da90c6eb2d5c5948f4da302278375bad2396258df93e76d533b9fc14b32b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25c5deb2a2170ea692e6a23a00ac2973a6b7e98a8e4fa5fb221d16579f08ca2c673d4525a17cd579c5b5baee8ea8a1239f9672f83ccda817f85fca83b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e8ccf2eac77c56a609ce1a6994e06617e1a57e3ef1437897dc807021dc9d56df45e5007622f12e4f85be1139c29cae8ccc38bf938c053caa55c34083;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha891582df542a4f792345aa7c0a4a820278c25161931412237231af6ae1a05a61157f3efb20a8000727aee5b4f2764410e4b1f91cf5be404afa3537bb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf26fb9853e3b86850cf05b2f9bf53a63e828216e42d260f72a29d13b0a5ac3c01d06c1ae125ab5664b75ed2d5e88d7ddc6be989cb7b4de211fd3605ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d0b162c78e4b21d0dadfe04fdb3594a7db95f323df75889e3c11b10124adeacb933c83becc596c4fba72c6d696cbda6b940b9767b07fb79ae9a293a7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92f8c174563d7ba79847afb9cd94164e62dc2b8ba22b382b8df7eecfe2e888375c6c7601c18b16ef6ff68ae7e263aa9f7f419662cafec2e2a0d9557a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb23f07e565e2b1d085b3adb63aca1128d5363a94ba721bce701f24717ac042c24bdf8ba41117742426512c3aef8faa0c1adde7e0e61c0be67e20b6f7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha43e76306a40b9b56a1087802f6537606e05cfc7be5f971c01d711f7605ea325c038056dc47d76effb0b287bf60eb10e1d1357d15fcdca3e7183d841a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc7127f69d6029c97dcaca11b361458b4d2ef1ee253706bd60444d52c4b1abe38affc829d7d737b0ca1b85ec1c2c307de61bb5f8d2ea525c660a19d5b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26895c33d40819b4d365e94cdcbbaad2a590ded69aa7a7aa8390169d17948e8f6afb79c35210da86875efa678562792d1198099f51029fc39db900a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8809e0ed2c43cd5649d2a51af03cbff45a89d0bce715067f0e8969bcd9b4638ca86bf749a26c9c7479f2dc3abada76455ea9c75391de0495fe28e50f1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h207f2b79890da7c652316718db8861d9075fa95e04f285fb0fa58445054eff736e6efcf4fcc2aedc627f147d41a1636c83fb0343b75c69acff30f80d6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b43c7a3737efe135ccd59578ddc2c88c1c7868a4b5c891f4d6744fbfba47cd1501e203da9d2a937550be9fc0b53a5f83657adf16abd7893472ab90;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e7955a36d8a870dac588ed48f296ac49911fe93436ac8b1550b2cc3dda7320c0b55ae9ee189ab0a85ddb4cb4140245f09a125e4fa0c949ebeb2e2af4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7fc8c0c71c3254671da2890f5a5637d0f4d5ce9bc932c865b42b616421b35b8212bfb7353664673bdfb1ecd0b961c3eca38fe6bfc69e23002860ad21;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21a732fc476aa0ba0aed4e737b6f6be75ad825740d5415bf0872dd09b772760f1a2fbff044a92d2e47264d8337741ca47c085330651e18c3609d00a1d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b474c9530069ad0bef882145d1666e8a73fae7d4a33186114c9bd66b83556ffd0370ed9468820f239affc7ae4c7774ed89991f13b5a0149e251d0ba3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h985c307d918e0f0bd4f6578ff530896b5a956e79dd7d314e18afaf9d85b2e48ff4515f655c880800d956656faa9890702ce8d4e0b54a8aa09aaa5c003;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94b70f9dedd81789cc5c548cb46aa6dd6d7ffe7eee1de6b839f30a04d6f7c317134ce9f433b7902046c8348cc37837c250667e77fcbd737f7f14fdcdd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94f5a84c7c25b576ab669fcc5b8613d73f8a9912e5cef24e0b780217bf7e7accd5593cdda4c8bd12d446c73bdb903b81ab8757ff7f10ccf3844fd980a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a3ba9c501ad6386b79b3b9751ebb82078543c3b5c0569036eee8dc1ae86dab285d1e762144d08601e40a10e13f5ceb3009a2cd2254d667d6bcb85c6a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he47a7ef1e335a7578b97d2fe69140b913101f30fe4980c1f00270df45e830418f5e53a2c01a7d6247e485f6c370a0f053b26a687c4fda90dce70d694;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe88127791c0d573802a1ce9b381a786363496f964a9649238fed8bb285f807b01c911d5e6662fbaab88d07cc05b1c501739cd739af9e0985c1a4be9e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac688f4627cebdc49c03bed10e24ec2c11a740b9ab8e0bd5e351929f7b702ee8ce6850b05bcb255e21c6d148a60dc2b7f3158072788da5b69b553aa8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ce4fdce942ab868ec2cc80c3a68d9f4c789d4c13c2e82f17278668f16f3980fef78959477aebdaa9a537c519a6ea6656c8ec67cf12e7122477179dfd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80ab1f9c2aa64d7a47fa4ed6e0560dc8821ec6d16a93abbfd855e26125c8bf4bcd4a5d1a223081b20f0079500d45fe66c7d8cc6d5c2209954eecbde92;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63802a1f9874a0499b3fd30e760ee3a9744882ba36dbaf10b5b6da5f61fb153b9cae8d63b46fa703b2766e8651cd23c600b76b50738f07c354d9eac2a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3e7782b6348eb216172636d8d99eb0f71e503c721628719b8b0ba5a24b8984edce69e9ebb2ad99de955b2086044a84f77bafe092ca6760e3c8974185;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72d17ad185de36f3137f83089c3a72265cd24d95f5284c0ef601f8d65232bcd86e484042ef8357261460d22b98b1a2f73ac7ec08f572164e015c676e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a17a1bbd44597649af68cdf68b420dc193df5f5efc1440316d297c146935cfb1adfa1e210b166a27b0d4b9105fb45d9e09c602a4512ff2cc52007ab3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8540282e3f50324143bf42e08913616d361a881e60277679275e87dcedff3144e7e9a87d5a746cad1221e7f94cff7968cfe182c36c632510321774e31;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90ed0e6b80d93b97aa1db26794d72362b24b958abf0cb100d5c14857c8c4377acb6bd0050b1c9e7574e534072b06d230bce418ba436c97cd2e7230bce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cb167fc7ad4f86a9108623e4c3e33a38fc5e3eda4e554392c1afbe1af1be04793804e51369846bc1d26e18f41c7c1746740fd8fbde9951aa705acf74;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb80659b5613f2a178d702b9c7f1393b946eb87e1e372483cfb665d07b46ee6c56465d88a33fd0a7a5d9b1324569e8bdb6e5bfe9183be30d82646828c9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heab23a64b4f9b40a2efb550a9842983df050d9fea9e78ee05ca575948362350a070170ebaf880c3e78e2ee13b953ea7778615c20693b4788efeec6745;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0dcb470daa53db7d60c16c9df050affaa831678c99834297c6c748b73f79d3aea88d6f7545c061ad88e729f7d1cf37161fac73392d6a8dfbf89bad43;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91cdba611055a18ffcf40c900c0efd224cc27483589382a156ba39a2908da828c43196e451eb0631f3388e40ec1c643a7f72697508ada3a9a7f09838c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha49a5de7f6030751ce4d2b301af72f57989fc0f97b0f0ff1b95bdaa1853cb755148bb2ba42a93a060f6487c673b2d8ef917bef0cbdcf639c4f6ca874a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7d17d224a85057fcb1fa4ce01f8ba2c4c9c0eeef9bfe9f3789e63fb52183deca02ae5090823be633a0d3e2c22d4a1d0a75ac32e6d6f3b79b3043832c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4e84fc9c0ac4088bda8f8fa5e94aeb4d3bb3bfdedb65e74879831c8c0034a8dd5ecb8242d874657fe97504ec09f28da2b82049225bc5eda51b0054a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32015673b12d81eef99c16d00c6600aed6cd232e924fbab178bf2abcb6db31689449cfa2ad0ed72e0ef948e62f13caee10dfbc304c791bade55e71b97;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0243a23b74562cc2deb4557b69e77820450be4c95ef48b65d9476803cd0dff04735cae7a87f23495f7516e98daa573a86483bbecb1595a3b9f68dac6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12e24190e306fbb77395e3b34d6f987614f621893c3af4a5682681c04a6b4134ed04a1590a135186ba838047faf21a0d392b11211bfa2b3045d9c4d92;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h263161e671a1f533c7224e4866bbd48e1b4c6db2faf1031ea4ba10862ccdd3731ce4b4bcc7d537304c8efbd936db446dfc885d1d509156899685998b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd0b3965091975e4b80255dac733bd71a0843c3cabf5dedc01648072cc848d5f056f43d28251b40b6f6a5f340af8bbe1810bfdf550f68fd193791289;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf61770ff96b7133365067182db6f87416098f7b3a4d83449d13715d776e3c4fbb8e1710c97490bb119a622b2b0eaaba796e893be9963f82915f6e0957;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h346b35cd1b00fec4fdbe721ff0d08792d411d77362e3cd589382d597054435943b0ede2e35a2a83254eae4cc7cfb1d548784911995e96ff772779a879;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha87630af408f9a59976ea5ab3cd8460c6381b3eae9c8c51ad1eefb21e4331ac2f08c1fcd3f014b93e3ef19f4ce39b38dca6d323c8c2c4d0f0a65896f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ba27f182db710f05006959ff3d8ca39f6fa91955fae1e379afa6f4af617796fbf314de19417a7c610e31e2258a68de283233b1ab0a9d34a79a421b47;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha47e9b25c2b9843fd9c32dbbd68260b11449791898e967cdef085a3fa579f10d561ad30d0a3b0b1d0336fee3a3e6588f27dfc978fcd2b10434e03a30e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf907f858b7ebb99554e8b4fd20a714a972ec76ec9766741fbe86bd4ea8ea3f7213256d36792cfd5210c9e46eedfcfde330dd9a8faeca73de1445a635c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cbaba555760d60d17d532bc3d845dc3b9637707bab384467ed9fedb78ea661722f1006325972c117fa2d27e8d2f7310df9585359248ba82f6060e744;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcbf4bf47f8caa573c32d27a4011bfce66d5cf4737cc832a466be9f6b5e119b1bb8bbde79350a7d928ac9ab2132804b0c96c6660c30cc2cdf703d2eb43;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h135acdf61e281a5e060cfb00f7860a701f00682d0422634958d4ee0d7c7892d489cea29b05b285cc603dfce900d5d1faef7eb07f71cb82eb96f65b210;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bd33989e15aeb8d965ae0a7cd84881df8a858dae61f06fc0697b35794ff9d0a4ef9a5230918218f0af498a4d9ea2984250b6684d20a55367089f3ee8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88974c5502c821f647491b396700018a2e18117a13f747a673e4da8b341dde756dfafb4a3c2b9c1bbd80ac9e3a7714abd1caa65fe109f12bbaf9e77f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdefd2d1b97fa3488ddfe7400c58ecd35cccaa8f35b85b16ab36d5cad676ec07e79897d5770b0c00bb9c314d72734bbbe141746916747f974d56a900e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62a54b1845a1680ce1e160e7aa7304e4f3baf5e07d14b3fe6d10f135ec460d3af057d436874149a1bedabc243387f10ba7a3681dc597e9e4b16b8229d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hddb5d959cdaff58b8848b836fac23498dd5c6dd0aff16ea0e74bbbe5890a2f2852edfac40bf867c07272d38ce18881cbcd7263899f2698fedb0be32e7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66be8527fdaf9790c30c743afc3b36753563ad936b8b57aaff819c8672fcf95150f057d143ec5d265895b01986a321e236705a29ef79decd4f7c4b41;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5032d49761b966f66dda9a72bd4112bd536e184ac4e84e43cc545131cce711a510e96911e556c7d0f2ab8099a9f4ec2578f8b276ebb37c5c5ba9b5fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h967085da7b558fba52b4efd02e14048b77781a563b8a1df473f17104d47a6c4a2c4fe72f54f52a27f74f9011bad1e5f752a82a9862a32111009f0372a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37857c23a80ac5bfaf81f0a34a85a9c741adc0a40306814c4874594790b4302e657039de851b7f56fb8fbf0f245db58231f84a297715b668771113235;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdda1bd91caef88abe9415fb65002fb64e2f2aa982c7dac1f44424069a4fc921d19b41a2425ad402f854a8156803625e2f905aa3c8bea0e72c7f28a4d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9e19e75735dd2cf289131e40a4325453d966f4c7f3e4d1357c28d0c88dc51807e571dea1cb595834b03bd8c5deaed811b484e348acc8ab1ecdf722b9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b978e63841e9b662d5c8cf9a02296187ebe828aa0ce9e0f4aa30a361e6561e073e1998940179163a3739392d4cd79a74da8deaad22072294efa07ac0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h966177d687fa067f71cc47ec24bd8a063f61bebff4390a581e6096e8096148882bda8434ce30ed7a75ff519a555ac327e2ebafeda4a89a5ef102afb2b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd29145a2bb6105b64012ebb027da352c5f855fe4e0c74f6590dfb7b1749b1e0202b019da48d4031b1d0d20f9c59ef81e45d5ab6f5bf4c70fc41e0d99;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16c8b40aa882b212a0a4c527e9f22eea31f708da36678a43ce738fd22868fe5b4659fd768c6da030ffb679ade7acce44f5d42bd84076cff2ffb550bdb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7761cde59dca7adf6af5e7d30b01f17646396eea97fc8a4e3231d5a594789aecdcb405d8ec17eadda6c1b7e6cd5f51bfbd805cb911e7f3e5b58fb96a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h525a2308c3478b608f560632f06a39d0f02e5e80d8a3b9a3013d83b69d47e219354b2144e10f418433db9b8d059e5779eef2ed1f518186116e207d02e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde602edbc2eab3ae9c9c059f40ad51d6b9fb367805f376c20511c84d930263d65e373551bbbe5bd2528b1a63c39473b3e1043e62c265ac8a75b524231;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hadc8299995d9498cb89bbda56f9666c0ffeaecc97431ecdd9dd21ba2637c3fcf498b50884b90bd089a46757b63a10feb109edd2e63d07383a6acf429;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3a815d2b4f9036f0edf004052875c4cffa82dd834f83b8187c7a7708bcd85713ecc0e4c7f15954d69e2a3f92401dc959633073917a397f111d85ce9e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h179979574a51dd8b1dacc14dfcd8023f978e361298a9517924a39b1ae26fc6cb996e9afbfd0316a8f0ab5375439a93d6ca70dda3dbeff02d7acb453db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdfcfa85fe351dc77a399a83490ac19fa285f560453a47310e622488f4abee0936334e474cd4ff827b45e4b2602615c403f228c6d7b16de6afb3bd19ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1654dfa6948fb74c03f141ccbef4b7348b967994f487e982f775f12fd81e2a7f83e3e5ca198b900211f03ff3b332aad10551c8dafbcad653a720ddb44;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5176b5ad9f5e2f82b9b7c83c68dafab13ca9241ae83295212c959bdd01653ba585d06c921b614b9bbe42bd1a7d02462d9b80453232effe279e44d0100;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a4065caba420aff89db5822778621fbb44b5fddc315c18d9613427de24103689d0da5ea686f0667dc4d1258ac260062927b1fe1060f37bd2c612fa60;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2550999248aa9acfd6758c0cb49b078136e60de0eb9664a56a843edf2c48872f61aebfcf98cd4906cd2ac30c68ca205d6d8f497269c3c78b2c98b786d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e33e7186a35514d4e2132967e27eb3c5ec2396379f8d5e874ddd0030774dafff0ca683dbe5b545298ec0996dd31c99664ce0c93f7d3197859e8d92f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h220a635362c02c5f1d59bde656b83048f94646e02cb2b95d3eac4bcba3e523d3b04bdc82e72628a93ad5abcac8b0a36a18e5079dac982331e6b631e04;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84d71221168326fec932e8534fa8220b7aa512d4a01659b46ee620fb4e947414dac67359725ed86f82677b2eab012a84371d871eb5d029bef2b4e85ac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5716b4dabbaa9432563477aa4cbc601e2f2ce222e78c592429b7574af655acf8bc2f69c228e57cb6edb384a8f050094e74c2a93d3fe3a9be4d6ce56b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79420cc6242ebc378957e0e5dda0add741039d877cb78511e26db81d3608e5008d3bada82ae173d2bb72bb6d8cc9e16cd6bef14db63e7c10d9367f26d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5cc82c0e7d2741ca9cc6c6245cd5bafd88819ff402fec812c21086d5d25d75cf07539f13bf34079d60da9c9e76dd44876893489ab4699336ee01cd18d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f25d29087156edc706a2126da05feb0e72974e38d83f54a7c3238ea7d568478abfbd4316bff8d6579f3862493f365492e96355a10bb47e94a0568e4a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7977f11c10e4e40c3b58afb661a65e44d8a0a4a3ef4983b109384c4c81d5fef7653f6eaa538604282190feeec1662d5bc205f7c790dd61d8e58f36615;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c15fc2477d7123c9929d8c9fa3cdffcbef0487b1252a764be3bdb055bf1a83e89666cbf5487c3776b280e74387e641e27e55aab66fff63070d0f7a09;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf34bec9bc301295ac8c27890af84f55d05d69b611cc41a3551478b291190c6c833c69b9e359c558eb66361e5baed9b017d08a7dda9750cfb9d8a519d4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hddccbc47fc916a507caeb712290b9747ea5fc93a59b9bec7236c009c68a36d3a3a74d54dd1f56629b1a67ca9d532f3d1748d5aad051cf246634592f90;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf028502e3f95f370c61d1e2e6371099efbab423a0cb6234439664560edafd63d4096f5ffca94d4e56f56277d31141bd540ac358e76d190f4e1692ff18;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h483d9a04f68a360df88c207279520cb7bfd1b44ab3808689b8d8a0a925a6794d93e8ab81cc0c99b160c68038be4fa0d673440106d921b0c490b2be7bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haefb278ea335bb55d6a2b6141a9b365bbcc8369d17050fe6b33ddeb8654a8d43726100728af767dcc70d2d67f4a79a73cdac871524d3c00a6db2c58d1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a8871bbcf5cf6fd32cd377d6dead29d9011e221eac341b36ea2d549518357376c92bffc7418cff90fc3ce7802f9e3a4d570b8d425e523abc1c2eee68;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h889cfc0f5e72d7b9348d219c3a92a19cba70ef4e9dca88633a9e6e29bac03b6552f4de542e59c91abbbfdfcf3f8942758f04b7056e946f637b0b65f29;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he02aa2591522b210951254bc9e47706f987e27c0e2ff5de328f47eb87db74cbdc47a40b00e921b2923e53cf0385bf8071c24d4edd3381d670a7fd0d13;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ec35535e743a9cb73d555ee9e9fd6ce369bcf4eeaac018f06b3fffa92eedd29f3d9a1f5969685c0f94cf7ac1abf78791bd1dc0bce9af978cf07bb6b2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32513bf204fe936649fcdfa1143bca5d5e02a14fcf0be5a5901c56f49da22eff83f0b56dde13747e582a662316071f89c5df9bb9b2f8768e2918177f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e4698ffc1cf162657cfa975aafa710794329102512a6124c1bd42be83b0f8b5d7528878ea7051381908357a6a552e61cfdc849cea957ad6cc74627db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb710592b2564a20ba50392372560b8e0d621350a47326c00fc88a7c65f6a7d01d8160c5fadf5a6272af26078791a4613c9162710ac9f1b52daefdf490;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he409ce8430cffded244cb597c9d6f420f70ee407e3acb3f6fb7a9503c06b145a7d8c5085c9194a784cceb863aba39e74b6d0d7408b8837bef31317580;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f2438429c3ac978626150e59e6ceb2ed8b721f0d75a6ed4445be32e9d389bf92e9a4856100ac75f823ecf456133e3dc508bfc4013a130d009a1805a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb76cc83cbb8e5e33ce3e58cf6e0d3ebc65724f09ab0ed39de26b466602c709d07c4ce48b64fcec21f3ce0d943b958ae7125094cb9ac7f166c56583c9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef6720140d030a1c20bc89ec3fa184ea153f77b2eae71afa75fde3327f5d5014287a0495ac9695961436ed6f98f0a9e13dde9aeb354bcac815b9fb669;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c578604d9bc3ea00fff530e78f0981607fe746183310ac26d5806b6b26b68c66236259ae4d560c949b132a0910cbf942d05e6de0622290d89b40e283;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb7b49a798ea004d1d74a4b7e6ba984150ff60c04b50f94b55d092dbccd2c356d06353e5ce67cc91f1d74612edec6becb4cdb1927bae90b186114ef86;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f77a3e8fe0ee89672e9b4e0178ff05793865ebd6155a328808ce1677df6f33ae742154881293ea89349cfde82c11886bf8b05cef051c38b12d122aae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ed440d41e464c3de36b85d02f638a16945a82ed953c5e25a76528bddf3bbed4809e71ebfaa1da1be4542ce2a7082e124a6f41eae7944e1a03e10a705;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11594d7c7513a524dffa4127d0a5127e0f63afc49213b9a2d8fb4ec11ed896895c2a1f405cf7223e25d6d760098d43cfa09c69a06a9b9730bc818b287;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac0093647e67c226b546abf945ac87239bff0fcc3a7ab9521f523ef2e757267411dc447a66583b334fefafc43a16137233e39705b53e7af967483c37;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h236119ce544c4073b51060ca8298acdc59646ecab80f527763f209f6c0c0caf7dd6ad1445ff02fbe8183dec3a7c5f88db73a6bd58709fe55be98ef450;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d8010efe0895127a4e7b5f7b0a92ab9b4b2b3dfa9dda5b742d720ae6eeb3e117e3a1639179b2105c8a8022cb36ff456d5010c75f7ec76d2f15c9c248;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14d01156ac0c70fdecbbc84564c3b7c23f18e5678c11153e383e4ebaa2cb0112a16645c6b510a5d47da580113a24b7a6fb0c6b570aeac833eba401728;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e49b609df50578cd311321af00c36c3b6e61030c91b85a667be42d78450e2affd3d580dc21e9db90f7f3d04c004d9d56218fe55d488febea9c688173;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb1d621e8a4ded0aa310f27ef0d8166279e70d24c9ba06527c70f39ce8bcd8461aff6364aa29baaa10252d49fe441856e8c22969acd6ddc4a314de39b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha047fdc6b49dc7dc877aa799cf38d8bea579c4d8a2efe6ddcb0b0c9a74c076ed12f92ff17d38a5a036beee9c19e7e85c056a7881d1af129a5bcb41143;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ff8a75093c1d4fad1da009721c51a2ddc30443cf2c2a2feb7a1830692c0cb3446b15aeb4f23a40e22e0d0d7a9b6c0d4e18b21403505012dd58357271;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4127a4d7b4ed31074a6a7c74aa44e21c1de1304df54f51b69480650c2e29654e1320298f79f92de15d02f838dfee94fe8e51f601ec0003241dda966;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h399c13d9fabdd4e1ceb2bdeb0cafd3f5209e14130ca60123366520f7265de3811f597f4420e3e809fb7a0c6af1687eef787d063ad02fb9320d6599221;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdbfd304fedd71eb9a4d09544d4af1e814545a7ec4be145e77e7e1987e5e34879983cd680e945450e6e479aa9bfa0b7360aa4c23358acdf11ec428b57;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5cf42d5111b054e038f4262468b3eba7302bd79b03ef56c2f32857d875f2c97398c5c20147f6018f667e0bdb626b58e229a8d55089662ee5d6adf437;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7efb0bdd44346a5ec5c17554f4a0cd836f86e8d268352b9efa05ff5a87201ba40bee53f2b315e0bf45a06fcfb8140b6ef7dcc9f70ebd97b6728aae7a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8ec8d2e1a923499ce2a91e6093aa46e875348eaab2e6962b691824a02f266e598e8a3fa7644e6479d5353399f86d82e4750d2d2b4adc837bdc356569;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha99b80cd109f1d9ff85e854d2fa7c46c8ce8c25d55a1de2cdf6956e139c0d085b5e6607bf6472a93ca22abb05e620947d136723edf8aff4275340c01a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35f2b76c0e12ea91a248903f54d4b5965cb78585636a6534cf78b05a2051a47450a28417ed6721a9f02ce98dc6735f94e2ce03081d66909e889ca330f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5fc9149339d8eef934787699aa6d9f6ab91ee85610b6f63b39dcf2931ef2bb1c2ae29eb29214e33ebb0fe73fdca2b84628441eba72c932f836c2d6d22;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ae56daf64ec02510762de5c711e6f98c2162f51d676ba693a76ec4a490d9011a26a55d85d8eab0a31111498c0c4ecd03071f7302e83254e4cdbf9fd7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc254e7a056ebb3bcd50afb85aa4a0a00e77c6d7ee20e883a50fe95594194b4475b771342ff37f1baf8cbc30ec2bd4c900052e305d6bdf9c35bf3a3791;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf92e1e8c7d2d23e2fdcc3bfc8e0aaf684b8e68e3a5ad5e27e8029e081c62b68d69ab1150f9149662f83818823b31ff11bbfa8875efa17cb60a7c62edf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb5492d3c301486fd2841f88c9f923586b4067206e81350f670c8fe3792d1464b2e66a633bff48456b234164f7c0b38fe454093e521783fda445da1a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h386500dff199f4d8d4f03e6e6ef1b3b80df04b8ea517bdd7e3b523440941c6250b16aabb2a347f6ad48f4d3da5232f38657a86b1887ea74ae4e13f6ca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bee7b827b1c1faf4c9ef758cebe92638c215bc56d4380d81cd7cc799eb1864a73ebe07e69c749b2003e82b7ffe930a7ca9052e7b1ca321dca6df0dcc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5feac99abdcabb3ceb534d33093317725917dfc162b1a40c4b17c330d8b3e527911be270b1931487472fa41954cd2c8b6232d2844369afaedc0893b9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fbad473c1acaa361b2cc201c7ea1a6b3f413d375b2130ce38c646f38612a306bdf317ecedf4094e1e9d722de214cc77d9d2221b9fe2e0e6b09cda5b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cab5671302516f6975ba2e675c018059b968cc6e98bfca36d4a5023363057de1e6d46242e826aac96a2ccff2975bc411710d43dd3c0513659f9a39af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb413534e9e91ff686dd319256ea10c200296e60531950e679505155348763d5e3fa3c1302d1f020f1459c15bb56d863374865613909f8607eea562a7c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62f7ebe16692b95dd11ee75e728fc287b8330cb84a1b66f95401269511f6058c0eb5fa53428be537d1ada52bfa173afec361b85b82387e0cae2b3fc4f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2220137392338492ded9f13b14ccdf9653717fc53fe0bcbdaeb5a9cf9de892d7e412f434bfa5a906ef14abef9812ad7ea75ef28fd0e89463b6106c040;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ef55aae4c89fde602f9d24d22c56dc9f8ceb4ccdad22399300bdab68812d9481777e295b7e293d462f1d2711c2d989112b2165a4b0cc97968ce520c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5311ba1c5ff97c4b01a1ff27a129811c9bf0d6413f5560a3eb48f916157d874fba58aa338b5c50822c17e351ac3df19032099db28822cc8d8bb75765a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1354b70650219e684edd10b622d56d94af88ce306e7c81ec4695d0dcb547164252a4ba0924ec4677ebaa5f33dcfbbe0cc3949b7d8a7754d03f5498c55;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b3e2a8734f4450bf45b59e6f9b983719daba833a7e24c6431995177dd2605a7a30466ad394e525a9e1f70108a16d6b669faa2889a7231cb7791e407b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d75b028b3543820b595be7472f5687b800f94efd979a10747dbf0cf85b5c2a1a831b0d9416654048132fc9c01a210f7a9ba06a514e51e30f4d79fe42;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13d5cc76a3d2395453ce406b525e50dbb5896bf8cfb3dd34f3c8ff8d5854c7ce6bc0a8f0bd9cbcce16184d8698a5592c24b2a0a8293d2f9390be273c6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h844ec6bee753c035fbbe0522b48393799b37310981a203b91ff6734da0e1a8676edcef1fce7c46d9d7c993c246485e36dd477ff79313f92fe239f7887;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ef9949b4bc577d05e4a6b1aa8523d278f10b9d19ca76ebc8accd954ca8e7ac5e37d1d7d72b9651f85921c9a5943f7d543df570b39f0251f881309f4f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h432387b40c27737b3b04a62057daa7f6654d165880d4ac74b4422bda2733349cb2555595726e731ab3694f8e330157963e13b66b53567e4f42beaa020;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h861514f90e80a81f0ad5b03d725fd319503d7a93fc409b735380940d823f18ccec730fab7205a8b7f80868dfa440aa46f3734a70cd51f2288d25f7873;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5951c36b81761234106e5fbfa762db904e93ddad562bb9dfb87c3f9af942c159c066f519b0c6c8165bd69b9ba94fd78423c92669c9da2d8596ad95d8c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6717ad9a3e0ee0b959f8d822a5d28d8ee05fb925854266150951cf0f04b69e4f6162d618469c4cc28735b0de4e00ed773eb53383943b5f5bca5e8268;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he72bf8c1ad6e6082c13d04f4c0fdfa9583a6961310f56d569a521804056837bb6bb041cab5ce5f6376c8a59589604033daa4456ee774365a9de2125e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d09a9abdd69b308b7460daa010949bbba82bce412cb57a932630d071891c52841e6b70c6c509e58e190f74c6bfc0ea7064322e195861477970abb074;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e110fce20f70631f60ef34d54d2042326d5ba7ef6558a3cedc8aed968add82c3f12068a682c8807347b852622cc19e596651a5a63ebb48c529f952a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6289f0e4a4b814a360a2a4fa8066bf5bf6e1c616db2061e6c268c88b99fad249d0c3f171e56a52fb165d4227d750459ec80d4a8300bcd375f84ce39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf682f6e7b2d26f19ef105560fc0428d8cd30fbfd20a589d64b92dff372942eef2d77f80537c48a72aadebe49824ae4d0697df700c2fca45ceb43956b8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee709f0cfeff54451eb2106640d8a95bd9f730b1e1eb5153fe3c3cc91529bb554d1674953ea8ee39c02987b36392d49368a86343e79ae3d582edecac5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18a42dde17d4730b6bed4923938fc90c5cd5f0df5d09d40c8d4cb0e47d0b6a1a6c723500bc366c050fe0a217284d0e8a1746025c3e2c7224a8ea60119;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16aec037a7d9afdf8d1593dd9000078166b0d8aab56b22af269b0208c35530506cab34f42f13de2da194de90733593c54a143fea3e5b95298b49ef63e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb30fedc6a3e632a82c749969325fa7fa59b3a63fc41da8fe00863e876709de2416b8a0cc465a4ac521da93c0322e686301a409a680da7ebfa08e0a387;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdebfa1e217dceccd921efd08967676f321852fd909ced1c2e623e764a03388d3ca1800ae0ecb1eb1ed3d9dddcf29f6519dbaa579bbf555b97c9d0b55;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e658211fd5b95665fc25a7afc555fa1293e1d9514485a5c69ba0f11004cc05307b88eb9f87faaa4db36ce98fe6a8915a50df99146c41d4988b9c36d0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb296c9018c743f3fcc47d45a965c271d9a01c23ca4e61d933e5284b754baaa57195a86d31d05a35e9b73f2d1d94ab621d8fe4cb5ddb56bdf06dc5c862;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c78cdd8e06315933dcf559499edd65d88606f07e445794e80fa3ce8915ad8c1a04551cdff75bcf6ff2f02c59c9f117d4cc10979d1087459d1a31e25c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb7d8a2d71f3beb8af3ba7bc81f040a06cd7abc5cfd6ba67c98a2bf5885a9aed2b176fd65bb0022190f6ecec9ef4dfeef3c4305d959ac14148b98c61c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8bccd923a5dab495de6652e9bc4cb858eac18352daf0bca3551833c410468f63278a32f6a1636f855e5948c9f759d82f1a78e12fd8162b77b7af75639;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c986ddd0a161fbc6b3926a65345f615a8cd0d1439e262e7b0f15d4e1221effbc873c9a784263d9bb934dcb0a6095656a34234d8bcac05caa594d7bc0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde2acad799826275a60bcc8f0aee7d9a4f2fa960e2ef23331cd56f16dddec049ecd96f089d0b41f1ff6a1bd0aa9e3d5fd04ca68e583a487cfcc8f1734;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99d4622a9f067c6503695295b667618c10209a2bba574a19b58d9ac02ea3516e3678b210311da7cc2373b10e978587823534e1d806a777f908fe4776d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdee49748ae1ff2581a4d741bebf29082e86ec16a73e6980db82b030b1d85ecb670b35b3d32ec1be3bc354a0e2797e30159bb6f221b27199ffdda19b57;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38e140593236fb04da4abe5c5c55e38398177b1843f5da8a14dc2483fd5feed387ae6c52832d7f36ab440ceddd0a60b7873c85945b60a9b231f439f5c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45927b99b3dd1b36e93d5a12a61e13da9175129379451d397c028e30e03685911ce5fe118a6f80934f31e380e54b8a0551855f7e3abb82ccac5b20271;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e18144bc2dfd3a14540731fe81e320691c9fde41ecf42a367e724c81a7666e2f008d856cf6e7a23d061bdd5175b4b77ea14e46612dc3685aec3bafb9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7732048800766081f0928a5f3139e924bf8bc9bd80c14c591f9a832a5c8fe1bdaeabbd733ae7c1ab188b62e7dcaae6e53563b7b7ce39f7f09060189cf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha53d5d94463e4592d35ba8c637022162390e324163df3503a3cdefc5ad7b2219c48908f3bda21ecaacdd1f7015c52545070e7039004ca54a67c1a3439;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee548ff0bac5c6e160f975cda532734ab0afdff9fa2921e69e384093a2db7dafa97d21df98e62de2fff87f7fd1eac3658ade7df17d8aac02fbe5328c6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2e573ef69d4f163823b52b8c8fc54111d35a006cb6fc05eea283dab7314d2a535be7209cebf825cd0553039476e99a999dce8f2be26301dbf8ea95e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33f4d141615930056abc51fdb3075f48f290cae9e54c0588cf652c25076a00b0f31f00e612d50ce642d8813b22aa74b89a3efb6f138ee8c2d48114bc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h242040b9081e1ee5ad3132e6976e8705ee3cf549ccf1bd414a8bd96be32f9c9421848a96b82fbc0a881dc93c10515495ccee53aef4f8ab58378f64060;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h467360d8de0fc0fde938e3e771a8c2c02e3d70e3573d766ace03221e354e3434b9ec7423134e6f348d008d2bf8eebf10e14b4c8d7e7c5559df08d0bc3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6da6164812fead9aa41fdc1b29836e329e6820fefe8b9e858641799a0657c72cf5bef1241f34083e6b181dbd6bd870238501b943dfba1f770ef3133a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda1a961a5bd832e55658d23a96e6b1805ad4a4414a111ffa7c2d8636bafe0583505abec286e50638cdfd3238f7524403795f0d4356379bfa1075c2c70;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f2c4d21265ee4a2301266ec1908ec99662df7377f8a8b96e22ce97c8d8fd3abff9e4dc01f9ab8cc315727667ade86eb6fad120f1276c4634c2430a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8d6d7535d0fc6cdc4e784808af1c968587f04b68aeeb47e5697f2979395aa911fca7f3df3922fcef00d97165e87ead6c726776c61dda966f52192337;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbcdc9cf76634f146205f19d979191e310373ef1d639d9454220cb820abc4da13d86fd8121835309b704ad634c37291883ac116bbeeeff01ad040f48ee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he43bb51cb0eeff99ad105c580ffbc9b2ecc8207a48aff33c0b3126235d697dd3ed3c48f79eed0f7a29c1fdb87d348579be45f57d15ce17654dec65770;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb00014b3f54c975592410eada02fc59fd46a7957f69aa0387b1f80fdb5997676694234fd0b89bf5c72fb9a49676e2a106bffa6b2c9d47478c692e4df4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha185d18036c3bb4c2a004b479fd1af097ee04c12ca40c64a7ee56d9f37e5ed97af1c949aad39bbc0822eda854f6074ca760a026a5c058ac4dc573ff26;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h493364f6db26c38be99338053eb28812ec4f9439caec95e9452c42e886c37f5cfca1401052b3df2feeb473d4aeb653b7a0467d5c2372ad121e59fd1e4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5a8f0444f18d356dd1b37d9e4e8e81a585f0536d5598176348ef2ebfd051176badc45296deaf119f2266e298a375095d5edc25ca5dce5c8082207173;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf002a49ce5fc81d6c8b687e486d37b5c44ee7de71c0f477fe602ddebcadf312356b370ba2e1459dcbcb35aa3e3bb34835a942915b0527e4ad4ad6d86f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h463aed3b5112186ad3cd75c2c116bf4d4cb643c10f25ab41da72da002b5ee9f067bef514c76e90c790122fe497841b0aebdfb5dffa2115055c20d0149;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb8a7ad3037a0fbc722f4201bf9ec9b46cda1248adef002efcef6db299f5aed6f3141fdde33efee54d35f61f6f039d50ed0a724bb61f83b3e174bed28;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a4d5c5214f612b0c2d59f5fc57f634be4633279a118203aaa45feb12a8a81e0e03871cf2400c79db0c530c367fde05d006b03edbc20f062c99e20c8c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a02c1c6c94475c6bcca52d2f6447f9051974d92c2ef2e800f16f02919737b41daf7ff7decc5248f2fd7daaad18e18cba5463e6d3e43c4d165cd4568a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9e088407019d8052047e073ee481591ff88c93673396026e90a028b225e3357f25e48df2ea5e3befdc1b2fb7f1b1d67b8a13a75cbca9f612bbd8fc27;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11ade6a2dd9ca09911e617050fded4d573b43d8477f4a7891e3fcb02e24a62f43e29cd407bfd9278717b46430ce62a71d6802f7a2447265f99a21454c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h606c5cfeaf8e9ec51dc577187701092910f05bc3c3b6c06429231abd8f717186f937888f376164b4aae1aa886cbf73b5f9befb5e2d85889116af85eb9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20694ef0e14e2b9380543a87cfc9b6f34e1e1b0c7bc943ce1c96c6f9a74ce162c299a909ee8031d556759804b2828751085fdcfd3e63d26530a366ffe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7e5488a340c729d2d295fdfc3afcc1ce1eed877bbf9ee9aa7764233b10103e1d030e07c91821fce599b7d29e830026248cc43ac3f74a4339e6569245;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebac2810d1e4302cb0de6226a7d7d62f635223a013a19e4d85d2d194e96c6c73bd962f4a346382c6105f47c3607ca3afd46a0d574a0be919df2382896;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71e3d15cfe3d065c8d97d2a542642e5006612f27c7e78cb730eda63b7ec4745f49b7b1446697769cd43bd05533bc115423256e68b7f7fc34eecbe8b47;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha67734a068d9c2148ea03da1984b8ad15c9cdb6ab31509e5fca0d83429a52b9051f7174aec536856e7bfb6cca3976410c8f6aac73e6518c531002c242;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7767a65bb00b1e4f847bb11f13432ce1d8f6824e96be61bc3440ec51b2eff94b44731631709d9bfa99cf31e9874e63117a2455b4572009f49e06027b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc445e8971d5dd61bb3181490f56fdef18d33d2c59544ac3d5cac20058e7eb880e9b868dca0be49e601b4ab8f2eec77a45d0f7c70f33f3f6ed282413b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8820a3a35480df2c8800455aac6e0b6a4c787754a4fb2b954673ec92391481e91060b55910650136b4653a779ca49aad525d529f9c7882d3498e0be1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h442a19691aaee6b489670fd9b10b7d33540ae4938947efe130ada7f8ebeb049d0e704de0a16d87a2070251847cf45b182eef6d66fb366f01655ffb5bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98df022353e80419a870418a150dd962eae9cf7c70105550e2c21f67e60fe466abdaf2a119f7992c492197b62b121ce05041f4d63cfaa4a6c8770a451;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84e8f8fcae64a6ff13e4e9c29bba45e2643bd4dafcc798b58c724df4f0d59dc648e20b41bfe6d598f37db777a87a643c0b88d148bc1dce8c55e68b596;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he20ed3114d5e69ee4a30167b431753cd64e99501a17f3d56a3bf0343892409c4dfddb33dd98b1fb704cca02c4bbbcaf61fff8ff873ce4a9014497a041;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc76efc6bebbc02c453c1aba24acd7f181d94adbace91c01e0de265f0e6d143f22b501fd250e3523cd172be7e1a19e59ea68eacf72b3ceb627a7a6aa86;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a26660d731d8ca8a806c2baeb876c3593b03827cd3fad90c1c9960eb6c0c55b19a77e8564c361668aa7554acd3d9f77874fd942e305db8f86c38e3d8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e934708d39dcd36731b9e9714e970ec156970b4e3f1a991d5f8bcb55915c34b1f1d9fd73ec618e637af2b00f8f869a75ac44b2f3348a55fde649ade2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h670f0ca9257cd8a312d483214ba59e9617ae3cc7b8390ad6b5e8a906f8fd6256805623e639a59a1ebc04ec8a035db3a38ddfe8b139f7d7c10369a792a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd3e5068f3b6b1ab1144287554b3a7b767cf4c82f55857b5bd37c75f76da80355a00b8b2c6df3f1e682830b7db3046a8ac2c8c0f261462e6f33c128f5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h980a138fdb748cc4343b2a179dc0509c02369df6764155d8553083577ea84c3a09dba5c0119f1697fcdde99069f4507db80c418a237bfb63996117910;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d171014a42bbbdb0fa1317abc5d3a79e8c7d99c066860b7021b3f1edc602fc71d638dec01f16683cd9b4ba04de23311a95b256cd32e3edb86d008b10;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8f87b89968d11ec7486617c06c59f4967cd7a486c9ed3f20dc04ef00d40ef8291a90f662ff7f1064a3f2481eff6958535eec45b031090bea825633d0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34d043d2fb8479c6f6c0e1dcc136ebbbd7fed8c79cba95a9df13c7e5ed7a32f56ae0b51168c46c1fe56277e85ab2afb04fa8acae5638657c44202c9f1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c57c9d270feec1babef49a210d2dafd69a44689aa190c5b4ace77e885e60cde6466e4c5fb5d306d42e49d9a873a63d342621ea8baaccd4e304757fa7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44ba9e7ee4d7703646f1a18776b18f097a4fcb5616e595b3b80940c477426e750cfd6184afd8059a30ddad591fbfe07c5f516c733cc261f2e737cfecf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb58bff1375003bc9c976987828536581f9cbe819a19adc0819f195e80fbde268b8bbfa2495293ba257acc20777f0aef6fdf5d45f2b06894eb25dd24b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18516c233ce5022fbdc3e6454e4067c963c9f6e84aa2f13d2a09baa367b7e009d4a4ec01c96b706da5902224b93fdbe34def437a003819a2415c53a42;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3097d3fd7ee2b8e3b6b7584f911eafae70895a25232df62f4affe0a86a780c48a08c0ad0f26d52e0f39386eb354079374af1fd4998306392acbd006af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd98e2a246d1bec97558b7e86e5b95b595b9795790ccea0e043cd2494d4e500ac1942eecdd3fb7106988e5c82c639caa95c932e409fd0791551664c2f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91b6a1c156ebd2022d807b38b2955bd260b6181aaf82971100448a9f5059872d767761aaa7f298f785660c672281fe340d94863d2cd4c99c9c91eba33;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd86bed217bf68076744ed774318827d5892f9d0c6f5ee80cf7ff0e0a2d246e7aff41f289bdb3c808609af5cf1cf82758c1ff4967558d41d5bac75f9f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11572468039c3a8515f1a0be96ac6e46e814f6d94bab74e72e654a0badae60503f213b90fe0e8b28772b461240cb5cc73ddee4c60fc6cf333e526f709;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f7fff32ce33120a61b168a6c1a708e407e8a4a74bb18e45fb0f98947a5424b5edb8e9add24942da1f30501f6cf9d32f31b1cfc7991889c68bf365407;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed498719efd90d658796bf1b28c1cc08da033503f30b31ceed6552aac7b45f72782e3a2c5af471a1398aaeee82a810e255f52ab1b177fd979ca3bc989;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5149ea9ae19dc3e5f0975e257d07ea41ec10d3b122eb30715a6cd8b9e0475d5dc5cb9735fa2ca2c94c19b2a82bd2f1ce4c1db811e66915a1968fa0e6f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf51528659e83b306b9f576fa11a32a91509cc14e4395c0b9276b0ec324c99ea99117417e376741ded6fdba8535e254660e429cbb9c992eed4000e5954;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h747845d55f06785d5f5075fb697de27fa3183d8cd4ead570950ce5ca75e6109dbd49a37e938759850f15310a0f0540d9ed1a38caa824d81bd79ea2a7d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4282a515b9cebca0ecdfc5158c89a313300585077919a3934b494d85fe29d79695a0a777ac9476e461e9afa13ad32e2f0d064ab6c3db104f33834932b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6831b5baa8783b3dfd83be0944f137a0d2fb14394b2b2fed47a31248cb2d43bc6af7e0f5aa8a4cb601d96361bc2f5c302b4b50f572e01a267413cfe7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h654ccd26cfc24d7f034fec94561c1d546f3c8c0777013ec69cde074617d03c6c3e1d21ce1a51da9b7c6279ebf42cc7f14d20c97a798238ce2493155b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18baaf85fcfb3abf46570e3ccf673829b9c4c1c77309e2d51d21a39a63729c0e40702b4b19b28a006c3949b114ce09920a733d6225e52b1e64c8adeca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fd2b4d13aec59ac9b47fc7903e9526c07a15ed020a2cd7b02db8086071c1646466abe91a23dab7ef9cc58df996e0d48af127b5fccc5632a8b2f90143;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2d58667f5c82d35573a19432031167013ae4d0429dbdb09637350b70a77844fa32867a25d686b76c693e5a63ebc623811e9c5994b6defd676e868bfe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6892fc34f1f97513861e6497846330ab3a8ac628882188408a97a6f92ff4586c39e9f12a03f077750aa8dc6023293aeb87101e8147d363dbe18282e08;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h335878af11b003c94712ea922e5fe2d5daba5747528b4fc1e93a50fb32219936f4140deaff3406eceff785b9194d74a70aceb091ac259262ab6a4c553;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8adeec4370ee6e13811f91d89bfd2481a280db82039ecfe56a1126631839dd1c411c3cb3d89ec0fc89f2c77391cfc13e4f7235afc4188f76c3974a2a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbab24c49bb7c4919aab275538de4cd72eac7363187d6c2b861cd41a82fd7b91101ba2b06f4bf61ec4069ed553d53e28164371eb5d6d7059cc8e0629c9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5a6d0ca5369ea32e87244257d9b107f77e71885dead744b345becc44a7e6e83c6619ab56629eb7fb1b80dc7df356e74478dc45158a2c0bda228508096;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he83f8df6bf181a951caa424e46a5eb1a32cb7c57211c299021d42bfec6daedc91ca60209e0d47a0394e4b007490d16b4b8c07aba258043da765cec04f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19944af3778e56a2a189b2f37bda4c9c3737d9dcab7000e209de1bfc54ad35b14b994c2f835af29c786c3e9dd522b0b7d6749cabab8492c240fbf0ca1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha428751610f49402b2727d5e8920ccdf4623381d807c7d7e0a7ae0ee26cda2394b866e6ad04a5e5da7b3dc65a5ba940db7326e25113a1345a18514831;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d3786ed4861d54737b87504b88cdfc9fe3c52e69269ca465bba4827ccb3a2d94f45e4232644e9c2ea80c4d1730e7dc79705b8cc65eeb55b0a8a669ca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cc425fedc3dee3a58e597c9497c37ac40591b222b004071d75ca9b1904487df2711332c5a6c6c7c11e148384447ac78b048e96b883dd9f3f49c988d6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5582a419ea69e7e3a8991316bcd840b9c9034a37978b4d039c2cc75cb43b08bc0ac20a0908f4ce8b1c1aca595aa3dccf6f5c7b902a6f7d2c8b321e9af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0937b37495d658d355adbcc7f27b2e0c8bf8c888852333fe446dcda26c609b50ef92dde0e023251329f2fdcb1f4d4447b6ff33a37f0827093cfe04f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81000d20d60b4dbbab8560421778a14e7c05d3dc5b96c380ae989e7293dc3debed857f64d607260d62d58f5b94cde22e9b0fb7e724b145e83d853c6a1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb5d75d9014d4cd952ae9c08a0beec4ed7a657de45c6efd4cdcf1e768b9cc2c72f32bb2342ac2153158476f4e75ad87c80019566dd547f69004b9930b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbb4dfa9d26b73f734288d5aedf4276ad3a7b1eb4820eb0858091dfe8f9a89fe5556803de80708684bd6ac791f8ef31767ff434c80db140544309fe18;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb070f60eb98abf9e892d00575d42bc0b09b918edcc85297c5c4cec3ceecf340170aaae4e83121c15bb10feb4f1cfd00d7839606daeacbf57783975913;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6871479c894dc05d4a23be47a1a067a658b51878f08879b96d6e59abef667ad656d5c1001fb814ca201bfc103141ce736cdb75ead3425bf4c335bff7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3a833748ecca74b27979b8b8dea22f63da1841e6feab2b0a971218c0aabc3c8a1e28b0b0d6113c604e9e6e2235625a6ee6ab245d726401deddd7b2c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h888dae7d9cfea64c1e16346bdc1b9ab16a52d6e9619ce59cd3147f373afeb59fc27248bbe41a40e10303a8a9c9c31b50a71314e6d799d4bbaa2e6a712;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea5226bf5f797929adc4b14b27bdee02a51d2f2b730f0da3209dda36d641ae5de4b8081b9f5f1b7bd2d0445f305a109e264a31af7a6d273385a098c57;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfeb14e8d694435182cef3634bc4cb530aa31ff0db91e416ff876107a2d3396ac66404892433f2e8a80b15b99c345bbdd5637a7781509e44caa61ba88a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1c5be554b36d03817abca197d5f46a91139b35b5f54f05ac3e687d7ad1189fedc51e554352a1cb134b65a7920c03b0f32c2fcda34de563050738054c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1dada1d177d3302f4fd5b8583d7c6a035116445b385f335b13c87d6d3e13e59a023f4dadc5ed7dc286686cbe3790ee1b457474ba85cdb4c5037160263;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b25ae939545822f7db0328a784aa1519e30f5f2474b0bad0bf516df24cf12357c895412a0b3a637a280a4499774eb3ca2f43d68aff1faca0920290ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h825a305dbb48164ca7c64646b69f246eef7c76d5be6a8adf1a30bb1d07f3fbf0f2a007f2dac753eed1a5f3ee69bc9c6784adfa3f453f9a0a513db86a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2516a51795b2d2bc8d8d135f5ddd9642a75bd92de1a892680da6da9aafede558564e35b29b4b05dae0a48b9b3049a0c15e7302b47a74baabfa9999455;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6b00ab831589f6402160d2bee517f03ebf4f9341c0ad282d3e686e092808caae5fc2740ab8c60327c34b0b0712be32aa990ccb48a729e31551d10c3b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc459b6367c7a76fbc8b596fd9953fb77ca9365e8bdbda22fbd4b4c4e88284a2bb8a4d2f92da34e2b6fc0674db28e1583ba860524bad0eebce5d106887;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e2f1656cf3b73a9f782f3bed6c94e4d53738906cca162931e5c12956db229a4fe2c113c44033bf54abd053dec6b1669130f163b2d22295276c4adf46;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7278b9da24dd59abcd5166200c33b48b74b24de6abd2d66e4633e67f2315979bd1482a30791dcff4718c48c41c3e6b5103e8eeb91929ae8a1716d0ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7eb2fd0be82e1d7143ad5e7f19115d1c103322609bc4d8a3d085ca6cb672c7488dba8f311c765d043d0cde633bcdf7c95dc142f77dea9e73662cb913f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d6af7465576070e6bf8e7bb11990fafeb7fb6ab43c068944ae9547dda0cf026ca1d22bbd98b247971dc87e30e86e9fcca57736436984a71e0c9922a1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6845e5b187563fc84958897381c7f6ac9b4e000b0c6ec91af252b7d3e769c627052bd267e19a7b74ce04e2a251a23ee582d4159334b90eb136895448;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9372fdb80f17c360661e110fa63c92b1eea7f3745feee147bae78bbdb14538ae72723926b8f89cc34f25958296cd63aa9e317430a70b85e83f7f0e7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43291bc7bd4f2f917fa42761af9d0e9ce747a57323fd97b9140f58ee43df3846fc49dfa2369cdfc9d0c6790ef7b524e03720bfd33065aa36ab5d9b328;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4dc135fcc5f14b493ebeb070457fe38838ae70934b977724f78eb43ba6594179a25001ec58513029de09fe5fcde3a9347670a2c0dbc2df035ec833a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h895d97f30da3692606ba8b4b2f2da5a45770d907cd8d5f1a37021da24711caf2b2d1d26461417174419a8216b720dc820f294b746eaa614eeea51fff1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf34dbb12b066390bef8f430c6300414b2afe272fb228879c20c3185ccba6c56e73c73fa7d033bfd270ef456cdc4c21cfba9b804d652f72644d2d5746;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4902b7c005cffb1c00e49d79536ea927ac0040e808f33fe50ab09e0937c4e2b5a0159006c949f441aaf57710526c0ad13c3aeb8331b9d6826fe55e01e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h217e5bfee6e03c92c691cf0e947eeefd06a95f9e3fc3ac84dea46e4bca40ce001b843048a7baf4b41a389387d556522eb9eb56b4443402e775dfd4238;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha431a3b910ee449e96767bf351d6148550b1fe99777d60dad6719be441715cd6823ba5afecf66bf876a5385334d0a9d3095021374de9199668a8a9efe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf40a79c676d4a0c128899f80bd22d9e1b66ee8dfe500d0869787103827229c77ac25fd08f0e49a491d908442ff6746081f030e5057737565844faf15;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcfe783046c53a40c452fd7a577bafd93367ebd46ecce13edd88b59e3782775e4bd200b8f925964d311e63c4ef57a1e349445d7faed55bf96e2664da05;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb82df892e43fa0e90c88674739d2a78dd6b614ba7d7a530f361251529be5e9e487af7b510c4b830bae1e455d5dbffab1270e6af7c02a2d66681ad05d6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfae39cfd0fcda4aa0c8289123a69bb1622e1f0854a5f9e2df31a9bdee3108ec1ce2cf87458a913975b782b881b67ebe803093601f80459b67a15ad2f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf795d4fe38d3831ba398c11dbccd970bec7cb497b713c509675b5d2bb9ed26b26b29920084b437a9b1e8be59749ac08272c9dff699b674e056205d45;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf82b06e26feca76b8a734061bd4b9423aacf888d6ca32697b3a0a80d994c2a8a52f2014aedff45974f17f856e0bf9271de89ce375f3ffcd52e14ef44;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b86fad1e3b63708bf1a9286f00eb23d27a39869274006421eb33eae9121e5edc19d5036c4e49cbbfc7280fa7d53cdc90b3c9da0c7de2514185ac4a3a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha01440f49b32ca096df7361083b322c32d821bcc964570811d3e950fdf24131e10356a316301a6906fccb3a3e8183ae0337c8503d7fdd7e77242801e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef1fb78c39ceb46b4260cfc5bca1a17bc80f22f9b7d63c1fbe64891fcea1770d6e50251f67a2d71dfb294e5b907a26c327217afda1652888cf2c674ae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b8ec4a3c4b3db36d64da447ce91bb7af03a13fcaa96aa59192d7aa26590a6b7cd306544170141cb48bc667fa98637164cb64b76606f4e724a5d665da;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4188e495a1cd10387d0c97eef943bca37258826325301dd08aedb097e15976ca80e16b82cf641d3f1a0c1bfce0b895487563ec0249794eb6627f228e9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h853a2c25d1afd12c3d890268e7677c8fe1d07b715ec7cd028b4fabb193e6f66db1beb60930207b7b751fa77141c350591523dff0180700ae7946c7be7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1adc4540715da6290be13da3367f9598e2a11df5ab48339d48bbe8260522b7a6b47e615d4d419af30762337827d0b204f90f2743b5220ba41033c5a32;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb80a5889416e46ed72ef03bcf23e25eb7f73db1f6e3b5e63a1909a7ac55d458752fefa79fee9068e7391d5af328174fe1a46d5b2ddfbed6b91f49ac1c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d3e64d1d6a2557e2f95cd565531b4683876b5665f6a4284d317346283132efe24953056f29b70ae831ae06be7fc36a10f7d6f179e2e66c77b0a35bac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48ef8c83297014c1533962473cc51db1884ad43b64ac528bf6d8c515603619887a10b46c661516d0643b9e3d32474ed9941736d56a16461d83da1d5e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47ff83ea5d8e03c8e4acea05d51a1509ebbb7390696a6de5fac43c0585d7a0ce709c3944e732431ff5fd19f7f9e1b7e517f12e3528b3300d860b078eb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd77ac3a465861f7c862257a5e2c7610fb5e6ea7691962c9082d5f58b44f82fce5ff8bfc591ab6a987b3bf6a41303e2b7f2406e53b92a280942ab11f74;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f32b4aac8409122a37f6bffd1962d2c7a72cf1c8d85577402785d0d4f9280e832d962fa455bd7a39cc41974c072391b393b067f2fbb35a895fe78d37;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd07b28bccb91c502079704c4dd32cfa02b702abef517e03a9d204b38694381dc68cdcb7f7890ae422fb00a2b7935404102eddc12653cd3fcc672cb92c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6593f8704e52336a77fcda8381f6be57cd1ed3135605f3f815214cd543bbb9b30499c2c32e2cc034e19fe4c22d2c6e427ccb1ba4f1f1d1f1674ebeaab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15ab9c21cc334dea0ff4bc1e58b33dc4057029334d1c6e4b7a6dc6738af694f012968bde2f47d26eea1dbfee5a456f3f7c436a6da4b90bc403bafc5e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h828c704eebef7e9c440fc5c5884c99108c7169b8d4ef667c592ec15b6073596dc4eb0302c64cf0f4f51dcc198016bdd3b81be2426c08f355dcc168185;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57d00dd32f76c8eff7f7b869f519ee967e09330602b1cd596a2ebd54c4c9685ffad3476e8349c813c9dc799311286bd36a4fedfbf8997e77fddb67520;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76c08140ff888759439bd5c53b55f2e1293c1d3b55fd478891140db6a682e7b05a6cf0774bd1001af871777ba67c29c607db8ea88a62bba55fcdf7730;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65c986ef69ab327cf0708515e582f50129a4bf72ad9b445f803157753d8aef774e0b8b22e37832b391f2d588b763c59f44ca05b04b65709730b94c4b2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h128334770cbc57a7ea3637f3a5812f898eaddb53c3763fc661823af53a84e85b6405e580a4140cfd8d345e037eea92bfb9eb83daf96eb45483ecabf11;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha701ebc12e3fb87e0894c8d43a5027f24e83cec999c750d9dcc9b91f135d93a4b1fbe80e49ae016159e917e8d8ac6710d18c739eae30984ba8bf96d5e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e2f53936b2a8c6e23d0bc75e688f6365a930b00bbc08c1ef342ad7773b57e694bd20b1813a279c30fa28c85c7e6cc87544e5997a4c795c04902a2f35;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6313d3eb7ad8f3984a96d938f66e7646c502e87b6952ea0438e9ec25a24330c441aca4a0a8ef4c07b7d550d2cc974cf073a82d1ac3c39e68946194b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc867585f3ca62d5edf37b877ddc7edecf61755d2ee64edfbf22666b83659cd436441545e8ef091f58653795e732493fb37cd0309762aec11d14d1589;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed9e69a7bc04cb13a2134d6e41266b11c5bfd64a6c008552477e776d2d7d1fa1f41c193823a96cc5ee08d7f91777b713d462d5a3d2ef5cc95f80fe597;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8f169c2be4baa45ce77c622ccdbab0a0408f63d41b7d835ea0f6bbb26c9a2bf64191693dc81c84f533fc5c52c6fefb9272890ecca46ee13b3a1716e9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee6b719c0161da694f00dd06329350fb560769950ed4fc123b61d17d3daa18985b735699c55af1b9994fd06eba9671936153a153abe7124a4d99c3a02;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd8d228664a94cdb50295def45142fd3378d83be229251c01096ce7864e136ee84ea0a7064c19a68948cc3a363b8a1bb255798c03ea7b19fb49cba94e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h963a5f5f9fde2a330553a89e80694d6db5adef2efd65b7fd37f37d7605ce00057c064861e440cce0bffcd5319dbe9c41c6cb742ad63f8bb78794abd74;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c973bf53d881828d2271686fbd4f3a9f36a653e51d64ca74a0837abe458f19cdd8fe1ffa29ad1ee6b6fd841546b51ec169dd8610f59ca072ba3f15e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf0a4c9998ef2b5ac9021a6d2b50ed3c7656febfd818854f77d3da214bd62a5b0f09c8d4907b9469f7beeddc9771644e95628feca51e2d5bf7dd98543;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a5ccd95a0887f549abed1a77a10d692b67db59818f1794d46611024a9c01aee9ad7b21e817ee53dc4cb2e80f2f1ea7754f8da3b1992472848b27897;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf16b702cb000cf4ea331480663dc26b9d709e6b3c94481dc469b355ba9f4d2395b1c2f50215c900877ee610dba7ab3851c2f3813a814762b6c80b1a39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1327f4909a6722d9c70672a1517b02f76b805803d7d829e6e06d602cfcbd299bc9420bbb0cbabf48a93f972c38b4414e1e9a1836bf37177b8bc3ff3c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h976e5744b33fdcddb012a2678593dbd7910e6efb49db1eafbbdd3f8a2bb6775bdb0710256942b323506aa155ca3a02e9223f6f675aced780a40d117fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd1864d4ac58008a5cadea62b315dc7d36cfcbbf361a9a09b08f8a1a74366ce4ebd33f2047b77c3bd72ccbcfad6c15a376cbbe9db7fd7c0e4f7cddf9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6304be0a29dfd78da9ce3cee134f9259218dcd20cbb836700b0ee0485c129c343ab3cbe035b8c966fecaed8217a20f120fa7b3472dfb0bc1858f1812e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40ba85846f2c7103455c411be65c7b0005b5449777073e8442168951652b60459b46dfa33e21fd3c0b9c13a298c3daab3b81bd845a4dd252f55cca42d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66dd0f52f69f910d68f2683c490c3ef36085f335d0269045cda060096b1ac4a1f2ec8a7f8310767cd09e70042e492b5e183caf5800074128004784831;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9a4acb44a1940c2485f6a15b52fd00ca74f3b77a8347102513b94e6987bb7ed5506a482b2e8d7378687b555178bc6a433178d5120c6734cda5d272db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b8055bfc2f07f3211af293a02b9aa1cfbcfc26e03a3d639b401e538fdf9228ac93a5915c4d8c4583ebda202d7c82c811715923ba19485a74323b5e6a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a56a2a29b8dad91ab45178ef23d829b20102847737555bd8a06dfdd6569e34c6d378022b1c3bc39a1af1df962769945b26b2da68d37230607985947a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2997d7e4caf4b00ce4050bd037fd1179d1396f4a5d6ff89f1f625ba82b080b017aaaa2a3ac5f9719b5c6960e59d7aaa3a0b3ccd45f83956d8bbeba603;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee939c7910a40e47290d73fe580c2a3229e36f8e47709b0b027f01db67691b4ffa83ff6139de1e966033b0258e9f36bba6ef9342125d9a9d835eba7f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4910f31474d957d8058a4557d5c59c7aecb513b36f8eb0284697419dff737bfb6fab837f821e5ca9af4ae2d6100a2efef292fbc6b0d4e12d5b97aa4d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e8f41c475396eebf355c0c9286548e3f2cb5f66d9dc63e8542d9ec9ede0e780e602ae47cc8c81380297c3a3f4d63b1885a0de6cd38d7e528e3273249;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb51246cab613595ad1c7e2682e3a4215b60281c573e6f8588fd13301ce40ef63b876f03e2ff5a025246470efad9c9e1c3abc60016d8eddc56a228d48;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7805b9f5952f6370fe66e47cf422b3572fb283c8390ec4b0fd4d12f1fa6bb7ec299635d749de5f9516462062310e1b4cb259b9efc59ba259879be6682;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7cca4ab6d42ab9c9b2663fe1cdc710ca26028a21f15d0bd7ebea400bbe05eaa1626d284f961be09cf43a2958c548abad22bb8735d1fdd791bbb744865;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8097eb56ab7a9580a26d804a252b56c5cc9ab0697df27b39abb9d993f4c4c54abf9e15f9fcb584e1b6d69fc85d9788050dbb39f17d9f2697ef81dd30c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h387aaa5d2563c4038249bca3cf29b36ec28bb2dc8b0b4451a6baaa020c2cb1917d96f018bff9b06f7847602b5695370044572aedf6418631db2224871;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h810529569e2e5af38b2accec14f63f30049b7b865b9ee9d8edfc8363c5af6591dca53cd877077a954d59aa77d6ff0c8b9a0e85b1d0dc4e5d0eec2ed27;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacfbf1408c57cda5046c4203bab445a4d2d7f113a42d558f38cef601f72aa7fc37ebe9d6e28bdcc7a739bdb4fff037b3882ae11f25f92619c3d469f03;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a90d0942025465cd359a79f87b942fdbce3443a3b6d31da1bab363319e81bde6132a7dc95ecb04434e1a3d7a10297a8f9b0e00022dc4b9338a7ebc55;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87ed4f530c174d021240e7b7617897427fbcd1173c86db70739618ab9e679c2b79d3f00fba91a141223b6f0926f0306aa173e94ab67f52d26435c0aee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h278e784f8c65f2e05f5dc001242909ec7531dad31743bf39548951be90a8819b86a99fc2f939bb53170440a7004e4669fc38d64c94459694c1b9665ab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6316914bfdb24cdf9fc8d62e4858c79292f95c9069004cf620de24575399f78b583716d69bc6f29fb119e0ed197c02c22d8895cec7984e0c5577d442;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90568e11b9a0232fed4ae1cbda8db1429d2e8bc01c052f93ea11ab33c3ebcbb6b87174354c1aa5ee5985c5b3403dc0f3ab548b031a220a75d218d1dee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32e2b2df6d54967903a037167c1b0c6b244156290f26f48d466705a680e0d5f75cac8b68d3e1ba2b38e6a45f519b6471af7e5c1c11157efa597352fc0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf689dbbcb0841a41cd996f159513ec5086aea37863cb0b28c9cdd91bcbe2a70bca7329414082af3da0363cf7eee1fa663f8b1a2b24f4db31d07fae41c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd4d2a448dc1fb708160b63210621ca83cb3bc81717bf445f58eecb8dacdd2956c696a7b55c4b56ad3ae7634d9285cb141cc513200e45e05e5d1f7e31;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf33471dec1f2f8429f6c66b7bf2271eedb06f03c2a267c12b28c34345f8e7b1114df92b0e1e13e863084fec37c571c816974cb9964cf1f239445daf8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b4f1f8545a3ff638de26ed12f709e44c2479278882bce6733acb859d1398a74ad2d688b79cf688be774be3ec65b61b3501bb941ed19929c38f5688e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c58573be938578101422646bc50fea879a9ba98420c86245b46128338e40205c8960c991811375112401fc9f9572bae4ab7604ad781717e35759442f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54f2a2e7f83045852b4245cc0a42c1c341e7e4b3830cf3e18d26c7c1df8e35423f19fc96ff3595ca0d94dddab1202973c824c87809bc31c43bca95fbe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38a745d28517e440f6ac22eaf7189da9aa6a214ea21f41601e70dbc82242f37d02bc6e5fef4dca70c4edf16acba97e37dc8875fea70e9b7beff3a200f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3ac3a32966715e45d807e66164212ecda18c8c624c3d173fbf165b1d00966563df0efd621ac8643f37b94b51769a6e1cca0270be79157108836b1b35;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4490dca5381853f9a5d70050cf22afa2ce404fd70cc1fd622c6b4052edf12671423d9a444aed568e7c3e567f9938208e13dc0e7762da567a4e662fe13;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ff7d06861dd09ee201f42f8e3979ed520fc9dfa1b36f1e3cb2e226935852cd838c12eaaaaa61fbee3a544573d5d40ab721243ed7333b9ca782c75446;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3f853cbc9f774ff3a966ab97b9d3ac74eb6405ddcadcf62830add1175834cb32a8b6b07bf61bc6d4669523e7cd1b69ac9440beab5baa57152c90cb3d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54017f1d9c5db78363be4a8f25e1043f64bdac58fc685fc275a50de6826f003de9d1eaa02833a6696597c62b8390e507dd7dcd4e3dfc71182c35d6388;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59c16b5d28bf712f29d17a230e4ebb6284bbaa97decf79d2e06c367ca9b1f7102083be70b9392d8297407d8437acd09273c10cbdee199e900e4857a7d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf83b907d23fd5e063f55638f258c985ae5ea9ceffb6013d552577d2d7204f049c95149d9237fd1dd7eb13a80c0e07c2fdb8a067d41cd0cec52a597d64;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h850c22f3b8a5299fb07448b67c56cc8e4d3fbb6d9d01a622bf0354a0b0a58d5f97bea183240a31fd778cdb5a7e4d2f1f381fe1c34e8854d060c0ac985;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c12fc727b49c6768bedb537240d917cf4418da70ece66b01d72bfd7fccf838c458e3a9c2cbd9b52f591fc150a096e5596c77c054c722d4248c972f72;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h159502f5291ac67d02942c980e8d3c996b3d53de0a34ce91b1151c9d65a2c22055d46fae97747ac8643a488b7a07db31c2bcc76ced372e64a7c276778;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h629600a04d6e8c72a0129e35b46171cd237420174b16855f604220da8ceda89f63111c96ecc1582240280bf255236385528699c06bc4c8eab74db8e61;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54448cebf087dbf817a53495535ad7c5bd15bbba8b71daddff230476972d02be6714c9c12f8002bcb1c16fe76f1d0148c0ab54e5d68ee4aa3e18c4a81;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f697b2b96afaa19360de7c9c70d0455a1f2e9e85073d5384e62832ec7114a5921840b8828cde5ac45bb40f2e5250616ba43687690ee8e4d99ab93658;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5d9c58dc7b3e94457c3a762b7172ba3b1ed9619b3cac705c2baaa15e65da21a135990e8800c50a1c9f0be70adc7a9ec877ec148d4b10c94bd5d41c50;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h595c2093cdb81e67169047a0310fcad83a2b8e9574df110cc153d5ebbf374bc5bd9da29ae37fb3252f360fae90191835225677e313324e7fa6f4e4e0a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c539b4823330ad474e64c2c87ef159b50f3d546471ac96f227510ca18ece2edaf17c40021b5213a94c9c1f2f1c7b1923fadc62663a01ca809d6c0c9f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4023daffa2b3b4a064a82ac087d43b8b0f13446792a1fc00079ce3b06ac3a104e7f92ac77e96e583b715394250bb467d5fa98c094bb1cd550ffb5905;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40bd015e5d1446565c6a4a9db03f690c8aafddcf80c84949dc604e19784ce83a1a683d2b654a02211fd2f6350c71d1cf955567faa0de52c6036633aa6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a03fd317c8f8ec50af8755fbdb47be05fa1a24a7373841a629e22e53c87508233c8ebbf1e65a874cc0b2c8b5ab17cebe8924ab875606f59958c895a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b3484f2872b820036fea37174bfcf79ca1ef314d153f897c496c9013ed13399aebf69ee5e9d96bc7e1ffa43573689e85dd497a3a1c2ecbfd68ed3fae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b98ce5789e7b26ad68145d0e5d6b3cda1479a6d34ff7c8562758cb58aad123bfec2a42ad7411ad7df157bc951f5b851202bd65f15d963bf41308b097;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h261f3bfc26b414df458eb39e43839b3536e1f048502d3343591a8d9579ae3c3d40425bcbdf37c364802495de3d25d3340a57faa27be2f052357bff6d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2deb1090a6ad50a0bb17e9b304ec34a3d9d71dced1d1822d0b2e0aad8be89244e7bd56d36f6eb2d536a8d4ebe26c91e3812d825acc149f4a7ab9ebca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c49e808ee962a70e84c01de58799060eae140ca0bf6475c4b0fb15e0bee653967e35d47e5c7e180062db198c0072d0b5b2f994d01a2d47047d8a0c6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hceee70bf60fc44f2fe046acddfa7eb1d28bd94da16343ca118a251680be1d5685f248a9ff516cee07017fe7ef1c6629174d4ebcd2efe53b43ce9ff8c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83702cf765ff48416e8ae137e9087594b87c475a6a4894602ad7797dd9555a7174a4d8d82fb938cb977b557ed46cfc3145f31c9ff871b086a2dc220e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hadb18f037b7242ac5b8d3500d22db7e06fb9a0536393565ec9853b42ac324b0f69449269e5ee07c8ba208dbae583ccb31f5bc3c9434a9832459686c3c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd64ed15046e2f7ddd8a61d0cf61c4b92f0e201bd048fc63299acd9307c1fdc382f5a78d460a216ab14f3432bd1361e8b0bb5d0920d1e17b73d95c8f70;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2281f20e8fb44c9ad7f6e5cbadb9b86e6132ea76c42ce055a31169f333b456bde34c32931ebccd3fedb33c8efed3dec91763893891003cc4dcf3e0958;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b7a4412b075d5aa5fc7afd7ad08a7df6eb58975f55fbbd98d416338fc49609dceb075b15834ff77b951bae7c1be1e9324e50f6d45208ad870d76daa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc888b4a3586cdf3cd00bbb4b1f26d2294900f72de9aef8ad7a4dc26d9656e13cb2e4204ede96286ba678bc28c2d36dffe0fe82366c651d1d255396b5f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27e50473fedfd434a36d8fa5ac9097433a5d0a6d9a6ba65d582c483c2690c4d7d7747400d4074241bcff2ac29032a9536d3e233b5400688b109d367a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2976f6cfff176a1d90cc182c79c42580acb8069d41c9e352cae0c71e12bfc1cd75665d6d6d6ead90719f9f36df937a03a87a7cd9229ed51183161b15;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9940dd6dc9f48af54640fca55be70900545c026c3cd00962e6bb7e79995692372d84e985da89e1de82c5b9a4b5fa0805409fa121b23c0ca7d0e80e0e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb392710351a17384b9d023850a7cbb2afa6372ee88942fd49918b8857ed80abeba4d25f3cd8cb61a51681108e65b1a0327dba0d99df9dff711fe8a15a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e68b8e19200915f1688b6a0e3280c204d10d3bbff2ae82fcc1d59b033571cba5d837e8782b1aa9ff3dedbe2931a433d316f3eb716952270b4dea82e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h618dd8a8d2a35c465ccf5a02bf763b680539fb9a6839bbc2e5ea3cb27957c7cedb6f9d44b98f8a50afdd40d948e678f22f3ac8dce483c9a9cd4667546;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38c0bda48a9c85a11042edc2851494da4fbc3e0afc0dc18b46a4fcef83aa3a1395d9594e61dff5027cd1f6320ba34a697a0d610c18e695326b6f434b7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e02e71e54ba979d8ab4b1ac64b8fc924b4d6851c03638be61ac78266ca805ad65b89ee7439175b732bd3d5ea7dcca7e38a44b3e27ce50b155f410301;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33ff424ea0b7b750f4ac94adbe1c9d8798951f73c32332d3556dd81847b55c79b58ababdfe76d5a013c9e35a56abfb3245f223e75ec13c4ab90501600;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h869955f907f43a75f633d1c8704ea25aac880dcc0aecf2f37d4eee7487f3c9ef109df1b7649dc7e59237e7ef3df0f33692de34d5136e79dc7c7e445d1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6770f31da36ca6a0a3c40eced14d8e2e6f8bff3202e11744823ce1413a0e70de583b35c378e60b783c12ffd2c3b17b6dd53e61cfab0a4a028a4d909d9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha993fece26dfb7c7bed04d84edfc73400d744ac88001b96b270fbb2e2b9d3ab539a7019fece7e8466a237f1aa7e1c60cb8672edd975adf30294177ca3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14405f8ab5323f894159341a213454663da15ebea24ce44e80bddeb73c8247fe4e54a1183d1a650f8b78a2e5ba96ee2743bbcccd95b6fe4a1a4abb083;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e11acb509f38a6fe28d255869027f1c33f1b573ac6e34ef1b0021bfbdcf5b9d7297e1c89ea772f859cdd277b4f106900df4665beb831ac6871978aad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88dd321288bdc8bf029ab64674c792fbf4ef25645333c529869c4449b9ae34d08bf6fc0918b8badc011a7f62fe22d399d66b9eb5a60616aeed1753fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4037955013622811e1333d68240e2ddfb1e3006c2a8fd8fd99235c0aa4ff83d479b5c5c1b59d38d894c492c322023edcd725d6f5d9506cca9295ec907;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb5df8734a5357589db9d68ddfc56fc7af21d62d54509d3b792b47f8040a57670378141f9c6c796053f58306f9370654dd8932b971b1d2e460e23eba8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac57da819d23184b9094522b0da3e0c9d9a8aa642a0801869a4203403c7b2201457a851262310ee13a08ea9827a146e0d782783242cea2f25fbaac949;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d4daa77e2fb339d30f06934c319383f04843cdca54bfe50ec3d896fa4820c4c9f5da318c5d697e0094e378cc85dd75ad76e8117d55d2b10f9a03aad9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65fc1448dd8d6a7ada43387a50274a555430eb98db83f763e3d03c55816618e4eee0ef39b54169608e90a292963a0aab93b2ed44376bf3892b5726943;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h545cc86b15bd6ba4fdfaf67344b45475fe20a3d119f59628cde793e881df46e40eae0aeaa3bf0dd4bf109b9b16c0a2700c32347020b8ea28f4d542707;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f93a93127e3114d4bf1abc75c9066d94100f4eda719e334b6e25d5c3baf288372971fca28a71ffc7c47d58c1938d9ecaaf21a7a05f1b8a92ad4ed246;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1578b0de878cc8a0aeeb8bdf5d60c2fa927a4b29c4d236469606fb825d81c71dce76f4c474fc5264e6f9d6ee2bf61594f1186faed56e1177e9d2af41c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8561cec9c3ba51281f111a45ff343da241b2e799f8fcd4c65b904f34a8452f661737d14cf6f081b51fd3f6a68b761e840f1c09d766efc9dbffcd80a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4232ae4596eadc36f6240d31d0d52f6fe8ee2ff198316d660d1cf1111f415484225c3ede23a514c5f21e327d3c73bc05504a08571d9c5917bf2ce651;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2235a6b2be64246545e5abba60c7f34c93c11353356e574396a74d7abcae4326d7ce37fd1edbf127b270c2d875f78005b628ec4df1e0729a70017d53;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbccd5669a656658b324261756418d1abfc75813fcf2cbe695222bb654c581974155c6d04a0a58dfa1b0d29d12b9ce2b961f228980e7fd8cbd5fa6b46b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb6a8101008852310161a458365e455c94b3aef48f0ae8714d29104db392ac2a1046736c00d5ef7eb4aac014bbd578243ad590ec63a4661a1e36cb4bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85fbf2970c3811a548c667acf0addf8998030f292f27477cc0a4ca8c917cc6958d9e2cab714932c85f435c73806ea5f1f365bc2143c8a7e110c87503f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb4953212cf35dc163c001acd3bd48182817e56113a769f9eaacc2b74fa67b19e8554265b8c64f9829cc17f092bfbce2ad88b6b766865010c3f93c000;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb73829c1df157b1181bbe384b595cef5d24ced23a43f1e3107ca2313d9db27ef50af71262de23b0bfed68e88a843c0636bc8a679c110ccd0150238b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7874afcb4e5de1e258a00b6e32b9432cb2d418593a2a0d12eb0cd7291565413602de6359f7d820b49207b0dd7c60673c551d5d2dbec96ae26a81caaf7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha80a876f1dc4d9390380037cc67bf0006fb8af736fb160af31a0999d32424ac3a836ba2bdea3f097a5531d546c70c4d1d51bec23152a1ece3a86194af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7eb66082f48e6ff7ac8c7698789c2712eb2a0b0d7d45c31ab3b749fa6f4e81b09642245aa5da2e08344a04d072a630f89c0f55a67e4e5eef69e954de;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf1378e785799d7433a8c88cb3c916ba76120abdb601354de960e9182d2098c4870b0cc5f1adf1c0ae7688a5d3eeef9232bb3f2b6f4f4cbbaa3bcd6de9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd99df6c49c6ff10b4e38cfa455fc29c72d3e4071b5d635f956ed16a3727dfbf42be3bf78faba60ca7f8052ece1642f74da0e5cc9d72ee4b3afd5963b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9dc4449881287c6276b8ef6638a4f749a3c491d7e30d6eeabd435eb8b02d7aa80229df427e919bdf2e03802ba2b530d9059d3b597a3c271273566fae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4deebe86543ef4ff6004c06e0f87772dd34b8fcda9547a32030e31ca194dcfbbf46d0a4247f9de4ba462f8c4a4d2cc57d565ade971cd87fefe82c2697;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2cc675ff7fe11ed8d16d6bd9f9cdf7ce2f0aeb2c9fa3b4e73c033749cdf8f89959e20d0388fa4d235a05f815fda826717dc559ddd5b50ab3cec0ade6a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56284e968d2b34eed5562238d6eb708c9af6dfab840c548617be67e2ae78dc0511ef5fa676b2999bc17c2914ce4519b6a687a53754b633b57af2ac71d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e5cfee0599bca43a1b9fe4d7c5cb8ccaf3533b32cee5b282759ed5d12cfb7244f78518ff20bc964fda766fb6bd0dd260fdf6bb3f0258619535e0169a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h102e8555bc5186dc98ade14c053a571987796015e1ea408060b4f08ab8a78dd3b8bcf0ffddde90d65ad6f481e4d8a3bab69ff845a493dcb3bfc82a8f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9aa986532acf1b0ac00a36ed3084c0b5e07c9cb4a0d178e7dc988b4c652c2c366211032c86412c4bb6369b65d63f476a0cce212df372cd18a135dd23a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f29b5a40da96ca8dbbe4a662205d8eb6cd18b4fcf0844bfb518b0ed2f58e83f34af2a128e171263365088d10800d9cc6176af2cd9c27206ec131487;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b957e3cba6919c0c398a28c4eabf06877b21f65a8d3915e16a44c2dc283a627258638c3fdde07e26f1e0d67a73cc4c2962c675ce5a842b0ea229c441;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h945c3b5efb9cfe636edd2a9026a6c7297790cdb90d6ab846450e912cbb713e83f3693ee6155abb371b591705a2c5f13d3af0340d9347dd8781fef1c74;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h636d165a099066ffaacf9ac2af06ef09c367e3c39e0ad87710fef7fe2fbff0ba1d0c4e368ff8e03c189dd9a2527a47d14493d07d9a7f42263c1bf4a1b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3869e4dcbfe67770639490a07a6a84d3ef72c6920168440030d393197e1627495549ac72938538573224ebc9958992639df7cd77b2e865006e2fa9001;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4a5a06e09f666443bc395032c7b8121c3bbd98742cee8f001927e85e21cbd60d7d81bb248a848c16d598983d413d9f28438fd0dbf052a0fdc0996184;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d0f75641659b2550acb2357ede0afd1a999bb13102a7efb4dac03d109ebb555016227210e4a31e40f309c47a9683c69366af64657f4614b5ac9f2ce2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf825747147fe28f1c7a08096cac4da0cffb92413d90b147ac57a1c8fccb62d5b6ea1354232657758b07200d047ce61814e95f1ec1230cf4a3002cfe64;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf3f586e8be6bc646c1d82bc5858fad84c60bf2df68c9dea8221b75fcce860e67c7f6d8ad1550f877d64977d93fb3b65d9a46bd2a29eb410540399bae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdc66a5ef018b5894995eac4aad429f168746e5cf93ea4d44af25bdfe572441964b0a2747c1e899ba4b8f655a0781874f9024f83ec0f3268766349cd3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ecb183ec08c888160bb9c4cc708f0b55312360559dd892fce3b6c3ce9927dee2d17b6d550b320ea004764a81c4f620ec1e7c020268578e3f80f0e325;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha93043d115ffc467904c231f129cabee2451735514aaf04775ae2520dc26f215a33508792ed8ef4deb5a722ee1888cee5b8625df5357ab195baf6ee16;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedc1df3cb2e41978909afa094c0c3d59c42c7eb4a21168c4b0b17e8e509c917438fb082c36b8b0f5cb01131b9f7ca957117d874ccbf925ec4085f03bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3b88e8aa8c390e76fc44cb83eb15fb9544b520fa16e4a292b7bcf5ffd44b94eff37845e06ddb587033a78f63cd957f49be8ce9bc60b4f445a97fa650;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfcd19866c501dda03c8cdf017f7b64e738c65fd7f87291eb4c1a0dd20ef67587bee5683fd8bae67c44849d8e9f6c318840258f7eaba4daf7eff55aac5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ceb04d6fee4c21aecdb12c1c9f9dd7776aeceb3ff3c1a655166c5f0226ecb8b6416db0bf62b05da41aaca4387b08c00d1c83a92493496707dbf50564;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45e76ca47c71c6dc5f976409d1ba5ca32ab802460dd0a41b92d2d85abae38af0f0ded9d6a29f4ac40b1a630cf7d61de119469155761991c34dcca6ffa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h323ad26fc955587b85654ed6fb4474852854290bac3ab16242227b9b2167004e12471126b444b03367729785080d1dc8b095524f2b24fabed6a2ece7d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3fdc93b4cf212e1e822272d185448a184586a62cb477cc0a11c2f7d665a80b1cb69dcb414da711036ef13c2348257d702edb28525d57f71ff97f3bb5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61cbf2059170636d0fe37988d212751abaa66be6262a257bf49c02d582b60c3233bc8fce3455c77eafd0af1ae7f7fa58675d56c1dd4354ac80a413ea1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc346d65b82137ae6c81364052b174c337e3877e3b3685b00d6b918d0c4a56d536268761f719c2f7ff3da1a8fff75b95f6bebff08a57b1f711acde3740;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4feb409f6e4302d9e4596e3764bb31504de7142364ef87b917512f04456c7fdc7141bca4f96f8a76a5fbdd4561dd0182b3018ce263307075c7fd02f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5de49360c7aaddee757b1b57323aa949b18890e291765ad339b565b3d71a41d74acdaf1fe8cd53a997de767a51473288bcb5ae658d10be4745954b56;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69182c665b5fc99d9595f222fa21c6cb0a690d7c8e5b1de1b6d66d166c7e5dd806a054c8082f4cc3c52a7a453291ef24fca49eafbe97a36d9ce77f4ff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h129ccfa037c8bb1e5995953754a3fb48cb84f9491b673b40a49c420308c54428adb1d893f9de095fa77c4cb4f297d2e5ffbb7c1e61a99544af7db9653;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha168f383a086bdfe3b473747faccb1d9456fd668b58a57103433402379c9866dbc03c31dd6664e3cb7675bc58034e80b0cead72474b826b5df5fcb580;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd55d0d30a31c455ba8f20f53b758a802f0489613b2ff1b6b05279cfbcf5f4a5dc7c43d1ad23d88a1b73c38ff2d87f243aedb5f6fd08c2108d0234003d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90454d4991c549a7d83a9efdbd850220bdf2242ef959680f767aa184f2a9e752b982beb1f0db392805f9cb1bb4677222b4768bffefa94ef6408a8161f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d03fc0436ffd03b6a23894b1617bed8a250b3688e8e3b3d116a57c5414a0c8c0cf44757c347f81cdd5e1e0eb8b13775431b36a030ba5ad4045182cfe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf702608e28a5e113b1a0fef842f5d1fc90ee9c87b35f1f6d5edb99dea8cacb585e032fa9c1e18956d6bd97690cfea5b4500d902461e9e21ebf6b9e27;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd87463c86dcb1e04849c98b68006d1655073319b5f23a08b68463f1ae8ffb979a77ea45b9b31ede8c97ae8c54eaee9ee9c7279e91ffb848325355efbc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h339b6b27376699235096bae66e80482c824c31dcf0ef22a0ff2478a8342d13c8fc572f8d48d8ab011b97bedacc4b0a8e9d4699b5fa2540f465bfc6511;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4a1a9e0842ea88061982312c91239eb589ef57fef7ecea030efbea311b62c3a86cbfbf090393ef7f9c2310eb7d78a0e2576e9b0a56b4b2f95f7ee3a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f556b45b0a7501a0757cbfe6b517a8ae3f4223d9eb7c394912dabd0e04bc2f6c2f484100b856929aa6610e6f95a051d49fdef1ca6333b6d3159463e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea2f438eada9dffbffa4e8de32163a5748584a9f4b294c24024341c182866f54cf979a73dd0ae8c0e2cf8c0210aaac5d46e10dd65114ee2145f9fc212;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95ef49d33bbb6ebcf304d70ed65e466756ef5df54833b7fa1089c4ae70de1ffe7e05c5441d014bb184fe5ded491024c7106fc3f547921c88f975a995d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29951b78347d6d69b29c2877597e1d84cf83a3837371034abebf6088fd925c16bd74d2866dc031620d560f3ec186d454b750a232abf17dea27aae00d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h820d50bb32cc4798d60e3fc4c46340835607c45888a88a475c14803119f24ae6b36c65d7349045ba02c86d9d0adf14211914feed96d3035960966ae0d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99c1df5b0146ec255c1d0faf308007e3b20890f33cfceb7a08f28bbff595340a30b55c097409ebbc4dc87c52eb719dab44038104ec8eac1feeb34fe14;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd0da296d92d8c68433fca7e880610a20fcc5c5030e20caaebec8d1767a836ec3384e42924c1e9872e1377d05a39a10145f3e4007440cbb70f6680201;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7636852f16ec4bd7446539c976a630d83bfb076671c5c1fd774655472f2247f3d44431e4185aed862db7d77e512a02adce158961b2b90d148796f86;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he621fa56441974df75d50a2713c214d2e2df5d3a87c3fdcd55a1017784df4cef183e41cc48529feb4681ade20db1aa8d96fd5652b961ebd1e131f5649;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e00303b539ff5f07471142df74c755ad56dd43113e0c1bd29e7280a09942d73cb770cabb9570e24a961e5f4c1da8621fac8507bff8743fc12430514b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefc3ea8c185f3ee7d255fce8ac12330f2be64f97b748710e720c7f51700cf4919abc097afe8c8a90a3c02358eb69cb91bd88c3748288e10095a44fdf2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7410650a589c73ea5e9f34db7970cf45463737981073ebf619977523e94c7fc01ca1f1c272bf88433b62d8f0a37429ed3eb64ce9b3770a399aacfb6a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h473a8bcfb617c0d3726d665f03c031352c14689b184906f80d1ea455a849db0da5dc5ec716bcdcb1cb6990cb0a6b2f1ffcdf71cd26e6eec6ae1ec73c9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haddbe1422535fa99a17d46e5ea4de524ebdc44f0e6597adcfcc2b51f30875b9ba89a2e491df461d40ef27e651809d35011dce2fb5d5353a74192dd020;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bc17f2e5339e15911596d8dfd8b7e7fe20f594bf6eec73d8de7bb183d3736be84894b9c740494bac86096a6f8e5dfd26d0549864275bcdbf20d7d3aa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha674608d454cdc9475b99b1e406e45f52a128d4ff9252e03b8391e80707f0f1e5be3cf458a197798592758ca7705c8fbf40777e12210d6528a33de25c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80db59f7edeb9237d01e16aef2df7a765ca5597804680f46253a93ae8eb7cca5aa0df808bf950359e533650ed25099a505c0b1f15d6e42b8d3521bf73;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8ab648fa41334a60fdac5749c1956b1925f307ecde24f09c549720cb2947d58c6b8ebac8035d4cde5e6b9c9cdd50c036b45ca95bb8cf4b67d7a13fb7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd192dfe1b7b87662126eeb6cf324d79b8e62f3f4fe2c735925c5992322cfef46a1d578592142ccdc8df7eb15910cb23075ecd7974daa15bf81f91cd3b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcac4a48a6bc82e7cd47d9ddabe23547c8fffdd119ace8ccdaca254c03d036d611bb532fae8c6a9798ba24c695b27ecae78cc65ce4d491c61dad033882;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5ede99346fb582681bcb824f145e0b5fb738e8cf313844a1108a3bd71d6da9230a51fbc4e40951d3b4b3b6c26d15dba8eb5724e096f440ae6839558c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h385d422b6ffca6afeda9a98ae5d8000af7daa52419a3181b4a1df0ae7479a61507088ad04fe365ca2161ea4cf8e3b37070876f467aa69e9b2400e86b8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12c90f82c1ba462a9865c9cc850f27aa666f7a342d7a26ce2f58265189f9ffaea3b2742235e48922e54f85d380bec46392b7d25b25a567ca0df83a977;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a7fbec55170353e76b2a5b32007d5e1b10d8a958e62960928be87593cb30a85ae61e68e0ffc235f23844d8ab76735a98e2c1c96bfc14f20c6f49a63c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b9acea745ee30323e8a3f5fba47f51abb295a2a6332a8b0b860efc3e195256147fae7776287221a09dd91b8c4b67fa7d3bf32af52a02b569855540a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77f2890644697731d709a36f93c130c24bf63954b2c8172abd6deb62dc131baafb08b03e94098c83297c5f2aa16f65ffe4ddea8d40b75afddc401da96;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h553e5cfa92bb33cfbb9d89191ea7aec51a816a4f5fe28ba19610d6b4831ff492a57458f8a1bb8a88f95615185304fedf0f6058508cfec72d9990a6fbb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43394901cc96da962df847a709ab7b5a9f5e83fac15d61ebb6095f3089f062efc98757864029e459697b7cb7695a37f8e4583f8eced5216c5a649cbd5;
        #1
        $finish();
    end
endmodule
