module testbench();
    reg [26:0] src0;
    reg [26:0] src1;
    reg [26:0] src2;
    reg [26:0] src3;
    reg [26:0] src4;
    reg [26:0] src5;
    reg [26:0] src6;
    reg [26:0] src7;
    reg [26:0] src8;
    reg [26:0] src9;
    reg [26:0] src10;
    reg [26:0] src11;
    reg [26:0] src12;
    reg [26:0] src13;
    reg [26:0] src14;
    reg [26:0] src15;
    reg [26:0] src16;
    reg [26:0] src17;
    reg [26:0] src18;
    reg [26:0] src19;
    reg [26:0] src20;
    reg [26:0] src21;
    reg [26:0] src22;
    reg [26:0] src23;
    reg [26:0] src24;
    reg [26:0] src25;
    reg [26:0] src26;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [31:0] srcsum;
    wire [31:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he1972bc710d861cead73ed87587502cc835cdbed301c921d1a35a8184b08f4d340968ffce92583b402f71d6e783d87f5ae22598aca6fd6a71e1a7c6b85b3dacbf2d7809609f15dd68383c7fabdf90216030e9c0c90f0c4f311b858;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f11029612419cb3ea0c31c3ec64fd2d395a095b38252e97ab038b67048f761578abafc03d3f0403a7941d800008b95fada9561d25d6d3151a81fee626ca9ae8b85cdaac3ac30f6ae30813da084ab82e988a5c8932067cbb6f9c64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc01cd1081c429bf8674fe6e6dbb1f1a013faf0846a94b8b51767380ad3762a29ac0b7d1df4dea3ad75335be1031b74fd59cb526ad93020d68b97c0162b60805e7244a363da2f7578140309a84009c475fd6c1953e90683f33a67aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c271bc1102221f85e2fbb9b942a806597c7f281a2059ae2ec5f2146176ecb47c07dde58052e8b10074187634f42d68625737822be8bebf33f9a5ada96746a650ecea9b48d048279c389067ec93920e20e1776966361dfdb7d8c609;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5a6d76a920454e2c3389d5a685923a4c855f0a331e275ad57978ba225bc306555afd65ad07685f5f0df8171b6c3184a6bb74032a1d0e2a4709e08364da4664ddb96055e616042c92bb4c3e39075c7fa3552842332e3ba4c166641;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10cb153c2df2bb002faef2b378cec8e0a577ebb050efb10ce1ec64b0ea4c09e04ab6f8ab695e1660f7116ed5f5d5ba49d08783d53a142309fcfcc80be18c5bf0ae05a8135b553fb29f03d877a7d2803c902fc572cf4b20c45813898;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17d3af2c853f02e528900fb3730514225acc5c090d7ee43bce3bcf366fb62a96b2e73488b862250204a1a8484f3210f825f58296314f3b3756247e67516d5b6065b173864137fc3bda9cf4ea36332193ad64c9dd78eeb97ec3253bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec46c8fffa343b23dc992f37394018b654719876df4a5396124c109429697e79ed8fa5d7a15bc54efb3b225b9c7383340e2082e1506d2b7d66a4d0e4b1807855ff44f3cb400c1827a21b076459a10eeff1bab6398bbd1888732967;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bbdc4f5b06cdd07446f62fa6928326a7f697222deade06c78ab43ef513a513fef5fdcd6db0f4f965f56459c075b4cfa79b9d7efa7ebe6d5252b3405a46f3bc6b7b3f99a1b4cc65d5447b725dccd586800a395a1ad37a5132fa86e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177b4fcc15ad1dbd3a36cc3a5e02065864790c8810c28f6aa919e6aa09a93fee6e3b6f114455e476036e8ac39a6a2223e6c58931644896855790c3d448d54e92da389ab3ff2d9f0f0df00f82a43fe67c710524b2522095f9093fe10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he629b5a331727da571cd0eb151c429a45d0c28744ee7993d7c3389128c73f2d0dca06e35a14f80e6dfc64ac541fbe6c5f1a22988d02862bc67f8c63d69df84c4c82ca662cfa9afd42f53dfa90e4695ae77a581adaaf4cb8fbf6280;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19852e17d6f10aeccc36771cf68177322b2ec7a99c076b61c42ac75317d20d16d149025531d4a4d10154d5cb10cc22adabaeee75bcbd1b6e98bd9f2e0f9d47a05a3ad5ef05515d9f95cf66b8d84934f8a3108364b1ed3181be2363b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf8915d4c99491aed7e14089d4001401b5aaed90d67ea2f80bf2d9a45f5703a2d212f5b5d3b90bf2be91d2d3423fcb4f1a83f2ce766435658d17507493564277187a201ee627116361ab756edaad1b1802a95a535303cf21ba9b069;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137af3b07a95b37265e57df20ae547472349b28adf260f151315f8ee0b12f10da40efdc0692280e3c4b965ea56b15f9b3159e82d51f2ca5a7a2b46520ba4ccb288609dba39157fea4a47717d92166c6832a8b23082cf68f9062a94f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbf3c8918b3bcf49134752eb7219ce0d3e592fcdb1c86d6fa0c6671c94bfb9c18d0719073fbfcf93fed4efd0741d2761347335a53656d749e8f49806fb1092799827d7247da47c80f02a4b4d86e2fa17bc544a611aed4716c23d670;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h68bae3ffabc0e12bac4ab77100067ac25e49648b2fe52f1073480acf6d4ea445f5944bf69d55f36c908eb7606ff2d07be88c1dd4f33798f15ad44219fedf3fb7da3bc0a364555027bd785f994311ef4363672f9dbfd81c8c45edbb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115ccd2711455deb641c23af92ca4a97c6fe4751410df510c4ffd203f514b278f6e524ef97c47010705fc9cf14b2f2e0e0e40fbee193c181aa136ac70f9ffcd9f2dc1043a4dd64958a53d138e072f8466544894c8b7f18bd7ba893f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d557113a3e5e660b5fb47a20c01a811616bfe21677e6a10475288f310085843e37bef7912daa44841e2a8be8d9da3401002bea9159c6b0b9e74209050b058b487023e5cbb79821ab18d823bf349dc3dde6368a164e8ef7c0045a06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc6097e8d423d02a1829671513570d561727cc6ee60d2d39e3d0f57ba3e9ad85c15470406c31effc514f66fd0943bda8db16f5e12c89adf683255c9ebfcf6d4947b9c955e5b3af42d25eb672b7649cf3ff82ed2d988684c4f1e3825;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12da3fb6c043d3949fb73bd5c521c62a7baa3fc8274abd307c6ebfb539a4f29dacd46e7aa974a90c1e3996f6b7a8554a6e5277fe60ff09284b3b84fa16caddc79ff42da2134bfeb5b2bae094c45b5d6a7537b50b61238b3bada1f4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h25f6c02ebeed51f7bc0f5a1622ca168f0991dfd8b0940fb5ba32f7345a17722b2e33770752e7fc17c1ad4b85656f967d7f1aea0a1467b16648fbf448a447a54420e5617384dfe7aafe958455ffffba1e43514311ad4e21ceb62dc5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11cbde484de2d9264d363db9d82b311fab0badeaef6ace76b59d9d9dfbb93a3dc5e9a42ce4e37e1967a60dd04239261950450dbbd69ef4ad88adf94e9a802e6dc14bc9310a127eb93d422dbfe55d9fef56faabd4aa2a4575d5f6562;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111ff620921800a21b2b21c83b6762b68d2f2c62e6b79daec82c6c53a4e49cdc8cb5d801f11e126c242a17365f4ebe225d3a1555b57424c0196ac6acb9ff074a851771a5a48810a81c0d830300bc851360420643d8930a6dce47b23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1069369ea7bd2f0f2575cce07636ba66a42f6d65420988379bd4ac4f57acf225fc71514554e0595053e9720c7efc981d6477dd429e13f11dfc2c07ad6f0d229e0f4e8789aadbd9b31d830b2c4bc121f8c2c824973048b55f30b3049;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fc730fdbf1f2c12152169ea6020c409eba64cffab166c60351b8fafad0dbc90fd74ae3250bd590acaac100e08736867c325e668e5a5158ca5ab9fd4fd73976741d0c6cdfc52f2236896c72dd72e1be8b2485c1c9bc543eaa471e59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h172a5e540e1d664dc64dcee31448d6f6de454e14a16c2e7c796e812d4a9cfe6fb3db38342e253d224043e9f03f80780d3fa3635ecfca0f6cec2f58950b4a232d8f0b8e6403087c5dffbbeb96d5227e21c2b065c7546a2bda6668e84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ab715a3b3cdb37a3f9d1f848a242838e7127c5c4c2fa6e5afbf1512c595ec8825975275ed4fec5029c31c65dcd523608eec2f9144bb67fc2019d2cb1955bd41863b9b42d24405c58b8ce4718fa5565c890558667c4b892416fa17a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f75e99563a7b5182b9407c19572615dace9f517c592c0c1db2e979053d8cf75e70dfe6fa06b79b9a0e7ad3b766a092e433c5c483792ea9cd24a96f902cbdaeca779964af037a7a93369d94f69f9f7308f1f81d08375e37cc6688ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h148b530ec5481998b7c996ce9a601edd40bb03adfa1f07e139249378d620fb9ccf7f100d6c7f5c5c32623d079e5226aa15339173007fa134437bb517971c3d49048a938b6e1b3fd04486bf0cdfeacdaa2fc2bdaa23f6bb734ad1e6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h738c77d6be9ee90e2761141efd5b379b34873e16a6cd46605964f7963e85a271efb97b49011b2344ece0a284864567b2c49349926c18ca88046c08e0779ec643794febffc9fb70df0179b800457b04146886e06f4c44294e464b42;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13073503b478084a9778f6379c4e79bae05b360c39be11adbf200afff5369e3ba5aeca6d1163e1575d35b309ec73146b376dcbbb3fb48f42ab770015340502ca043147023e0c13b881d72f2f0aeefd640074aaa3aea9b430bb1bfd0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1952e3c19bcba87ea3741f8a2ba19667b2486f184252371fed7a171d2cec0bf1eaf2ae1bd3f5e455cffb0e4cbcbdd48cb59bb71510a2bdb362c39eeb92ce51b98949b978ea3b902f21a6a6d60ea811640a6f756f6e3db0623d2887f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a82bd261e1460d7a408c6027605f5180069bb062e4d8c6ce816f46b882a0adbca70c91afe94c59d7f27b0b4252d49ed4d0b6059cd1c0f17dea039fe01719b309f5d9d849f64b2b94741fe35deb1f77c2cb6de6e254226bfe03fb6f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d9951be19504a875450d7c0b1264f55f295d97adc1ccf50b4d98a0faea922b27a9f6341bb58bcb4c819bb3d263428e29fc66e6af0b612a8ccee3a65984b0a7f23d2a099b1c867457f0b2d4c683b34c077a14b9ff3a9ff01d923e06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e249946c73280321e5747c7dea971d35aa6ed9410ca6b43de5a57fbfffc6281335e8192e9562817548ec73da63b86074f77de65fec0796955f7ed2ce4b190ad96842308cee80f8220ad2f1e1970aa67c1bd10621056f00084dc12;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1627ed934fef591e689a4c603dd18691dcfebe5aefda4dea40d02ff1e958eded50b442508f0e3688ea59198552305ad1d5f9b7a0c5f536da693d0416f487381b213207374c041c9fd76c716c3ff4ae55153bc710dca8aaaa61a2307;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ef8302f98c03253f6bd5458b006769af07a825ec5ac483881a87daa5f57743b860218d56db7407959b8a85dc58a6dc9dce00032a71ed7ba3a335f494fd84c248188c70c4d60669db49663fb9c6dfbad610bacb945af44c77ca5509;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h38ab2ca48263ed504e55a604097c6ff64db349507474f1139b9cd6a5ecb585b7e28110f95c39a7f2f3c0560576f920e224b8264266cb8d50019aedb57df2d2b923cb2d9fb7b136d971b323aaef21d02e988437b2cb0024b5389705;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefd69a5a93960f41be9f61629cc6b3c7d210ff1709485dacef4e630b5291dd7e2d6a4dcb66bddd233dd6a38533a20274fac54b2004b16e1867a18c744ddee8aeaf981ada53771cd0a89b84cd6fc08fd6f9dc38f3d0690b5e1383e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9548fcffb52a411e7068a94dd5c2aefdedd3361abbb62da35da02f1fe87996309615d58522c7b14fa8811cc024ecc412b6da4278a1b8d5ee745e43da352b940f3c984fd27a969913f9b190c394a615e1a766c6aacc6dcadc62951;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd06e44724ffedd8dcf3b2c17e4ff42600b0c5a9f72e9a8ce30da8c2160d4317bdda533c539eb3a283703b3fbd939ee7d2cee59613383a1f549b49baaa5d928df59552630455858acf0dd16de832d0c8a7178661330ed83ae400d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h71e0e84dd9ab0e33bcfcbfdc183ce2753267df8000dd727c26d578e278b9b08ae9b1167757619152391b1c57fcbe47e63c82f510d407b825d0ef93582a53b2956072eea0c17f8bd7a119eadf62f193ee877d2fcefd7ab9061c8111;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h154df2d95775ca2421253f76534de4d31c560d3e91186961dda119e14b6a3b5207c6bb2ede25df703b2974d8a23f09bb9e6095d1a63a5102932ce526660fde0a74fa2234a515f0e68691f3ea113b35bc14119c968d0369458afb4a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfc27ddbdb8065353b20e11392095d3bc22c2a511554bd062dfa984ee0c9d2aafe4f39009a0f5d80b9d6678f2156fe4667f0b0886d686d2bd38d92698f88dbaebbf3943907dac609d1a8039dea83f53a8e96541a7f3c9937b92e269;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hea47cd5db246c357701a0580a2f9e5efa3add3517f11325675698eb7e57fefb49fd63e2c1c2d9ffc780d46eb46be4d22cddae0228dba70fa28d095f30eb087763f856c98d03897052b10d4016c43fc811a4d65d09dc93405e3affd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed566c4efeffe445864105305db4464b8f4d7fbfa8fbc7ff8f03c3ac80d2c668dca96cda0c212b6857acdf4dd1eb996c08fbffd62441da9689f636050c2b0c72a8af2f5fa7dbd1348e36b53c655538aa98881c98dcf00b6916ece3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h236ca6999b2b2ddc59344f82c62a7d24e4b27073a45d4655ccf5abf054437c6659cb92487b7b2e6c1f2b88a3259ad354a92dd7fcbc7cc9b6721b0d102995b3cc058ccfa2005ad781155ce369d557569cd430468363cb388d9ada95;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha46e305487e18a023f154c7157278c8c4be61d039d6b2dd374581a844f605359d340f7ad574bd1c6f18169bb017fb91ecb602e38b4b25789a18c40f0592ed224e627325d8a8e6890838c2eef415320c9b2eae43dd0432d4c9698d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d9f505d2cfe65e58b57071616f78aaa3f2077741e97365c0601369a4217dc3f60efa4a26607425fc2493ff4e07f7c6c2095bf4e1581fd6e31d37edaa10e8d5670eeff8a721bf2056d0aba651a2a668d0119808013b2a3504a6a116;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h196bbec4691b6448097ee1855998acb63870c1f6e92cc1d0a7794664eb2fc22280a1b2c2a14d82d976a2c93b5bf00f4487c7edc4b611269cdb8aaf2b247174b42c405e6b75f3fc5f0480ca173fd3a01fc5db13c3826e19647bc532;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15cbb91fc03592119ec1c4eaa86d5ffefcf3f56e7bad1f7d28698ca535dbba88d59d76a89bf8f7d8b0be93b5cb0c583964142c324226a62f7a88bf58c56f1d4d5e2d887f8a054318c89217666444fb1e19f2416a09b09d6405c7c0d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156fbaaa1d3a9009b1fb28f5feb681c779a6139a096a1cf152a4b0f8bad90f572ce5f6efdd5e0324e559df88d89997b7a3f607796aa367aee53931b6be35e05f13b245645092e7a289ce35181638fdf710932c9207ef4d0e7a5e480;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc45062313ce1c2c841b48bd708bac0a67bc864a3099bb752ab944e5fd1ad0350b96c582cfff3cfe71431129857581c65c3728bed5c2504efae3429cddc8b466979195b5b9b90f22c8ccf26cee37b31076cf534d2592a3aedaaf4ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h189b85cda64d7233e4aa3fb231962611ab3e7a46aa45531058f7fb8b2ea05b371d35c14ab1899902964daa1477ff3613f4931ac46c1d53260d469eade809c12f15f2580f22fbf4b44b093771b0c528efe078e50abcc21a4b5c77e1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3a05977f88efaac7cbaef9c85b523aa6d56d5ab95fc5584feac0e22da2fe73e3ab2aed5224f70495234d40efda2a742a413bec06f3e5a430d08b0ee97a9e1d30c5303949ff7917382441f478dba032c35c86978ac7b918aabc9edf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24bcaef2810b5d1f1d72de4e8b0edc6bbf165f1f0ec26463335343b5405e3f2a72452ccd201d62d0b13bc13ce82e33dad934d01f254011110b272aa081c642474233f30e4ee619d24b764a99c4c86a296d075b407716ac68a48190;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hee67506aac3dfe67be11ea71bc8b909b5c504214202cbed4ff04f5a02825688444434b416c58409dafa3629ca8da2346d115b9621e5ad07f606765baa1f633b93013bf98cf8d8aaa366142b8430fad33a01cd45701617035a6c74a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19da00a52497ea6c977775d15be4b33d51a67f5a8dcf575b0bde3e1598160575105f709ed21c7c5c52dcf006e1d785d72afaacbe0f52d89fa0e7c8db947965dd4a9ce158f1b3639eb62aa8f09761999ab19e6a2c5eb6b009b4edb51;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e57b43b7d1d3146a666e1550a94a5dfc0a9be82abf5bd6c9c744f499cbfc64da936e944490df4b806f8ca5f92e2bff92cf1a5f9552ed378cb27ffa4cc93e750aeadeb5d5dfe90fa6735cb4756f8cf93fdca7ea9af0c91f2bed689;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd46a7d3f4565f2032d2e7be2c8a097a76ce296a993a3ba349dd632e57655074c3142aab992b31cd5770a201555ba55e3eef474711378032caf1f4414a1474ab1463fdb58536b80aeb9520a562fd828277c0eaa59f8dc07fdebb7ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1477bc5c922b99ef977aa25e15d38954b499510aa18e5ec570a218a9a09b2034cc4d0b3823297375c5742584d6aa5322e1b2ee9b7f726457e3236cf6b6b3bec03efd84c600f7a87d8456ce3388d4a23166fc1c6c8ecaac6b9ab901b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'heb94efcc1cd1c77ab3ef348aedde8c8bc3f822c3f1f540684f2f7f98a7efc6eac6f284f80cfa34a616263d8b31648555405596ff2b8db8a94b94e45626acfcd6d38c8815805f73d179640b815f877fe7bcc92c01440ff0e5c924a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a596cd17ed6100ad1b2c7722c714f1f1d3e6e6c3182e155c7e14a4f80efc4c2aeb07c3a8cce2dd5fd9349d05eaaf74a4f1adbba322354766bf9445dba1fdebbccd5770548ffaeebd555f879dae226d32c2c309da1e5a30d57d0e98;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h65ecf34b19f95ca157dc6f96c6055b71d1de67801fbb9432e62cd06090533fe91145604bd9495648aae4b39377a4fd20b84312ddcba24d93e6a48f1089d268236ea054c7342ecd932fe513b7ae003fa6cfbde325fc3327cec6db22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17eadbd3b532c0b243a11950a5852551664f855d2eec6551c2c12387213b1c63a7235c72ae5345d79477449fa014ef79535497ec62a249681abbe763030274b19b9505f7f7be7a0453e61e237f8bddd5a4c5679d63b943a4fc2c69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h96f65518ee6d9625a4659873cecb75cfc17d82770e6268b2eb7f638f3991cffb91d462ba699790ebe0bf95f69e1a27d6fc23a896b668d2eb8e22c61d414a9671995848a3f02c74f1f1bdf08511e5b06b238a34a43d27392201ef8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15afb066e13e6e7464e1ba4c4088d24c07fbc038bd78859fa1ccf70b59178923cdb68b792a657eb5457c0715fa9c6f50c00d372b23ea0c26109c7b844727df4fb2ed7ad836e3025a7d15ecc08d4e26903793c44bf8294a9f8a57c06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h355058093814c8f5b1f954dbb4b052a64181a0f35efa13de70b6c95927f261ccac7f03aa2d4d2e08dd2c1e03ef3af5252a1d8b5d068fe4f4096e51b8639c2659e7b76173dd935f7dad98a586db81ae2ccd54629b44d6c5555b4ae0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a74a16d0e908146daf59a0033382d13c185ab312f243fa38c78ce0a39638ab6bf40fd179126d3b33bc835ab5c222ac01c901282674100e789389fb1d16918797abad091bac0d85791d13c467c53be3e94c014b7ef1a9ea1bcc9be7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c20bd9605f8740a071a3f98dbe50d5c82d721ec3a019f1735075facf826a193f6c925394031bfc2f7570a98d33f009ea0935ad75b22ef48f3596e14a85df3c6cbe1cb530159f19201ead1fd3b2ec5fc4070f795d65e0d0b6216c68;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h20fb9c9895bae03582973b2c1f43cd3e0770f8d0b1609f17c3fcb19850fdbf618eb467af81e192860add11c4ce49e9f7ca4941621c0e628cc93e64614c2703380021d9a663d46685616b10797ef634bd498f6ba748089ef710d74a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf23d7e6cbdb44aae4fe82054bd2b75cf3f5e6a70455f3ca8ccd06bfd5a3a6e36b6645f2f0e5fe520d839f3c6fbd66b79082a7333f3ecc616489e63dc7a901839713bc3167af1862a373215f6ff6eb7e5ae3e976f332014ca30d0e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b18d68c7005c71fbc9143747cc3f497880aac458c276567bd588f2f4e8af7a75496da3cc4f2e4281b257a5392b4dcc5b0b030367bc2feb4b99747f6ad8156f5a0bdac30dc9eff5b5b5c5550fee072d249ec3c2ec534e6c140ad767;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1409bb89139a04dba4385fffd243a82882782e88bcf8587ad6ee4a0f57716d6073610fa7d98d27ae6d99c202d1faddb0b838851a60aa57ca191a42132ef28940685d366812d6d5f943219b530b3b2f396978708b9d02a8975e6d760;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17e189bcda58790034ac80800a25c800827f5905b26c4bcdb3fb59480a8e978d8fd458020078ca4e3b23abda0e34380609985b0d905fefcbeb2b45204966f4391ec80f5e77a6d2a3159d23217e889f49db5e9749980acfdbe0a819e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c0ff5d0c613ef51a8f244185ffe4266e03d446b94235689c0b402aca41389872f1b08fd34adc51ebe10d43d3ce59a6e2488dd6e18a81e7ded5dce55ad0b470cb2879d9ede03463b34ffe9edf86f64856bd2c0c2cdcdd89d678912;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb21beb563d7a7950998aec84b19c2eed93f27edf32489396b69250dbdf4a80e0dbe45cbd59d3330f6c15cbc6b1950610c6c445ab86f7c6475386f8489267e29d2907821df562288b336e0a567e85268be2bf292cd7885a2ef54f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115b8d526a01a85b4b40a81daf658752b6f66ce4c97e21a85a4ed25639f61fbd24d89d156e2843005a31483ee166a3705812643d415e52ec7c6fa5645e2957bd2c4d267817b6f94ecda7f34c3f70a1efdce7141a1abf56d388c8ec2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he6b2b6867d0a7b815cb7079e371810f61dd846e09c1bbd826ddc5d0d2fe2b63f8fa6ae718bb931e0d45c5aa7e261a9eeabcfaca670af6198ec303bdcf864e86f70230ea68b070b5737eb16ec7c71ea2b2cf6a3446690ce1b09e905;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbfa6826006d738ce73ae87894706450a8474352805f7b7a55f408156ff4ddfbec84c247971e3d21bf56ecf21e97bafc18ee93e23934b55ef6e9eaf0c1409903a9cd71c017de6b49b6d7fb383e3dfc7b5acb40ea8f2102c97479e01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4fc5ad1f4141d0628db53f9ed4377be9d5846649bfb7266b956839531ddbd4b24df7f1d1e63733286daf4335b8750715f5552fe92ad5b8475dc68d9d1f39d6c796121967629cae56abcb193de853d63d0f5125bef9d189426c445b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ba3c187b52ad201761738bb3fca17050daab7cc7d8e98fefa3fc8e271182806aa10f59291615de16a3e9745e6140d276cdd2f2e8b22da4122f1c7c13c0fef8e9b07cae55675d71b48ab6584457d7ff57a67d855e186a964d6f1eba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11787bbdd10db4442b5f7d6e1f7ef01981bdc980e03a7cbb72790c65f028267fcbdff0973a2dc308a8ad401bd51da9b4a51237ddf32540550e32b8abb06d3b82ecb6128324c6d21cb216c183c588ef8da16635a91ee169b48ba39c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e6a3111e30ff911a1f6e2fbc65d84fe00a5e6de666d82ceb2e55dc1d522c200e82a1fa8bc0f5bc9773dcf05862d447e094e1fdd29ba26f3c5a006d524921bd4e2dd1ac8883bbcdcf85f9a13f931345b60f42735bc53c7b1c08104;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6b78a135bf1ca980eefa7b95c7d0ee52a8d40083c5ba8bae204c281a264267f8189398edf95bcf13d8ce5d2b6986286c7991814267cb65df722f10bfb123a67683a596179ef0a0eb9107e5395ee512b2926fb448343d57f47e344;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h30d50bff33dbb3b0f21cb7fbf87e84984e1f8f0fd4801c635630249aeae4bf73a3d4b3262cb27432d70503dd5f5113616b69ebd813b047726636192514931ee27f5a861b4a76fb0c10218b074158a70b24a0081fa19f592708b615;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12a5c5db85e941398cbcde1b262ff9dd586639236bc3f0a1e04c3912eab4c159139e76e00c2b15d987029b6467510559a38104bd81624ad1bd6fca056846d29ded3a7c54c7cb0cf03ea05594145464ead2c085b78d04fa609ddc11e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb3ce5cb15310051490f6ca7e4d1a784c6edf4c91ae516d91c3e0e28a59f2ce3c1fdcb9264b8b34c8b65606e7ab64d49315c3986d22369ce0e64f3b168a81e25f9f9b8c818b13604cc8bc071d9702196c5570e231821464b7acbdf6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11c0b84a6284b380e19471fc866c585764db881500a1ed20af9dcc6cd6866aaf10dc8bb76f73b7d4ea10e09613dce49d6560ac9e1a045fb6ee5dbdc2b9fcd21b21403c17af9544573a9fc3aa8a53e1dde2490cea7e77d3d1880184c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h69cf4112dd99b1dcd6e927c83c5f2ec8e3d3e44675bed02de2e4c1aac3431b593f3a71584b432d898ec38bbc7515956d064f83c72282658983bd0d7c1643d91f1d344f42c4908c3b14d04eb1004d2d5316d55bcf299628ac89e7a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111c8f2c2615c9cbd092e77250d8932172cc5f4126f6504e1dd25592fb3dde9f982bffc647c656b66dbe7503886d48a9f0bca897da29d9940f5aa2a2307230f86efd809ef49c15d356b3e6395b49158d33b0710b2e5cb5c603993c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h869dbaa3bb98d26306038e91ce271e338b0a219e764c8f35f0ab713e35dab2696ad5b577c4b5f4ca277d8e066adbbe5f52600093c881fd0ffe205057eed3912641470c1ee10fe11b4d52d1c1e96915987fc2962f5405126a353591;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h611ba1451227fb323b5ece23f5cece56fe150ff04a10992cf03b679247948b0c5ab625753c688da68acfc78aae433dc060c8590cd06d24a4881a38b676385c199f21bbc368513e741342d26e3f74e35b40887272834446a7d8b3ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h698775dd5bfdc2f09b4bc1a1709a497e32d1ad0b5f1e76e78ddaa8514e569e930dca2f8e6f2ae66b7a42c1765bf0b0932c65a2f49336599ead73c708d18c5efe06816b2ffe21959e39ef5cc832dbf866bb7aff6367d011464d029c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbe25b6f425ac4a255696955ccfd408388d29a9c66d55a5a931f343bff96dd61ad2079a9af8e202368f7e1b710e31026c1fa5b2446bbadc8a4ec82924cd46663b0b96ae2cb3195565561515ea2df5580177a482294dc7b80bca1a1a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1273e38f4ab08e2879eec2ffc42a9daf3a30381e811c8d1d578d65e8002e9183d4c722b87925f4dbcc468829dca1ed0c9734b70ff87bcc8465a6df5edc66d9f49005625e89a20fa002f774efa238243078ad9eff4b20b65fd6ebe89;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b78f61d4713ff9c4a02dc48e51bca2aba5d891f761396abff4f4ab010c21a0e8d341882bb5e936c8f55b13a510cb4a8e736de54d7cd108df31e85da9b507821273e897bd3f2686f8c446bfac70653ca99d9ad3a9d5e00750be0ebf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18e9ac5ef4cfcdc1e5bb639aaeb64f76ef037a95231eb729b814535f4584e86826107e4ce18c6fcb9e365e168f8247a52d5bf3e7293a6aac6f7ad8bf1188e5a5c0a47f64c8118004e45b52deefedc01d3202646fad51238b4c187b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4427454d97c96acf9f6571c80121a3f4044e9bd7fe1ccd80ff80dbaba10204160ebff2a393a1eaea9ef3dcd08af64a1073addcab6d53aebb314ddd70b11ce945e1888f0ba32f39812d3f8408e747294a2bfabfb1cb20f3b6c1331;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h138f802d7fbbecd286af13b0f88658c6794d78cb36b6017f06d9671c105728fd45e3d912c6dba2da05a4a1b649d2b5c650f3dee3578d897cc36a14ee8dfeaa9006e0c3a07ec3a88951158ceaea7851b2b5f34284679ac5e0bac7194;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1479574c834a08d8575a6febe7c8c64278c7865f5e7719797c98158a562feeae46672849f7cb18a9b9cff7dd7d6c06e7783855a654f3dced8ee05a3047545f5ca54019f557693ba94367152dc3ed72c398d040a9552909c91bb7cec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10f9f9c0b77c369309febd167d1a056f37a9dd96efb440ed647d24c5b281b2942e4555b108b9713296d73e9c045e370bdcb472b5d8340bd5925dc7551ff9a1c29112f12e2182a7fca8ad536140e19be20479ac518a5a0b37e15e28d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5be0a9ecf84bdb3791ce198a380191d939df8726197095e9d11a88583c9391592d82eb9e00af5a01e5c2726595d711662ec7a6e3098318e962c68420dbba289f1d4caf8e49712e7f7eadbd80490fc0e6ece39264acb7bf72e26bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4f886e46d02d8b9e0fd34dd9b490aa310b0b10666f70a3680206fa14791c9ca8fbd50e30e90d4789d57d009a0c65e4eea71bc82572e76fbe96eeb353a128fac5dc63e4b2eb807a78c7f1c95cae3fb9b7d78613cf86d24489404472;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c41d0094ee94b824ffdfffc4dbb021705ef3ce55be64bffdefb2592daea8ab489373a80899111f461542bd5038661e217a23c96237ea1cedf9f57905e2930a590fbfeef540ec3782c3d49c638a58d561c1f11bacc1b2e955259bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf86d248184fdcaa99698205ab07f90cb9167733a92960c0bb7519115a557d56fd644a1f0cf28451c0556d606331729d9ee8dac3be4330416f8b5351c746320c66ee0da2796986e208275eedaa87a5be1bffee4c08aba13613b776e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c15ab6bfeaf47342b8129c9cec14397aa0212a84c2118db8959115d0b994d6bc6406133664263eb4bd297ff6d1b336fd631ca9cf6de142f6b3c574c19948f6ec3153cb03245f72265cd38b31c0aca5db9c364ebe15d851c6f0905;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h123182ded74273e2fff2d5998a5c3846e8187d37ac69725a37c5e437c0fc2db27fd0ade8d97dcb61975efa799b5d1b064209857d6379ef2c38934c225aaed8ae2dca24684525fd8cf2d993006e5df7855db3ff4bdda6640488c840c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e77cab86d4a802984c4da4061c3af1e046fba3a34a8da818a643eda83621b105a9d8d118222214aff66c05b228c8fd47912813ec655ae772c96282111e4cba548f2166e07eec7798e379dc378fc3bdd607098cc95a09bd2d40c404;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67a91b5d54b4d9e6cca14a25b2128fa2204e8381790d270c46b2956068cff2ac2f5eceea965f3d82786d2f720f850da8790d8b08001df8a24814a7e9b9610d46a39cdc891106d412a7d125f64c4ee1ccb417784a40ce60b58fc13a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h176ab746f176a26c6faa361ecf505e572cb639e2074aba244b0678b0efac22e3f035d708cde380c4e045e4caf911481e18b91ff5046cce1d261eb007001a64cdb79b3cdf311c8a1dfdde1f76c900f70709dbf0249ba46291454b9bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27cb48b57bdc8ab878a6cae70db409f35533048a670a3043fdf65266e11118f4d25879e0565ddf9af81d14536d725e9af944355a6b6d5e1115795fcced91ecdd2273ca9f9390e8433850af22c6240638370f723ef887c82dc5f25a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aee01c4d95d848cf6a40c964c9daea187b8b8d41c5d4633d9ff9c0202c8ade6765efc550780b6a2c2bcb30c0153e7e837f10a4766defa0c029176e747c36cdc56800fdbe41370d7b5db94d365ffaa24ed35307dca4c235de3c2b59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha720079e71f63ed10a9ac0922af170de0a8dd3ed923b04425a20b573b2cf43f497dd0ea90ce674a78e2a183f6ec5ce7a022a25a967972ba032b696ce435f5aaf6973e80961d719e8d79c24200b857c8d5c7b9195ae4257e640f589;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a9ec45558551dee6eb73c1783a6d0583f864da7628fe6f85911e6d3973bef1678cf6cd73e1691dec9995de6a17a6652d1ca74a274f62ad7c7f770b21ccc751d13ca0b2d14e4518ab5e1062437f21d414a97fed1e914d5621a8efe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c675ffdf2f493b7cb4fcf3c3fa2a640ddf0c4aebf534ea78f912cfb520e147a4a01d610566800dc9616d4b041ffa20f3c9f5fcc2d321d8caceb729761c22412a7af076fbd715c93362991e7b02cb1fe9a5ae78948a0326e6e80c96;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h158f149bc6453e5b7e2fadc040cb49471fc99cae7787c8c33b9ae2d58351b8fb5e1ca6d9ff6282cb1e9b4df7d37ec569f71207375502d724c556064180666b3dd7df4619006b13a79efa9c38df193cf664570b7e7c4527aca045ac5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h613856e50c5c6bf88f18d9d40a8ef0e7982811bed0ae6ea77caccfc432339b411d9433c5171142d2ae4aee52892d5995006dfdf22170e558e20888cb9ed01fbd681fc31a3a59b1daf537bb7d849bbd49e3e6016af1ae29896de3e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ba930eeae6a3f11e06b51c9e85da55d1e479aa18e7d5eb91cccb22abc1027fbed1d8b2a16a0d98183303ab7d32dfb8936e8bc734dca74ed9104a9839f15a8da72eaf734b457bb36372617e9d0c9e31fdaa1292ae4dc70e5b569c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136e2fa41aff7aeb8cd401779c451daa38767d416ef748f896a8df3bc288f3b80146a2e94b54ccaea877541d53081855832bd9f5395cef76a90953846ececfa8818bf073c6b3fd8ed959dc8b6068b6d34e2d5756c0e6377991acdae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9ddd2885e373a53967f2923ca917541e472d84fc308236a6d1c066e353dc710a994ae40f1fc59dc02f29dc8e7a015fc294044db3820e5fd02c5f94af01a62d2a0e7b8495a6e990237f48a694a16cd10e54b119f4162d0aca5964b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ac14b11bc29e55dbe467a4cb09ca7f1e8b6846bd96a68b523aa7506fdc95bee9177f53c69a79277e1fe899e2a3da45ae958e36548f86fd3e967ca58f4e5456eff092828091f8e6383bd1c40e871134eb44e2c8688f97b7f6df3d7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb36e0ed7034d2d331ee0cb2cdb5243ca3ccb04a944de99df2a91b13f0d3e96d5841961a5ad286c9bda66e10ef0e1e8f579dea9024dd04a6858ffe736277d355ddad19033f07c40596c8b92b122d852e0cbbf6e9a1d56ea2f659be9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3464f45ff3776ebed27b97c5612fd51e0edd6d1f5b55d25541e41dfa28686fe0fb10370ce828db4ef9ffd9301b497fed0df3859d43479a7f17fd77d935c5215686f4de9e24c32b9556a7810b368a4a2d25ac9233700fff1690abe8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156ab4f76c3b2d46d558c74d8f75a92976163d1fb051e6a82161cb505d66921007390b382259a45b91d447f67f31206cc0285394ee82ba718e773f45cb34424a9ecaf9563e2f37b2bec9ea030083e31e36ca097d187da5260cb60fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h139423398a5a547eff0a784c115feea0e05fe242918eb02ced229e3847b67292e672b81a0a93d17112da47556c455f0d038ecbcddd06934b8f9db6b8746329e6fff6d42bf0099abc3de700500204b366ecf16fbdaed2618e5939c14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h107fb2f48cc97bd5a264d5977c25c9391cce78ba7de6eead4dfa5ea7d9ef6913b404f5c6f3aca7c4ecc5c4b20f3e2f9af233e9472f696f620cbfff10d3d0994dbb2c980d3d4424f397797c2f2cff083bfda2a05c5cda675709f1b99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11a08dc9997e84639fa706727963bedfd2fbebad61bd7ebd41f21af338cf11d8ca41b65cf0d5258ef81168aa730e074b4feb2456b4a22ebf501b0f4d1a68ae62b36df45d7c25feeb7cf8e2b9acb9e2b11b5f049fe2d0e380a70045d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h337011bcd785f577b55013ed8aaec8457e1f7fff84c03c780531f19898d62cc66e375dc0ad22135b0c9a7bf794cbc157f931d7ba69a98a2fb1181fe3d2547848e13220e19a667dd9395a85ea957b2826e6f41a9111654f186cb8f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c0ae1f984ef673e872b6daaeeaa89992c97a3ab7588260f38621741c787756a7b53d3f7fd815209edf04fef7deb372d6c14d5b99796e44f07d620b89b411523ddd187030bc69420773e73bdfc5c55744fddbd620ba86ba836f6d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1234a7b96c37d251edb6f02e23f06e847f303a7b88c692e0ce39861f58da43f206da7c528b1d0c7a87ab8fe96bbe83a822c0da5481464ce216c5013b64c27361864f5f25e1690da9706f7d92c40b6fdb79eaf21af6ed54a42f75b2c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb865a9f6b83ae171561070f5eca8ae43aaab7e54ef25dfcc35f993b187aa4ee78665b3ce3575840b0aa76c88d233b3ba8c9334af47026a89bce120fffd08b761771268c301765127266513a77d21a43ad6de6a117ec36338801bd3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b5030d2a941ef65537a962b17161f1275d4338b81576b5343345b4eb727f847b15a936fdd5f43f67b2355ff6c62c814cc71c759d8137136a26b6716f1bf9529c51c46b83af4384406639c19f7059f74f1e9d484463603a46639bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7d7405aefb008f394af4dabdb3b966c0734c74c32709eb76468a0aa9e3d1e21a5c25ad4b732e0408f3eb1673f2087f549fdcd8cb7575204b1099171652b834400018e6f6dbf86bd0907f79910b05358acf29da61aaf307b10cf3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19160e4a89783b12a9e746a69cc207cdc8864c4e1f6d7ae2edc79169b16d9acfe7e7e4d8ac5e577f49e5b24686b75faa07643a5db851592f00bc31958fbeef6cabe2adaf957a1acedc9cafbcc31b0de2e8210573a999297afc387bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a800cdab42b958b72b7398255030ab8292d3c62ae9a7bdde19fcdf7ff708565e315494332198231479eda85007d2c76b5772967dbe26b821aac39e60a3017adb3f4daa22bee2f57099b36ab34ea1cb022d8671d86b5703cce1d4db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1edd323d38c5de255e476e0f5487fd4fa132a6f2285db80a1104cb5177e2072a4190b937188b8c66319657b87c55d402130c7059640830077d2b1fe84e659556b7e06cb36491f19395ae4878637c53317d00c93de0994ddcf1aea14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ba04fe7e9b5537227807474084e70a219dbdbe36de064c2f117a6af3a8441ded4727c6b6ac7072a7a2196efd73ab6668569d4293f69ee30dd792338aaad71940e12f9632d7d2e5a49e270c585fc21a3cfe655448ac82ebff80442;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h54eed7ea991a7a36db21316b93330adf0b6fc7782b74067137cff5aa7e03ac798e5ae124048bbf79a4fdcba4151936a2aa808a9e248c6b7d199d6ac13bab56b403f485a5ad8c78d74566eb5dab87ea7109ec0a5f0f6304cf77ae57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18229523e66634b97292bd16a884c521ae5c559148cd0b6358182dcb6f901fb51e4f0bfca6ee8015563fb3bc4e8d88f581bbfd84a8625af9105170013fceaeb1701fa0c5d2d2e1401627056906f12417472086509db30b92b295359;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4eaa4df8d2c6627ad368ba18d86cb4c8e82fbe7d832b8cedd8d68f75b29774bba8b68e17813798e7ca4ad08583c68943aa2ac9cc38f2abc5dcbfbe2ab8c6931db53c67a1bd843d1482e1be3b375ee3b47bd10339b1df11a61b162;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2372a4aa9a304e89dd440b70f6c3589a44cf31719efccc5637e1fb2f72a1a2661e4e0e13257b84453ad6b70ed0fb30025bac82886f825f5f2a3bead8a78eb5fa2ffadb6bcfc7d92b27ebd544aeeceab81d1c40f601daf273a31ea8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd6fc14955a4239db90d25688d3a0ff82eed2c5334393b35fc512caf6f49762f32bc1ecfa3eef804b0ee1c9c2150ccd1564ffb8861a48a8056e447eab04fcd42056242a99241fe33c856942f6470fa129516f0ba869929b96c66bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2f2d20e262f3fb995ae13318a58e83d9c8ba96e2f8e0d588904960bdf20ba01b25666c71bf2fed526456844c2f455b5408ee5cb155d294822e0b4550b72ea104beebc8f0cbccf373425e63d1667f517085b31bacc38e827b65c9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f30105c94a23298749d4d968685847c813f847236ab133afd472d19e4ff3683c01f044cb9619a16d24f85a8e9642073e082dcd0e16acc6a18ffa3a3a40b03464a5a12b83726f5a10d47ed39a4ecf51a9ac5066118c9f8f4821a5b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5c085cb197d3c727ef432b8a7c956bde921564eeb595435bd7a98b9d3ffaa555f9cf96ff410c2bc76ee66a50004c81a983d2c7eba003ebdb210ebd33c36fc2f6a1dfa5763e1f299d7da710dec6c9892c0d37bdc4762c1b4043594;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haed56fece2a891da60e80bf85a4557a07fa719ae524056061be6a50a7917d71905b657f94e40f969bdd0061c1d80fed1995285c27dbfa36bab9d9734f7912237d54c54a3d0e02428292d6b4685b71bf9fadf15181e92b38c72c30c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bc61808fcbb768a17f2d9ddac99cbfe5dca00a3c53d433ff50c6e0a72264dfd6a375f933343360ab7bffc72cd8314e640ff3d9f1c760bad513e8bf1b24f545cab5018122fd61810951c568b07550ad3d7d0b2e294e991f8154fd81;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1003e5552a54533504d43c4bbf61a36d52ca2d2bb0568c96fc99368aeb31240766464a8e3c16c575c793546c6c1dbe4676f25c719fbf83221233bb9b9f3b1225bbe5f73490d043d62a52a85194b2b512844ac86f4126287ea799dd0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dae7b891ca4f92ea3e333ae9bbe43a0815abd20b2c4a7a3ef27983145ed93a811478a205d767bc7e1964f926644525f6f81ea4a0027e6f6ee32eefddd54264db080b8c9f5849874ca481ca0a901e99759fee26bd0637b46ed6e16d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1628f447fcd55c7b5a8b8e5ede49e370f9798d5fbadc12cb1e15bfeac1971da35dbf6cd4180751fcaf2df18cac1a18e1cd562d6a499459317b824dbb8a647dbe69f48761008c61c68cff3ae20334e67d716b2ad5b89d1fcfeeb0f3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he04a09c724c156fbca29b7a188466ca76da1b7e72322232d6efe121a68d298d6c721df651f0c8a47feb180a0874172267394d344ed339e4539a97f5b9936895a5f37d6976d4fdcaebb37f4cc7b75ea110c033b7f9ec91ed7b66bd4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12bcfd09c31dc130be7efc997492001c92dd7c23609a82689c0a3f8f1e5089871d7024b7b98ec20ab10ae0054029ba7e237863712c1df3486a1124e78352f18610f785d4736d46ee3412dac898f2ea2f47cd613380323f1cddf0a2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115c01c1f19189d4d6ef73fd94ee8aeb4d8f858fe587c454574111419fd1536d3eabf698216ea8bd5b0dcf8b6c709a2202c22207b25feb93e0c0acf22b1cef35d1924ac731cf17bbc14d4f3b2f7761e353dfb2aca0efd99fb17c636;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hba885a798d9d8cbe2f5699e2b46eb8900827be56900cb5c0b4e8686e2b3cb03d2fafccdedc69e88788fc5b45649b705bc5b0e4c8eee20a8c466a491f809d9c7b21b5b20cb1306bf605bcda528d01b4632f41ad3df29e44504ccfb1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10f9477896c58586aa14ffec148b797c17e1694f4d4a96d319987710f7534d05b870dc49fd1e2a19675920dc8bf5b2594d6082125b348812d159232e386fe2500aef860cf537f29acfbf0c7d18ebc65afd2581e34048b19c7d75c99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12428570becea5e5eb4546964580b285f17e1532bbc40ed5bb32ac52c85d8ba24b78bd7ac22795a0132975927e3a3e29beff38868c83267485dc896799caf42452d9efa1040ea0f54b6d4c3c8fccd9891352f77b309b21dd460b586;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h152efb0c70f59588effcf75971dae2e9521037ff57e41085f8b9039afa4e9be4f4eab6d862a0f01695a58fec5f2cbc306bfdf7e297cfaef42c95dfb66fc36fe33617ef51fcfe10f7c0265b4de7041790db7dc81054d7dbd9b3f3607;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53424c6e2a6d4d832097873d13cab1fc8f29879aeeac91546b030a5f5f22ad55fc12e9c3dcb37aab5683921e24782f7eba812957a34d079f2598c37eada53886b5fc0af7b5eaeddb3ee8cc09d0fddde3df8eb36cf5683821752333;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfb2884459ff0e1a4897092da4e3937209a38c648b64d3aef12d228cf0c0b9b0740bde4b28d19c05ea1abb8d98dfac8cd6566d29f597c8e01024ec5d2df6ccbcfaf228c168eea68b4117699198d478ce78fe54d09d10c4f3912d8cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb1874a3f1c52c59d0748e0fd8b771b8d2a887a59cc031c41d5ff0eb4881e1d493a2b296de9c3bdb7641a044274aa7534393b4ce6d137c0d123b1a0d629b59ff19d9a985fa5d084e94f9092d049571cae83df8fa01c2098c80078be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180ea35f78a5b12d7251db6dd44692f033b6de005a88172456ae5bdae134ca25a0fbb0fd4801f6c3fcc9e559f2b3a1ff1b4a718aaffdd6496cdd4b3db452cf650bdbf7f414eba01bd98ece0e19cedb6c9bc8288373eae325bae01a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d9e0dfe15ef9f30c258e35b663491b5846a061585c89b842dd99412c89c0c2cc61cb003ca198bca34fd16ddf09c52e5b5b250999c1db599b06038b5303b7b61737dbb26953fa8fee11e6f2f6e5ce9bd09ae610460cad487707928d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h292fd52855dbc2a588f061e8df07178f10b9c856d7608d4b0eecfbb2a9af1c7cc797e71423186944e6912d67c3f8601e717c0110fb1fff7edc30106484b107e6974acdb94487c6f2eb002de90dfc610d88335466c6fd4b035cad91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e103cdb84e1201c512bdd03fdd33c5123e311939aef49ac28c454c856749843f58f959398131db3ab94f6301f778db521f740d9475489ead56c707d509cfee44b33fb86554c4ee72f3d1e311cd953cefc4051bbbee7d26e2c4360;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hefad2246263e479190aa04d81029e04e055052b907e865d10409775021b2eb9d6df0245d0de4c5289aa9a8048763aa75b133c9c1bae1a27f6ea99c3048772c225b67e9a2685ea9c08ce8cfb8a50708c7f8ba7ac56c62adddcab76d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h74f45bee13bae89bb1d58a8481627bfefbb1c3c0579307fae8da0a2bca700b4325034bcde9d7a921afd70d08401ac7470431781784dad5b40c3960c0a2733f2d8b156f705ec00b2e9f434072a24c24cf7d80e737e595d66983c4b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe6304f8c1d35f6e4b3be529a680fd1ee45e71c2324cd2587d0932ed5065374f1d7cc2a1cd5f30645d1ad45a76009acde872dc23337b3b67e80ea6167d8fafa1094f9aa6f95f6028de9f03eb13bc8f93c786e39aea8336d824575;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4bc7ebae254a06b79e7ff5e359d6bd0e1ed7e21fcc4ee48a10f54ce213ee6c01125bc433e6c1f8a589f5bf0b8e1fe48103c008ec8240849279bfc161e51dfaac9ea4ea8611c41967448f79c94c956cbcb3e12638fe466be1dec81c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13e7e0c82f1fbdb11b34a3dc29297cef21e4a238df3fe41cc177f4a2a391401a431ebd2d82742270261f684b4ebbf947a3f1d5ca453841ac437f6145fe1dbb48c38e9cf7d443ac97ee8728423b662e2c46f461c8fda61accb33afb0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aaaa37d77fdfa2360891f2ca57abab1a79dc928594fde17804e885c60b3b86a9811227cc685cf7396a901d83873b6f0d184030bcc9d79e2ec1f2d7abaf615f88c971396728f0e455736c4d95b5ab40643007ca1d241cf63d1ed410;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h118e2fd81260bcf068459906c8646f364244dafffb82ecf1b5f5cc251421b78b605b0da1e2928af46eb974cd8736c41fe9e8a516db5097a580aae2a1bc4bdc4cca7a2ba5087cc860907d02203f7d54e742c71c57245034a8ce62746;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h42112f724db039858180f0c28ae5364ce18e493e430aabbaad13a653947b33ab728b43ebfad4e6a1eea358f1f6b1eb1dc8a9a6529a96b13433b0907204192b26234f7c485b2174ff5617bce36a38de2a618f58a701f4629992c451;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hec5e29e637e0b87bcf50dcf84eddb2cbff67148eab08ee79d1851ad560a96e2f4f11f02d5a401c01ba413f234ea2c508a95344b9fbce89769ab8528cc8b67668e6839e23fa08ebfdc664615cb46d0d149f6d2ec30c11a96a100066;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8c56e84c32d3897b7bf624a0930abc5eff89205fcabb11025e6168a9ba5356cf99076e4a22d71d080a3454e041db4447336340f27ecb19eb7922a2bc1d54730dc5aca08a30507af4037a5303bec78d629a1ed18d654533dd27d652;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18cf1123cb941d8675cbeeeea3a9c0dca588e76ae970312570a751b40f5d35d754756851ae5a8f419ba9e1706578d7840691f96aa132e3dc0a361f0f11efd88a5895e3738a398ad5063905838c7544b964f27407e62156ccef7d44d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9886fe40f01d4822804d16a6558ece998c0807d0f7925dc26d0c8843038b721d797ecd29d74a7db11034a35195c1a8e840ada28bde99951c8ba9259b3e03ebf4b66c151c866db3b5494b41d672a7d5843db96324b5ca27a1f5bf9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a63494adf54a96f35438935a9d485b39da0ac3c389908e1c1b59f89a15625fd1ccd61dc40c051da78335f4d1ef3a1ca08040cdc0a4624428bb6816cae6bc2631818236da793e4526d64069d87ffdbb5744d7c312ca3a3878be293d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcaeddcba125c179b1072baa6927939e6804b68d81352587a79aa6d0e6e5519c4e73095a5cde22685ee83e0532a9d0a10a743672f73ff72cc96882f8357205d7e1697f5ac372b2fdef6578073634f677b8b77ae8418e14f0f0df0f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e09913ca8c66177da80c615c2b1d495d9695ee396dd87447cac837dfa33820edd4f7071697e16f10ccec94c56f6f21b6537277fdc096a805cda2dbffd7d82ce5350b3cf37213b652e47642b6e172d90e5ca341a3a6b160379494b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f3b4f687f647bdc6b0b2855b142d65dd2cb940881ad5e705ed671188415ba925539f3eeb2bcfca37f1fba4c020b370ee543f75f13b86726f4ced4cac2656b038f85de37b99a4c0edbf8f466df81fa16743cc67dab47ef101fb9d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb78ba4d63f6217a666c6529fbe823a8e1f097f3fd165d5a4516aff31b1dc17af40cbe5741e918fc8f016b15cb97a1ec5b4b5961595fe5978838c8000b0b921fddfe816467b50d28c7cd73eb9f03cf3774b4b7f9287091d1f58308f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16ceec24af674f34672dfb05a4fd26f854fa63e3a9461b6943bfaa783c046fbde187fb8b496afe02ace8a992c2de6fb4293bc56a9b1fa3ff1103814f73907ae98d8ae3b32fd7544edc5eee098f08f05603b3778eef6fe560e5c1fd0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c48ad866d844026523f968d3b92f0e0dfc99c2925b73e0c203b7991a9c53e98c416315b9ed2ee2da03ce5ed07ab9b94cefd35015b5650f12d8a4c16a69dac80632674a80204b1b83d0160891fc5f353f52f44609f4843d9f1e7913;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7885ee51da83cfc85cfffdf724fe7b78f4f6b0194317e81be3e8d0c0fdeecf32435192735163cd246e05e265a158b3eb7a9e62538c814c1a7a1ebe39bf3bb329dc6fb5e7cb76fd44cc4dfd5ea0d5552a436f97d4a1bcad26787b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3df1234d3c6308986a4d273600aa3cd0cc43e438d13a2fd8ea3037fef295179b133f7c162344b6ebe3fb87afffdff23cb79ab2b12002cf4160f725a92671c005de6fbe839782898152a6e438cfcd35ac2298f984c208b6872aa2fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf8a2820c3b3e80245e08e2932aa61c4a5681b7054ab1f8c2b9b9fc2779b461c1ed232973f78e3367373edf4864af0e27ea460a8f8e56c356180c1c77e739e8afcb44b1f057ec9a8f4a659d62011832c7913a2748a10369858ad15;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf9d66c9f424d30898fa1984b1bec82806e80b1628c4d2d6afa993665cd987b0d4554c938e554b823224fc4cb0bba064920a5d46255d7a3087a9c53c8db2044ceb4a8320591830e3aa8cd74d9a61920058e830da8d427ee5bf579dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he2aa28f0e875b2281a07b9054c944240a6c68866ad532f3692468000ab910fd02b6fa3bbcfc54b2faf8b45b6a92ccc7a90fe02d1d6211c5d69aa682542357c7c1fe2df31ba85279013d506fb57c960a03cf458a3684ab111e13b85;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1db9506cc26e56465f5eaf7ef3f24f6e0e044e926f684f41ddef3c7d9a5b76bcb52ac0cc0c7e5bf5725a38528bbfa9cead0b3362ddff6102891cb9f08442182121d510ca3882e8710ea26a1e87968af40cdc692fb0465bccfdae3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16afc65f61b23a2345e380da014165ab647be882335eed0749a4b064a3a5bba70176514e31fd09dcba5878397ab313d343160b3f506d2d7c7297f82a0f25fd922070bb708039c28da55c40b56d242587627366ff7b8c47c30c6e1d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5cf2a0cfb69f4f64f629792f2347bd5edd112bc3659bc9f8b847b3034dd1cc770e079f9c1ad9334cfc1bf919e698aecd157e31318d2f8a91cb9806ea29ea0db01b96430dbf862a2c6d1a05863b0b36efddddf0dd0621b9ae89e28a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1125c961206ac188a254dbb869526711474fa7a2598de70668aadb76d2279256f5466415a0ba08532131848efcc3060688376b2d16e6dd2e1b501c5ffbbbf08645b77477926c9a76551138967eb062e825893e7dc7ff75adf174d8b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd854b86951bc62fb500d680916c6e492326d64fe38718ce79ceffd92139fb14ca411c9c7c9552d1fbbc03e0e033858e224f9755c821851f99355c74cf50a5b00fb136d726e71970309d72b2eea791d8206390ee76a6d3ea3caecc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3db72d3973f8bfbab7e3baad1f4fcb948e613d8de8810e69d17a1f79e634472ac645a3ac9865b1731b003e0b31667b71b1fa8ec796f08811ad38898e0cab047a5628fa2cca52e0fa5ece36bc3e3faab1f6dc665caaebe5a75efcf0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc74336960a27ec7d59ea24945aff3b920ff6159f5b01f8cf70a295c3e2b7d8e04c63360278f2f57762d1df0db34eb7515edfe873ac6e146fe71095b0ca4a1c980feb15f45598690ddcfab7f0c9d9512f79c8b08d21da815812b897;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14216434a8bffe991e88219aca021e24c59ac44f221070d2fe9ae595e83549fb7c90626eabf77d2f3cf1fcb7976d7d6eb240cb049efbaf994dc36915cced2d6d27b0a29a510a4669fe8c79253a82b82cd8bf7b443321727582e01cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h628b96e03a1f568f51306a611898fbaeb4f1324794dd46f6920472b91b0c1c1a2662b2420c5f39c778455d65ac33aefade4439997807601a7ef1d8078ac3ef4a88819f34abec061887f9f90eaace1b547223223b5096014b8b45e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12bcefffa8b1815e20c2ce6e031b2b505e492a636c556281e61850ae38d1fc8f12815eed48aa59ac19d84ede160005ac1e4b07678343d4377ddef0e155310d9e72c3b8e52a64ecad45c3b5be43692926fdab28859eb7feac62f7ee7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13d93b5c27ff55d5a2ec022aeb7c93cee204b638846ac44127b5ff134428ec3369de26646868ffb29755588f9c6cde55d6988ca34b5e0caf4dca7466a008076b17178dd064367d96c32b122bf4a64adb17d934922e833586bfc0872;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f85fd716c0c4d1b23892c34d37dfa270b4d69772d395cca358aa209fa692b14a2ca8040fa7e8b0744d2f38d2e2d9e17aeecf171592e12ea60ca4a20878644e3d6809aa24ed2c81a16290924c93d7ede5f8ac8a338346c0cda854e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7cbbdc3c9b56950ce58d990c71aecdc933aa571db9cdd0a8d36b164f2ab9e0eec933c45df791289e212917919396d5cce2cfcae11c0272955eed81848bcba0423c7e3bc01b54327b07137d660d1d73292c89891e1f52985510ce4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4699345fb0fb90fda293ce309d920786838760fbe570170165266a8a35434915b3eeaded4a63b530920fbd308877b67fbc2c8b6b60135e678e82e9ebb4a79de92ca2f6ff92599b31f6f4d77258d7adc4322a455f61047f2e79165b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1debcabec717c44a7e4058529d76d84f277a21e132a63ef1520b52836429b9a3e0dffbec187d084348da3e30a55145ad5dee8d44d5a70c3382dae220cb94d446f8182dfa6dfbd2349fb8b98da7cac575a74350fc7a8217cac3e3e87;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c65052f6d71df101cd03d09640d4e9d1758419dd8c973590b2d54e30e097fb1a1ef4a49e3f1b26af7d35b4c843bb22096823d2a61d7232b59ac371cc9d677d0f60a02bbea65433211bacb112a57eb3b45da5af22380c714ff3f2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h100ac98b6651bd4674d32677a44e337eea2dd7a363367f66e3221d534ce483c89fc2e1f4743d514f8ba93aba2d9d53cc197cc527322f4e649082dcde755b41805da305ee61cf100a7e85f7f65eb55b268fa5246ac7d108bb7fef5e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f849359892666bab7e0521143c85d04a62eb18f41b205e1d5882b03f022f78df4cdf99905535a5f5537bed7e9c9f9483f8ebed479294df0254d03320bf07312967f288b88e9ccad58b40661bd0fe6bec6cc1cdc3d60266b698044;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1468b5ad95a9dfb1fbdf6c6a1392e52b1a09abcabe3f6d5dbb4a0f4e538729beb24dc2b73b086422d4f672f494187ae7c6d7afe3d68fa68fc26a90b6c614b2ae9928455214165e1acf1e90c7da140dc150ff52df29aab05de4279ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f8cd3d71b99de79c632b124282f47d29719106aea2daa48e4a02b9953f2970cfa3e9500b2aa482ce3177463daf40b6dffe673791efd25a0dd63520305f310d3cf47758354310b922f51a056fa54e6de6f0409fb11d1efcb4ccb476;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h990a07d21f564bbe2b3e3d515b05ca1ad403c60e19916e1439cdba534073ffc11c3a39b325b5657db8fbaa7105f9f4e716bb12c0919b79589682a296cd5364465a964a65d1693e54c09823b5c45c469cf2c11937f1d86c94189c9f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h719b71dd8be9ce64ddc0bd266bc8b80c3b65235a969a5687876d058014225b7b587d500678e2bb34e628654e1ed8a522aa71700dd7fc0373cbe6eef937fef5efa1f9792565bcccad26ad5ca65d4396388834191d035a4c3a2f892b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f3a7ed8d13a2d2ead8987c1e30f04d68d09a83d211f8eec541a7647d430aee86272a2fcb240f28a2025a3e4d35b38fd3e53680a06e1c2a49b022f85d57c4f9178a7a1d0223bbeb128ea3b2346dc546fa03fe26b72ab5ce0805c91e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13c5d6c8aa1d42c0f1c97de0fa2ae95ed425222a3ce8dd9a8d526a36b88837971d8d715e7366d6aa5381c005c4201c23b82d5f3c85a5b698be12fb6770dfda06bb12bf1d4d4a1dcf39098e6a09862045d982d8f9f0044ebd17eab98;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc20079072281c2dd6377e4b1cae95e3d51626aa4013f37681f7338db21249ec82a70b38c44b6f2cb80cf27c6c044f39c123eb2b6583a415093ded506fee1052fbc164ed0d577636328ec258c3077a24ae59c8bebf6ce6b2d0332b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf7e25a170ac20bfd5eb0e7fc5a825353f92db0ac4a8a0363561db1133d0ea137fd000cdbbeda2cf71761e8dbf8c4ebe7020c4292880836c0630a9d90970ac4845fb707e63f14800575dfa7350bafad365e75e748b5e7b307c3b4a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h282fa39ac019e81cf1f39698d2cc333831936312edbb4f675a54ebece79ccae1c40e72d5c9b7d5661291594b1bff54f101b1f7803a7c05baef698e7399dff2cb5772da6b4f9503bb33aa9dee560939dee54692e491e0d7f0b4f36d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e7e3fab7e7e4aff1dc3fa4fe26a3f016055f4808bc801d56b01aa6bb4473d95b914f7f94f68d1fff6af47d441a29082bca82598809e210be607fd98e64e897f2919df69a01e6af1513cb5c65cf1786025b919ab8c14bf50b259d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h89c6ba7b5031d20282e0745d200b5bd641163c9749d5661818c88847fbad2f617fca498693e76e3d7dc0b70c9389f2894c766469c459686322b866b39d9c7fef26e25aa8b5b4ea2d25bbf9e2de6cf6ef1ea0de91340680025cc473;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11675feb4afb88b3153e1256e38f7d4c7cddfc1b0a015c247120e4c961bf8d2e4fdc4acc5bfc0e89953b7821ea780f0c07470f45e356284054bd25b83ed8ee46f37fed2055edcfe32ea6656aa6fdc9e35857f0c0212d4d1b5c6eef4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13aac425af365503c620f351e2c88bc0d94aa094919092662ef25c93494a4c486f899774f61255c513b34f2963ab930840766c8f071fc411c1aeffa7937ad3b5de4ab4da916af6bdc9166deace5abba32c6f736b21fdcce2b4bb045;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1553ab435bdeed31a39bbeeb292b07d07837b90cd03262dbc74d943a8639f41b5617689baaf7cce6163dee4ed83fd5d2cf1c1ee8495ff75d69acad3d169ad3547f0952916f0384929a9b5fddff4291f52ade1634061d51acf5775cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h465646ee044804e669bf78e4595120fdbeb0539f16b0a56bff9eaea03b894c5c2407b2f4b7ad59a8098ba8ede52d79f4087bb79cc5e480746f13d524c16a3f2f6ed3a143f10d7e27e369ae299163e335568c952a504387de7231b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he5e7c4fcd6af4b5c08df33bb84e52d3e7d357c3fec2e305133a5891276b995f50fd244fd5c8368d19de065babffe1ce1e7466d3cd0955536e0585c1159efe63258b1712b742336a07d7ae96bc6c1ef89490b543d42dc31aa323b65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2fc664a74cfabb479ae1254c7d506868b1a59ac63480c5d49c3ee3f3ae75347f79043f8602b7228ed0aae80ccab4f3e2d4cd85a72c512be8dd18540292638648518b6472239d4b0911ddaa0abba1e8a4dff2eb929942744b186c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfd78e32b00d7012867e37da5a7e511173eeedba184005a4c02bab1a8194412bda257cc1789ce7e01501bc03ffd94301822c0229d6bbb02844eee438245d262ccba3038ba4fa3114f3e964a03952c43d219d52e83ff55822cdcd8f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h199379426ca740b4cfa6fd3aaea35538ba42bf6a8d0b0477df0a6534172fa884541a5d11b3af4693ba32ca3fd306d642ec2af3e4867379d6582612bba46a828ef01726ac564d83e16f5deb6da7bdef2b8f323e6b880b367ac9a98c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e9c79765ef45acff3539b7f3d352a4b332d4e3c2defea30158e93e734076ffc762a8ebce5bd6e58819320b79d905d12b6874e56b7710db315cc62f0aadd60ce09d6b73f404ccd82aecc7e254a1267d346aec63c19ab36cd10ca787;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3ee1e73d7233f47f2bc5d7bbaaf7a847023517a991d1f8a78ca72585c2dee374c8a3c5da72174a4b2fddb429b57ce603c7809cfc42c2cacdfe444ff4e7372b735e99bd72deb3686e51d9a0acdff3854ad0c96b6db5f40f5085206d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15ee1be64072596e631bac0f3ff5469f8379b9c52802758364f1ea9c1e5e270bb53b8c7a13eb05b1ace5bfdd54f6d8173d9407ce38ee13081ea7ef7831ad0c01845ac68368da4c964bd000b6313e107e4376236b3d84af6e3f1dcdb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1250c0298d8daaae3ab3f2e9c344dd2a67f9c8cea7b80f38cda6421a77b6618864504706cf7402b3c569d7ff3567846583032b514889578f0c628cb25a9d61f962b75c246c013ef43270ca3a67eceb5be72d4e76bb8142dbe253d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h157f528c7e355011b46e330ed281c5710d3bcb43fd7fee372afcedfc65b8f50d015448f01edce690877c4b5ef51817835597509e9111a22a63c93266bf0f9ee7229c6330bf6da94c84a3b771aee07edc7fbc0f84ecd2785fc7833ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1471abbe81788a314bbe7b5bc1414ad1bda491258d4e1990834f369098f041b083d15ce33d99ab61592f71f678abe3eb3885f9b6517507a3516334012c8875cdf8e52706de6534a9ca347f0a12268c9ea60cca3d9c25ba9a8418944;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda8bbbad7c16df46d5d8da3dcbfc6542da013e3ffae67ee6360024e5b52a120618fd9871d56211a5eb978f5e2edd8b180977c78246d6406bd7dfe2a780235c35756cf809d0d692c2f1e1566500854c6e6277328bded94ab1af89d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h21a4d820471dc0469761f569a54f943ed91c7c21ba5a173a0d6d09517bc0d78bb8e75ef17789104e2acabe9de0d7c74978f57490b42fb4b10e06b451d22b18d2d0ca17097d58a14bce63dc276ccd3ed535a352a21a4f918fbda8be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h172752f3f8abdd6d62b698018d78c766fd4a5e545a7ced275ec6704781e76be757d5a8b9cf391f79d280a4c7e43069f00b7d84064bff02319496bcb73d95f1f576270f25bc7b143a5a7f4527641fecd774110abc9723635742bb6ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18bb4c8063a396f6b2ea4b17be17a5c51b5093e54b076e7795d334f521e4136e06ce1e4bad10b0234d1b812d05fac0fdd8b87d35dce5a7a1330ef0b9eb22e13518d8d62daf2b06ec318b38e5b29cfb4824822677f2ba4598e513842;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e54a3a557e8ad2bf68dd850fe507cd4ed854b3dd908a1d9ecfa4ffb1c01fb938cc3f2773b1daf7240fe8b47a6dff3923d46c1bed594996b0f949e0a16f7f3d1b16dd65e0559f3d1633840768cee145b3a26f1207c5ec0cb59f97e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hadeb8ce82b28c31fe4d2aecd038103e15f92acb62f148807f55e52201cf8107977631b0dcd60bf30f5a0a277b9fe69ee1ecb19b9b4cd7e803613bdd84162328a02ff79bd1a66984dcbc1d26f64876a75d0646766a3f786ec15a460;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb63d5293a9f601b2eeae692d90158f11659e30534f6bdbdafd60ab6cd3826a9a4cbf2480ba57f7efe6b278c8bd09b75b1438ed6033fbc0476d99483fc8755440f7ee6318a07a4f76b7711b84b53a5a6cba6c902141be50f0e5f6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h394752130bfb417b996e746413c4b46eb0636e5b96b7157a89609c89758c5e7269195ef282dddc417a69f9cd855dd768ef75687385d836cddb0e0ce1de239e75d372fd25f7ee3f48af9df3f84d50d32bfc9f750b94c26aa85f36cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1398d5afdb32fe3e97714098c4fde3117fb9fd583bb2f37a65be308599137833e0ac8a388f2579b381254a40e715e03cced68e4ff71a5e465d7a6340904d49affc5967a5239e6306061d22b8083a741344ce192f2bf706b709a0b69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d0d48d11c6a09774016091a7e50bd5676e885719c0296ca8876d5987e3e7fecead177dbe4ebce937b3bba17ee3bfa87ee945a8bd5308a3d9529878de5e3aba27f29673e7d06a56399395ca5b1fbf622e3d7e365b33141c4b7df02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11c1d70e2ff174a457174828617539ca0afcbe62011df20e9fa5d2b3ed20f791f446a5e67055b25699ff68459dc28c8bdff3ad3964bd083b35b10132d1157891b89358d3c40c209dacba9377e300a111fc9871257e30a80504bd20e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd7342154139109afc8a1a0db1e756bd1464ed797dc9e24014bc3cd907c70446d1a717fa80b4f0f5046796359e81de0e92eabd06049f35636a7670dc62d2bafcb090f9451c52d14070db152c722c876d6e8b72317c0a40152027f19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6ff6614492c4920a7377ce9fd15c91e7c4fb43f03fa9e31ae322ee6efc40ac1fba98449a19c4dc71660fbfd161cb1771d279260605a854849f4a13505d835fa07fbbab2b830f6a62c2d34214159dfad9087fdf4eb66c8de83e1a0d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c3803d13a1ebab4dfe2d39e2a2b495cb3b3837794012b1c4e04d642a7db2431c00a8334ba650c5494ab5e81663a2d2a578b3da56b68620d89dce7bed88211a30ace5fd240d1e96542390f80782593374a8479e1cb4d5ca3be4543e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c0b5b78a2cf30d8b9a48f0b2a9479a08bdfb7217d26cbfd4aeca478dacd6e6ccc214458c38165bc0effcd404b258b98abc3a0672c590cf0915f6cbbf0e81ead4801b871505a1f0072d7aacd6ddaff5564d64d2585b80e1a88a264;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d18fedbce6fa863513a00533a9f3b70cc93b68a08a44a334a117d8653de6dd28855488d3799552ccc22c29204a961ba4cb0357f924ad5dfe2b16da01ebcb5e4c9ef8e761d21622a823a5fa56bcf377cdb846312c8970d95cd92f3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf4b828af1c3db1e3b5fddc73913bae64d5b3e4dd5840df189e5dad6d28e1fa3089f559dcd14e3f257425dba7dd1da83eb36ef183beb231ac6e9ea76cfbfd2bda016fd938c2d5275be217ebc405378029a220af6d0871b1b6ecf432;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1526fd0ee812ae7b7e1b2024c2568f573d1c8af7733cf4b68834edf858376b062711512756a4b353a5efb726e4ce65bb5947c392594f2c6d029709803f4b77574ea696bb64045ec9f476ceb28962be249240fbfdfd0d25ad2385fdd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7e0b432b2fee3142004c7e467d1c245bc116f435d88d0dc4a9a9d10ead8646b770d7b69860639730492a4acc1d4552a8b1a744f252cd2ab9f7af4b1edf67027382246d89ad9fcad3493319f5e8e179a8a7ad3c4bedf7a49db9644;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1113492c45d9ed00cdd054a7fc86daf9209194dc54d698d2bcbb7f03e26fa2ba5de63cc3b61ba88d8345ac9abfa1640ddf2843a086b39f61a9f0d2d42d5fdd89c1aa52f37e991d01816d50e8a60870ef0cd06844c84f121d0e238f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36d6320dede8479fe5c1fd0be1e08df64d7a39e7d64d0803f4dfcb9cb304959eee2bc8f10f82906f23847dc68d27ae7385e2b74a3f84a7104f0fbd2c7f0e2766fefb6d98d22d994aed1cc03ae66e1a73ab7eeb4e49021f4fb209b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1416c9b964d6540832ff2752edf447d174028534c5ff0dce65824502a1c8222b6e1343f28b3b04ebb6603be43ccc560801931a7b7edb8abc016bbf58a369317bc45640c9abc7ab52c3d867c0e2fe54cbfa6c5e151303cdc33325861;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e370213357b0c40e3b3a0bb27185ebe6ab7103364d062d5b52a6745a7634490555b577df0702393ce68507d4c3bc1fc26bc519ba8f785cde017bb29c2df14ba3a6e8ef55ff596dbc369b351ab3de2b564e42f6c218dfdfa5c0ccbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h89dcad587dca1017de63071412734b0ea0a32103427d8600aceb481a30762f80c7b20a3b6633810032cdefb5398847ba7fae7d4b81c36ddd768330bf917543e417bda8e58f091337b77108083811872faf1a1015984453fc59a581;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he2db41a86b725eae4b9f3c1377e30293fc203e69484c9b5d1fb22231ce7e72ee98ec719fcc98035882b9df8befee69cbac1e2df280b6e8f8e457f42b5a5a1cae55cca6404f3a3883c8e17a431ef3f4dd43f002452440c54a2cdced;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136484f03de4526a52fc7b7fb8052fe7ad0ef3cc62120b8a153ae3aa7de88d78b8a0ae93165979633727e4a9b8069c9d00b475801ce5dca3dae855aed826afe6cb469cd8bcb32061a2f8702031254c40f5d405128cd781ef66e1ddc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb882c06140c618b5bf434e9f811b06293b68d311302cb7fe8685c3bb29cfd79b73ea4df8b0adb546ace10169f753999fe23ab5663996b9ca663412f18bc3bb9acea8b1fc48f5faadc9d1b3eb0b06033cd5f033c0cd7d83e706d5f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he4e432300af9c970e60aab9bda6f454ecc35d5d73652068cbfb566870e9a370251cb3c79a9bf8b56360dc404af222500dd66f7683007404dada5e8597bd22f3904f970a787e89e3551029fa3dbc5828e4de2e005224a2e80cffd1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14c1bc7b98d2f23af21e52a917c3b3afcb0f27bcc4114781e7ab7b5b3b862c83eb86e29ed4f3ff79c2509d0d24224100affab15a764f2bca897bd68e40dfc3b62059276535f49ba8cc26535f6d52442a8d7c2e2b51e468d0d631165;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c354dac1ec60f55ef7c0f3ff3ab0f0866052bd3735b5e566e9c21c6ce08f3590a8b3e054d89ab04c8b272d498c441ab47cc19ded979918f3bc96e5905ca82d4809a7008a5ce5ba810383b2fb29bd21072af6de8d2df1c4cebd3d7e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbdff0830c236e28f80a1f395fd18957a12e9a5fb60640fb36461cff9eab6e5483b500500eabd353300c568591d8cfa7a801f9f8467288f4d20b72adf5479bde39382d829d653f800e25ac52314fcdbe6063552fb0a8ca07223dd13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76e186cdf437ea85a0a1b8c90cecac38afe5ae1473eb134d44427831ac7876a1d0a7ddb87391c606040f32837253a0088d18d1e250658cf94d720f3576cb3243d64ef7f9c65bef132125a560b6e0144f5cc2f63a2b4ff73fac6bb9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17cdf6f3ae1287ee8f28a04af8c4c4f05b650c7cc613501a72eb067ea0c75e12a789700504599ba3adce89bf76524713835746670ca355573c1ab6525eb69c5b33a772c5d8cd5c9da9296f924980ff8ee499dcc7b307f412c12ba2f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db5f9d999c8c910d070d8abc7eb46980814127c8ec4eb5738b112e2335796c83ac27bf80933a03f7d7a18d76748b00fa4ddae20d32631e706ef05e0769f703eed572221922171744cb9d76bfdee3b3567a96c9eabae182354479dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3ae3c87ea6fe21ca0995b84aad6fe6897ffd8d62dedffae34bdc5b27f980b43974ecc9bbd8bf0db8cf0117f8306b3def6172cfbc5bcfb331eb2a6f6e677f4ba77714fa34cf3bf4f13e05019487621df69990dcd6024f5d24fe9d53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h55dd625ae7447613fdc564bf9f3df6410a57cb987d8afeab7847b301babc2e848ce779af3da3d21dc7fbdeda6c5a1cec44ed17eb881661a4220ab5f8ffd1d0c2b506a7241652a6009f9e65bef1d8d402cadc4f10ba1bc15ca7b8e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15c9dea46c25ca33c5c712b6c219e5f9ccd83e0c7c474fa10e4104ec919de06d751686110f9afbe1f65522c902a57be7a5f46dd4fde80e0283f2caf3716ca6fc41be49ce24dabba6f55c526d8e1fd044d0d5cea9185e76917336c7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha6de62b8a0f728578e376fdf934dd7946bcc114c12bdb328facbda9d588fab08938e333b222e88efaae41feb8e955193ba6120ef7ba8251823458afdf90230c2083002e5d9194c5bf5691db646d81757065e21353ee676b47d5f7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16f507e42550f4c742ddfb2b1d1ced36d8cb8dc3160147360aed468a4c86a5bca4bb9017c9470424c5837d64a89374e100616e3da11b6f34e11d56cbd9fb9f714ab913fced4268b03af3660c5feba172dfed3005691c508931b8962;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5d385abca5eaf1eb6db66d6ec6810c4e92ff5d4b6985719c3abf9e614a8d2cf38210d5ac78a81a37167c7e7bad55f945d2e3f918eb58c41cba9909182acb2559a484b744d77ea4015cb0b8e5299cfec9a4cc2565a641eeff546c83;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h78f8a2914348d9a0ee40939b10598939b162a62b56c3a937573e679756659b5dca0c47d10e0ea8fa61c6db5795441b2f8005c05d2a3c27c4f92fb8fcca008a052314914e47c569ef02d934b73d83388ecf5e27cd2f6065216e8375;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16fe46530e1983b346571b9b77b98b8a431514e9f2479bdb9ba7d5fa4f5de96892d6972a3ffb9cd322b946b2c28f8f723841775baac313170170f064a6ffb0b7da129e891cbfaf2caa2c28338114bb838a2b6d85a75c1f99e2d4f56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h556f47ab8d6629a95dec3974d9d0692487b9cd20159b407b77404c1821a0c3220d5a5eb2968cb67502dfb6ce2a47a7fc6465cbe48ce246e673a0c177773d3454d4084258af04a8d12de1c23684336ff6c33da7afb97a7670bf9fbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcab9aea4b01c651f75285dee6cac115e13f9fe49ff418eb308b8202936a795fd00415713394e69efc112a7e2e03126a0dd0d2ff9921a00dfb8f1c3f144c71c3f414eeab13a0ff2e0285f11fd509ff7c8e6299e71fe574d48dc9895;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdac672c24bb743d465369dd973806ff58f741dcb4c48603aec85c4a1ababee0a9907ec4cb49251023a593f54f3013abca4d5a869f66d3ebb93b22809eb861bf7027d3e9301f2b284f9f21cac0d85b5b89a4c43062a765bf1b967e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ba8f03d06052496b0c31426673353897e909a718aaa48529f27aa5ffc92d1c82a537056bec98be8b6ed36c48fc6386a4bfa0ea2a33a838f0a44256ed86620e8d34349f2b0c44193c44307959240b2700cdf06282237ac4943d7758;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7808b1f0d5f388289dd632d3129d768811a382298d3aad99f510de458ea32a8e589249097336cfbab60b1ae082392bbc8478869fc23c4c3aac15da34d550ae417ed8ba227739139c27eeac4b6ecac325de036849d2c2887da5568;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104bd54c4d3ea51074dbde50f5a3e1bd743d91af431375ee97a49d103ee1e6b33592754fce833005a86a0cf52171e8075e86944dfa6dcd77799fd7ce0fc2e50b764c253d6f42ca54be12f0beeb99c7ab9616af7759b2b0de110df1b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15cd55cc96973f972299b127bb61e44ed782cded003595505f931c238bb21c14297978949eea41c64283419610e58ccf39deedb5e1680954d1771747b1d769f1c22dde98ac949848211076c71215326ff87128e1858e6a1ece2cf86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18752804e616d9cfcca1b41fbc79dbce6485ec57ced1171a98764c8b08e7071305adac09e7d3dc39e53de63b76a5d1beb0b689af98857ae0387aa2278f372700fb337b65ea14e4ef92e96105cf3aebbba8ee479399d3749ac157d30;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12937e91d3e22aba92b76c02ba3ae3bd5aa4df151d5a91e875ce2d3f429bf7404d97760350eca2344504339869d21fc6bf68e6f3539defb899af95c661f384782abba6342ada828942c82ce8a69911b474ebefae86b396de5b51053;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1749eb6d49c6c44568bda55ba8d71b189633f362b85920c4341d14ea32680f918748b39c9a98e966e6727d7daa0f02a2700d4228b9ed5613be98179b0c266e99fcc5a583b4ce4e25011e35bff2bfc4a734f9848045052a63a824027;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4ff31a20d1305aa58068d7f246b3c08d1374ad53716a02ab1ee28adab1f0f6994fc999b9ab61c8387eb44d20f1bf08281ce9d9801cd373d6877692cb965a847e52a2a2b21bca5d1ba1a33e3edfc0f3f77204ac45d31d086bdca476;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2933087b9cab97dd3d9acfa921a63fe33e1fb791db634290eda400b7fe558388d01fa1f76dc1a88df97f2e4f87da1c9befb69294b9c9ef33abda10e0a3b85b704d7c66fa880fa0a0393d3b94fd39013bff1b82418f401231c82a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc8ac10ed395729e742afa5549de22b6eac6a4d40efb8df8f66f3f923e99e248aa0cb648270c8d1c9bb5569c90209ffba72e5a0825b2b8832f8e1c13b17e19ccb7c53113dabab30892d602297f52e2733a998d28b6622c05b83405a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h58b1106ce6a2484a2a178ae62b958bd14ac0522df243e34e38cd85de62c3653975d85968959e4e841ce9e240dd9ecf4e38d7c47e29063a51741b5ed4dee7eea1ba2e35c1c59255472a6eece61ed6dd09e3b39537a1b749597765fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h193635534b59943a3c3b367a0007517f9d2dd85b40ab8aa48dede2e07a8fe75fd6564e38c7162925c606688f3699069e0549f02ea73685d2d6bbe8ec151ad5c8589b5eab5412253c2cb15dad1490c2692ce86b150f512976b15cf0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1536bbd333a0a238e0ec68afa4eea2f4e8b918057fdfb006cb4e43b99668d6b0f6b8ee72865e65987336591c09d856a8745027f91cc16825dce093c0338d30d6c5d5f133dace8fb286d2d390ad9d6cb5cf902a53ac28ab7d1885;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f644555498c980b42fe89a864d3296072b25c43aa8e039d7da8d81a9e06d5eb3573d638f22c41dfad9e3922e56ac0fe3272afccfc63cf1a5437d470a5dd1cd3b9bdbe7cb603c9f3a85b137a8c481f473d4e5b0c537e17af305e48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1acc2b2b3d387899cc9d4b47cee3a073217a47ab13d0ba481d666f8179f035eeb71457b5c1ffbf47f4cb343f367b85e98ef5591df58c8057a8ec79e8be4db2e4632676415355ce90059080f00cedafe42a582150cea31c7d673ccf6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19f23be5a2cc306a5b4a13ed3badc7fd11ce29195afb23527b9d99b1a5fbdda75c6dc5b217c625f98a7c906aeaccd382609de4bfe537e8597dc77553739bc6b27f6f2b091c356a4e2474168e6c8a92c89d86137bbf4a33a4cf1738f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd1e64604cbe180e9adf189f800984457261bb6644fe44dd41bca58203c2762f3dbbc421f9488b59f09be82a067541db30bcd5bff3eef0275f90f403e0c44cb1351c536e4dd9204e1f42d8a451848c1543fc052f6ab8e31d1162eb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c83b0f8a4e358bce443032159110758409c533d6a54d3c2753808e883b92685ef88e3256d3532ed5f2f311a5abc36dc5678e642a9035831c6db2a40e40718788d970bdd36b704d908aff3711cba4fd9af7899df573bbe825d6a485;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17647e2249714dd72bb1800a4f9db9000000633a11f25c030af091fda2594eb9c9f427b684ef8dc9aa9c2c583c2b2011400e87711639a3f6f085d49069b3a809dc61a9b4358ba483eb288a5c5b03138e847b0939b827b6b3ca9b013;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h30250e868e84fa9d97bbf244cf94628424014f14cd51df2d1c9834f223d1ee32869ba91234b55cae70fe188b4f47636fd085a02687d3274de4fd876182c661874c6260c4772f7617b35ed4691e1d71b0c152b2fc09f6c00eeb2d26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10df399a6182110bea1dd898b14a70d89479814e859e587ba2b97ccc97eab23dd79a2bc9d8336eaa81ba3a8a939fa5f53f1d598599798e3bf19b544b52ca4ce468dfd07c48a19cf792058ed418931d8d2d62f192aa848fee8020e0f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h180be0702bc8eb92918ef66d0dbbd9e35621b5974732eba5a96245c2723c3c6635a8194f680ff9c74aff206489efb739c9c08cf72781d40045718267926ee4c3e15bc2dc55246555e79996b519fd26042e71aa5b67adeefcad07bc8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf5d0c8169b05a1225026c51071168135af2b972e9cebdc95ed5af684b39615f201c3ac5fa8ff4665f7e6b2255f3b1372a91b6af66a50025edafcc646d8e6aa3fa3665bebac282c1a3026bb94f60d8cff0039d299b343bab4487e46;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b10b64c87152094ae74cfdf7a6dde9564ff32b622e4f9cd52db41a0b90cbab4e49f13916db3a821e0b26f19999f1323fb9a7adaefb6ce4a9a78b07cda00ff691637626bbd2a5fda0949e38bd069df4f1377c67fe96f7d78bab42ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76f50d0f3c596b446ae3e08fe359bb5b6a7fd4abd76460e66106d3161d44acdd4150bfacd452f2488490e87c4421b3c28a5ae5b2ced65a4429fd4af02483cb9f2787b7010079aceed1b8ee3be75277111d12d971dae3591e00140;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h616db9f394ebb9d97dfd2495b5758492918adac845cb81b56ffab87ab83aa3361d58b6b55ab71997c43a68e0decada090320d5d517671ba0b5726f9fe5cc7494f350df1caf711c40f1bed17ad313a97036a72ed55ac687fd8292c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf92dde3862de9a1593955e2e5c507a0fc276230627631e8dd0d62ba4ca40863eaa558405823320f47e51165c8109ec678d450136008e78d8094211767d9301365ad5bc03c03024ded57e4cb74e4f34e0ada17019e0a2024530d2bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h550d7192079095768886e448077309f1f0d6e05fa43909a1db926c84812eda6447e5863cf3b27a8a47bd52fcac48fb30430fc9e41444e428d98d226a8489ae805659c9358a15f8ba65a467bb096d28eba300dbb8c04e453243c4e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f5511cccb4da203dc281d5abaea013b46f467518f34b76e9c273b00aa326333b365f814e52493d27226985d3e807271c8ea5f57b2ade3bb37fa783ef23be9bb793fbaed4f689bda8ace3716d25ba5c0cfed70efc0e95f7fd3cbff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h93c1b756a0272d2dd2ee2b663a79bb575bb17be02574553b4178f0e33219533e15e5ddb744eed91af72824ceb700551352e0022688dc454643abf8f32b5530ec87d3f8548c2c111e656bc2e16bd2f222e80d6c7c147d97f07f0c60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18c8c166b8536b4668b593bac695c43406b4f4f8c3679bdc748a597cd6d87ad0447676e75735be9843a392bbb0574bdd99a2401a8f8ff1ad865475f5e0016bc05b26b067339c84a576c3abd4575e08a57351123d2bc78fcec24b9f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb24b030f86557120de2e3d0091f67891d797884c1322770ecdfef758365076ea7f3bda4897a9922e55f2a00ad4ff6c2315c45b32a2ea88ca4e42845e7c92f5d636026210d0460945c3044b4743789bb9533aed0d538744fedd28ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11c659ff47bf27e6daad4827ddc2b97d418e2491255068c721b52a90c7f39a321d9a5cc10d45c94a0722e693addbb63a63da66e7d5e10e4e85b0332204e506f8920a0d813bdbe8b861827bc7b31a76591a60a19e41e706667a086db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he4c3a367333bc1f988199c329e852611d9e400f087a35861d8d8d3a19ac99f97b54c317485173c2a66fd8d219144b7d7f8db0bb3b48d0d145177e387f1c715c6c96c77181bd6a2c37f2c2f3571f56106d9937b7e397647fb02b089;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda57f478c84046d5ad8ad353d0b27359bb5b226738cd5899f194dc959ba24043bae3ae44c88cb6a210870b7bfe65011370cd61f85199802927a759e7d17936656920cc7f506b1b58b5e87617bf2da9a6b875385d592af99765bb2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4482a967615616b89ae91a1ff7f6eff0e18a869f2d93ae3d4f7fc3072cfe6a36248c23f4b4d866fcdc7350e5f5d86191a790b0976536e9421629d1c8d3f750ace146deed0aa8323f6b801e8993e54e8168fe264ae86d330b068c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e6d45797cdb35a3d9c5807ca4f08283be1109fed892cb467046a3b3cfa6ea937588e3cba221acb18c30765cd53d0a1807771892bcc91db26db41fce82a4e28684c6802a862b9d5d8a4897d983a6d2591305c34ad9a4f540973e4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1828dc14535954cfee2017d49380f3d37215d5f55d0b7b8f6838db4c0cdeec3d95ceae7a744beeaf0d31bc3152dbfa7de2b665bc9406fc6a9ea72ff8157722eee5e7086d7eea2d9cd28aae7c39cf01796ae322fc93d386a2baf41e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c5a296a0f4f6969a6835ff33196ec869c89a88fe93379983b3e511269e78d9b3d29758d38c2292b4ba875c78fad685030078f70360f04cf1d8890ef7bbc789d1f04a5f405693449f7c74348683a7aa630867a124effbe4c5d76c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f4a206309a46db00888842c8dac277f787b1726c3ba1a091fa4e9f538c4d3b732deea4023c56f34654a2e87d049a87e1029012660d7d1d1b3bf25647493671332100077a908d367e71aec16af28a01789e847731d646593929159f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb283aa3fd761edf90092bbb5d67f6200b62d4f6ad5b1d8058f793c9598cc307bad429f11a37aab98365105cb3eb3a638524f896e98db3438462657d625f61625e050246090972998d978b2e1c2fe41d6d6d92a74025552b48eebb0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h128221d81c2ed5bcb052931ac1e75a265ec9a85ceb1efe9d22997bd2371315f7f42dc819c97405c64d3a684c18db92b2e187bd95f5df688b4ec7c1a4d8e1fafe3c4a3320ee24a0ddc6c28e06d1fc4c8775d2f690f90848c4d81f82f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc28f72e75277d008e9cccd74489d6e66dce213bfa0854f7cb17a1e48b92e5a5764b3829339a4c0662653becd854b522e85958a136e94adae536aa5d03a5b2dfa9e80d90e1e9f690ea62004da3702b763b28d00bea9c45f2fcd4180;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4e6d94793d08b99aafa2ca44eddf407b9cca5a491b4da1376cfff6163cc86fed2b67d0366f74c88a3f917fad71425ea865b77f7d495392a1928ab1643517a8ee4f029e261c8c8ecf72610850abd90f731d4f441bf35a64440b3bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104794b6dc47012756367a4b55d79a70fdf283f7847493924c5e9c9c312ba177402e208bc181b53392e774e399a17b3b59897e0e9f2ba4a65db8f7588b8cd5b2f5210c66753b5dc6dcb46de48c6652e62c3261e9d90308e671f9dc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h983153455a8e083081494a9e84d955c12803f9e3d2f4cd859abf2383997c244d3490c27343343a490db6bf66282503febb1bfd303866d4c8cd9bddeca7adfa82dd641a9db59427167af55352e6f7db98e7d7f33831b927aac56b03;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1399cb7c0e6b5f94804067762de823a74990e592b2a959d65638b6598d5d409c1cd7a26232071b5a8937516c3ded2821254c63ebc4d535bdddf90dc158d10cb0d37adea1f6bb4f44c6314458eae7b6de9530f1ef0e56f8319f10688;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6654a0d26186c4f08bfb0e436abf14d7c7d0aecec071640674003e5394dd24eba9c4d7e186782c8549bb45b0cca54ca8de6180ab9d56e662f6df4c2867ae1573389e0da2cfcd07a6db5d40d9bb29e079ea7a14e47276a19927159e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha514d369e13c84701559b89b6c891a4c042b82df340e2fa181e7019d9acf23660a10732d5d228cac38435a0e4355df5d8172f4fcd0b98ce9510e313a5f482f8398ae2825e6ea6c73927920990cf7b32cc1c3b49eeccb31027550f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed2f388a22aed5bb915f0057a6ff3ece76f85926d0b579e6ed1de0ff31759116b147d457a5185882b2e625432a4d29d6ba75c1647d53040cfe828900f824c4c9a4902e9aa8ce5f42f55c686099fc182c31f627eb2ce61eb47c4c3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19b142fb58a2c4b15150083fca39dfed65fbef3066346c0f48b66cb7fe8137c546267539bb1cfd1acbf8879c1dc0ede109c8c9a431b697d485471c257429f31c434a35f37fd4f2b06bc3c27eb97e3a0b2673d76e8ce775d250b33e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h39f56e44d588e71bd0f890a49fae4976e2fcc26730df6a27054342c574c924041c13f6b4a2cd063eeddae7d798430790e980b00222ed3bbb615d27fff1bf9b9f5c3864644f7a10008b7d1dc3d90ff12ac5b9e8016d02d49c2c0440;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1538f9822e6a615af99e74c2929b99c86fcbc6d417017e285383d8d320a13382088836cd4eabd976e5b57f7fed0654f231d47f896d53ce3f283d477bb13417e58f41247fb939a9b49af2a216677daabee260b00e1982e2666124f30;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b334ce0eb7d0d6936552b06409cac88e0178adec0d21f69461bdbc214277b0523b05fae77140ae1413b0c36a5f35c165ca04d95d649af06ca60694122023458e42e7479c893f4e6bf372ed1bf57b7f32de7dfdaa40e1b7da4cc5e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a047a528ddb6593b6fc5ae33b81dbda64ef376330f7441b1c378381806370c1f3a2dfd1e7653569ede3369e1821f61e290b076755d87794dc8210cb1e80c7e2c357a98a1637a748cc4a09c2313407036670797cd6693118aeffcc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hef3d2e9b20d3dd3973138ba350624f8a7799ff67d300f5e587610fb0ab4c5b4049bfbfd90d8d528841daabc087075882d2982c1f6280aa48353bd26316f0df321bb5c3fb2424642ed6b8afd39094a75e49e7ae6bfd434effe09ff2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8692191926a883a36ecb41b2c7e96560807af06b41529ad7056cda20726fed256c532758cd8613b19d4f1efe032c1cf2ff5fd31d2841d198bf35ddcc16aa3eec0c30ca7a25a8117c16132111d3a63231329e38bf04eed544c89e3a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14891b748d1bba7d4da3a49127bcdb349d14a4443a7facb21c65c0181d1bb6fea0f745157810dd27de392a9840ea514a6ce3324d8b7156e87450d0ae853f798ecf157fcc6741e004c162c6d2223bc4021aee73dd90a139dff516d4f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h46c5aca95f06aa06c0cb44ed3aa8eccee28b4c018bbf583eea2c46891cc9648f34b53c0a1d91df60670d88712af4b6b532a8f09ff21d7aa98eb1c7c69ba0f5d5418ff3be43a3bf4191d5a60f0cb6afb48dff0d7a53879946e5bd3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h153c986424da833d9541fe85c53b5e76a6b6beb9c2bc9d6fb8fa2e14f642e65b6bcda3d6274453bff49892bae5ac60654e453af4470f4f0363262f7c664979e0e912b5dbb70f1aa52ae06c7d611d9d21321e671b8d3898a46919257;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d4dd70c48f7d73d14edcf6638131a5d5e0c4976a2ae10f92353f25407a7db85f7d15282e43ff5c140c918fbdb3a6962b8eb29b49bbdeeffff39ef59c6f7bacb0e781b287b2fdfb3de02042242cad3953083a11f27a461465d4e87;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h54548afd228ef6db9234702aea1b033049d2103c6579b6ededeb976120030f249d2b8afef94595a756bce13734b8e1c89f9371941cbf8d95cb75f76b10a8e9a1a2bdacba97165d29483e85d04c6a14a8fc288bd368859210111bdf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b2704ddec09e2877e178c02cc2d3eb1763562eb28306c1cf34d86ba950e4beaed0ce42d778ebf5a5ea5f467582614e3de511ebf349455a33e29ca42a6a5899d28043513ee121ea880a8c604cbd356e4a0d050dbcb0142fa3b81b9f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f7ef70be608760e574b55c106704ee520268628f00196714d4861b24feabe8adc8599a848882edc1c7aeedab302579fabd28ffff4c755a37eaad5817b4a3a4a6e79759817fc6e8489878461f03c266d18f0208bf8d540b3d49589d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h119587b0f191e710a4005e83f20aa3415a692424cde404644cc350878b1ada37ff54c01c70a68e3e562d4cade9d0f7df136e635fc6c948434e5eb2960d2f4eb16a9ba0195719ced2d2ce26638448662821a9283ba7e16387b495b0d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h125ec4cc3a4aefb2a791a5c69ce4f152e144965ed48e63b255411cddde6c303d1c2cb7aa9391ac522ed19ac1bacef5def7d03f21171740b5c23ee304a02320ba8f64492a07529f7452576a16ec4027356959b3379641cfeccecef53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14043608f63e259fde709d55abfddd190c4d58fb3bd5d7d411c846b2de0fddac48bb00b81e58c8188e9306d3344aee795a89aad500efd49ed8abf0c81d3a3870f0edb7c9df9771df2f97034f6d96e8d89ba3d7e3684e663b36278ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b0e896eec2679736f74ca2ccc962d3df3de46b617ec9370dd8059abbb884200daaa728d3b338378e55888a1a5d20c95716ba64327881324f21cfec6d51ea770097dd5c5a7a299c616af6c896dd88b4f5afe3f345bf5025e99d56e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb7a0578149f339c4f5d3805d9e5a550b508b05f437393cc6c6942863815fa4ec96fdf93dbbbbca1552c23cbffd361a3fc95b9c0f1d3a3fa13efe9186b1ca32abc8df24b9aea08c06b3e8bf4d615e613be5177d9f5f585d2e2ea42e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3f28b7f0f21e3daa319d96178ff0a3ee1a23c7ce2dc4323c0783e34312084abd32007f9ce18afdebc58c57c0ba9a14206f403ff46859de0014d7a3e1d552064863783e61b656464a1b8d726ffa122bb2ba2af08ac867bd21e6db38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1efb3a6baf2950cd3e5130b629151c2c353d8aac48230955dc7c35a2e60a178cb28dbe60299d38247e933c407d9ee59f39903496f33c2803875b049de6fcf095a71968650e431fb6fb02198802e31e785e75d833fb48d3eefa96ae8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd883b014e925e74aceabce7b4cc24e9dbd35a84ff8193f3f2476c3323cb431d0f9f50dcfb84b45e5e61e283c41e31e8eaa068011e7c947454dca481b053eaafaccfbb59c87e0c96bb68857088840163e7e2882e28c262990f488d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0036df073d5827af9a253dbad5c9879230cad2eb7f30b965ea972b781328c72940efcd2267a10fe6f88a115a9146bb5a4485c0214f5e63a1933162609354ac44866d9bd9c8a840d55399f54b616797586ec9446c0b1c9df8f85a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1be71084403329523a1c057571588bc900672283944eab72ec65f58715fe01c003258c5acc649682632f8573cf1727c5ee2362554ad8d19e4605d2c0e160cd2af699d83b76b57e00e1295a7ee3981a59875fd0ca25dab24207ab580;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h33ed9b5d5a7b06d687a6d719f8532de268b43fa6c32c78119db44ce44a8125f55a51f12c918fc2cf88ad1c20145c00109116144dd1bd8ee29cdac855493f04348be8ddb235c5bb98cf49eefc7624fbab337e7e9bb0b1e96c1d8249;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f5f5c99b1b3c2a2f23c2195cc495af4970d9c61424ade2f453c4e1e761ddbe9ec0632902cee1a096e0a6a93afd9e725c6e3da742ed2b70df72fb33fbcf611ea08b61798998fe78b3db749077f5bdbae70958af7031f0786ca5f98;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b6cb8c1d9fa5fef2c125bdf590f3c3e485c17dee79b420199d22f0506352ff88bff932ba90f0801e1f270ac07832008805dd8589696190ec9b8070a86d75d66b6975a719d58032fc441f54c7ff37446486bc828de3d7f96062d643;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h48fb9bb4164f09bc3ddd6a8ef4a5fdb816dfae910de15df52b79c1961477de9561fd4a889748b9779e20728fad8f1d2b7b0e3e27c88bbc2c9e0982c057b543bdb138b0d3bf347e8c4637209cc73fdad676fc113deb0726c95570f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b64566bd81c7eb776ca96d61edbc42faa4279c199aae2c25096fe9ce9ac89848473afb4efa371ba0ba7d0df2aa3433fda67465fb30efc146441a34d4ecf6547956dab55f60027a474eb8eed1d3af40d30c7066af30a6d3933b8df7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b391db24f5597f4c676b352c696133eeadef0eaa3410dcc38153b29cf7e5b8d84b7eec6d4c8871bf8e8f536829e2b8fdc949479737bd06e640453fa9a7bf163e119fbd7d904043ab726e61ea51ab817f512dd61bc4f952bd1ca48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd9ff87be111efb0ea856dd4d858900e908e4d2f13147071106a63dd9faf8d25b671f740d5f4ee5a365b48dcccfe611c6f636311ed3e6eab7716e0b64a0c0c06a889c2dc3effde7b70bc05eaa2d41081a270a872b30325ea24584e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h170e86ddb3c797e74ed764e04d66dd67bf531bb1837c6aa609a30e8dd1b84d63ceab619efcd020a654a7a0f9438b8c5d3bdebbe9d32f1c21cd3e7e7542597c89c50da6238bc291dc88d86b48b8bc27c55c606857f6870e063559df3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b130ffb329e498dbd3779c83c6e24133ed70c35046a45bd7d12995d29042105ca54bd63242be3dd0793eef9181378e5f50b444efb0a5d4f5c2cb6a8ffedd58421456447853c208630e0d84c588b1ddb887c971c89418f28ec90c7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9417e0cf0e7f590767d85293a80139660bcfa4cace45e775517963d9860b9cc05637d39fb95c4a569e3debf55b6e06cd96790bd5e585bf5909c4417fff09bf784baae6b33d25df9d2b36bfc99283836d43b66937e27c57ec908a38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179a24befb2bd082183ec98908e58533732458309d8a0d187c797847cd5e9d5e7fe2e213b657e6173de175a4d8cc02dd6f6102d187508e4524f990ca95a0b7dce2a1587e787bbe3210d28761336e06be5964c65e7a73ed2ca72be43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbaea294dfbbb98213bf4ec875da64a880595d2f5b7a75fcb8dfbb2c3039d3d8a42cf68ab8e8866958d833f1c4602f99dbfa3058668af684a5ceff5750b4c4fe2de483efa97fb70a574d3a42692fc71a8a629938f73edee25907ca2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18ed0ba3d821f12dba99823e88103cdcaf919f0bebd69bb23b42ff3807f1f31c61c773010dcb72ee4b0a4ecfefff7a92e3fa48c8da5e605150302b2872de13d838761a53e6d1bab15bafe8a3184c28d8e63fde1d7225a215de65ed7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7eef4cd84efcb43c80edbdfe4b711256997cdeb33cbdb5d4104a19e84614d535a20c4122bc835c4b6fe4d9d080444d746962b42b2b8892aadf0958c999c0d92ec0fd31dc053edbf3258fa977cedbe96a34b47166b7173895f10a9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a6ca5a811fe5dd19c2bf36797d4590bac8e13cb9da56c63acaef8ac67368ae498a9bfa01222ee0895641eb737a1611d683af082956cab1e32d517ae5e73120024153342d2319357438d24988a5e7e138bcdad34dc8cc39fabc0c39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h101ce475d272314c81b2715f2f69f7ad484798072e255bf3f83acf4a4eb33b2186b5f97fc7b22e7b78e3c49f82876897e40ade8cfeb3436a966e669bf47009a9678a26947541dc14000ba9388d7f90c0567e1d7db2e947eb544225a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14f474130e34bf305a0e49cc5f861e0a81ef3d168d7fd329f47b3846708a7c83494edd6579c9e1ba19554166903daa61d578d2534e8a8f3284f7731397821ffe3324e991391ddd1b00c28927876546cb326936185bdeb6b0cd9682c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b53d097a2313c7288f11b0246f37ed0b4663c559dc3db4e85c0a08c245fdc2c7ce2a9712c2cb5a87aedee72564468ae1f584de453a40c5e5602ed8318488dc265d11fb8a11d4dec642951a0bf54c2e963ae81b9055a3f4bb3a13a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h131b4827709ddd7d0c60b253184200335798a6cd5579bcffe0933df66e17d523aca7e1d936de64f4c9b9ce7558664767c60f10996c5c29f3430ad99471f2362b5a6110c4e811530fd42114526295eed6e789cb824166882ce8d4e70;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17cd619a58c0b212215649885f7c065e9c23eeb70f4520d8f5cfa8ca692d8f42065b66d585fb305fdd118e0e73b6b82866cc26f195c689468dbc671f16656f84d1e9b1b72806db1e52b04e8345ab294905076c7aa9c93ee80111dad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fdd7845e88a378eb7fdea6af18a922f2a8118e62164dadc674c95c11bac7295212a8646d5b4d2c0162eedab6637f772203455a75c653bc1240910beb49e22400f57f776e9a37c3d3c02621764ac09b2803a35b438ccd17d06da6c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1737246b772e85179c0f2774cb0d0a86d3ae7cad3edb0aefb8e19501c7828baae8f4a5acef5d6a153cae08ec4dbe11bd727e37359104b99f0b35313580dd49a96cc100b220602253f010a5279fad5f2077bcd52e61dd726c3ccfa4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2819a2edeb166263a50962ee9c081d0b0cbad586de2b38cde5445a5f77274451c052e199bc083549f904cd0e1de1a2b35051ab9fdf330f21e31eebc7e6fced62ea08a3ae57b53da9c673e1099a3c5d6daef8cf35f96e27098ff706;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1aeb82e94110bd2b20605feebbf9e4b13267d9dc0a70379a24f989a8210c89b91e64a3667b5be3559d45a919e7b3dc1418cf8bfa06e8306b0be3dcf942edfcffe6e43febf8428d38f1b6f963c2d443616eec8a9c760fc5d3ac6ea27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd70b86faeb942954c0742a150fb00a2b95db50f480ba66b2dba78de9f90a8ed6127ce39d7163f3b4da263db655b7f56bd64e802755bb0f6d9d4879822fcfe2f94dca6e71a1e2d14ec18555471c7137cdd65c31b36136edb53c5ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15636b1ad62127e5b53171ed6a3a6ffb8d6595a47a97473e7418303b72169768a6a459caa1eba148f153e3d50e3ee0693699bcc7c5b3ad4c40009d7a7b53bbed73f6c983b9da556de4fbe7c29c123c088b46b66d8ce5d6e349fc5d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h151fcbad4f0e66f204efa694dc0e18bb664b7c48a6ce4d7b1f49d6da267aa6c67b84a22621c6f5c2874b8bf97c19c03e2e773e54f070d7ec8309d9671f6393c028cd3a481810aef8425b812b5433b17ba3f3f3119363afc9ac27fbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h75482b127e1231be5cff5d2d0f170ff1d2f84c8d7f8c3298f5b94a2a5c9a50a8b0288a15e3e40426558e0da5710c1450bf323250ac4bea7128a909b44f0f66785018c4d01e66dab8353e2c248ebb6b597634e33a1a6295d23b89c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfc81b7735d99fad9726dde455d5a6ad8083da7212688f961c157ebe164e289eccaa04ef8fc3f478324664867d4b88b4581923675851f067c26ef6a60f6874aa6f0046cb6f83b4da08421ba86488dfffcd71fd9e939048580bb26c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16dbacec7ce29b039640f4d95a0114e44698824a3f281f16362bd335129aa0e275c7e518cc04051e3958e22ba5af7e5cd2f97b42fa3090d398c74a8e80a9994aba693f59b15b8173831ae3510d7f03a649051fc34c896b1a84082a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11f7d989af3cf38cae312ac547ac176185fc114f2e1f5de3be48a914d0d5543fce950351111a0eab9cb2339dacc018e42829aa90a2e2b4aab7af053e217b16ea111953ae6736fd17eea6749ca7784d42730e77cb49966ce04d92698;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1edda54516611a3c8487cfd2fde7966b1d64aa1b3a7d436a7b76d72f9ffc9217105ff20b05d7e3b8678183d3cb051dce2db7262be2ebc5e6d52849ce8d4bba9837389f7d8f41f0d8ed9930bb18236d6221dcc224a2928ea5a2a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hecbcb1571090555a33efc7e4ad9594d237329ff9b9dd1fa6e0ecf7ddd84c6a5d1a3986c50add28c42a5fe9358e692e4608cf8ab4b02f02d5c8f11a69899d3dcbd4be0a52988cba67171fcbc9396c88ccab7645a0590dada0e8099c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7fe99c6d973dd59764f3ec32dfc95dd8c643bf50d986f232d2df1ed05cd0ba1ebe50d80022006c3c98146c74cdb84538378a4b23383409463a442b1ddef3535c56c15d310d64c513bdeab8ff5416070b700657137d4e4673f5dc35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182578918a0352cba7b311e84d8bed54060f9dc7b2544cf76116d71a50bd5844ff33e681c2294c5f85177ebef5bee9d6f1e0caad3cbecfa3af2f0d76e50bc53dd866ea83f0276b2544e00b252222313fa249d59f691986f701fd468;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b7fab9b1c464b46caa341746592c35a4356c0fc125a461d23a524f0d782747eeb1190bbbf1576136ccafabd9cded7275428517b64d4e4bacf8fe0bb5ea265435cc0d9e22105a2d33b9326fcc8d57043556eaa1ae061d41e03cbad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6026bb84abb8c8f02420b58858377bcab40afd893eecf75e4952a07bd72e58306d941981c43556dbf0938fb0a9efc87e88437c82e7c7b4abe2b6cb0a8dc8c284c70215847df3428cf16c867b0af6c4ba0979c21abd4236581fa03d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h613c678046de52f2a7475fd965a62f125688cb7a2c1676f7d117398ed8df0249434042eef3d81298ae0a1dcd9368e0321e60d81b96c9981d9bcbe5d2256c4c3d820302d22cd7e034044d63816a48c724d29eca49bfd51edd48c97c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a39f5d37f264ba71473812ef23747a86980e99ccd9f3504434228048ddccca6968bfea56aa811745f421b76aac87e301ae68e3198b042f01f0aeb93887b1cd5cbd443e5101b44490b3de02a31fdba007b8b7f7f3e5aaacead212c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af6231e7e7cd676573b39e589993b3b785c5650cebb8d1ab98dbbc73b3f86e21508b00b3571e78e406e40678e506216ec621c1b2627a10440f49349fd067858764a88dff4346fbb2101bf69bdab06b0422a1651b55da7436b78a8c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11b54becc6c59991b8c0c3acf08061cd68bad6a19a5e55543ca4c86e11a0ab37444b2683256c35f511eeb68a9f4c1d0e2c7a6915df8953d3ab72d2619da68eb1fe0aaa413de6d7a50dfba8cd5f7c2f1a08742c0b1786660b2b31462;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13912a57bdc8994fb3732a400aab1f82a794fe54f0d687145007aaf0995a6902411e8ad730753e99b5f0a50aecba22fab117272d826c3816294156fbce538d2f7d28dce02bb545a1a5399c678b47f183ab7b4b46b25f4c666755370;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13a78d2c29c472261da4b7fb53f5f711608ab262b4d5aaa73e9f595e374e2fd2f33a46aaa3ab2cd94cfe22856ab94e2033e86d489161a8974de25be581570900d61a2bb46cf0d2e53219b6c70213ef5937c14a25fc7d5a4c0b47fff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197b8846463d82e550f0bb9577f6187b564a712a36c80b9a1e977763a75a857c873d17abd24c4b280786ac82664c19343c611f475efca83a07502f4ac298172c030a70568780ee44055068f46dc184a0cbc389e0337417aecd1ea84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h107a3e5effd61f50245db8dd08eef1c9b439d8fc579bf6b2a359d47f161f5ac3c95d1d4b428acab786394b905b5cd2fb51752b913ae816957f459fbc6bf0cedba172556e323d482b949e4ab63749907a0dc5040d1e123c93406943e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4783eb7c579fa37a24682ca62d13e872806042d6e1d6e4379b6916fc7b73bf0119ad4217400311a65d99eadda47905a36991fbbd232fbb9c4c21df6a6827c3179d1a7e5117b326efc25361b32f105d0e6e4c89b08b3ab304e61eb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ff5396f03f757d49badbc250d697397129f9b5ea12935d21a83eba7bc5a8a7c50df153d6b91f0484e17689fd6e01cbf7789e12e5488f01658ca4b8da7f32d9737bbe24cd34fba243442514298e7acb3ccb9ce84336f2b147c71df2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h99627eaab9d02455fc3bccaaebf5d2ee354d5def72c68a7d3aee425c90a0b2e7dce1e2847d92023286052251536118eb9ec136ef065a81c8af1d0ed5db26ae50a7ee0e5395994ce25a89cfd1e13497e33df436d01b27bc6da53f1c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3a900aea116c02877520c615889254af4352d0fa5662503a3fc476fca76be19cc841eb25b06736731d8b3a61af8640d893ddf04ac8e38de8792ca1bc5f182617494997a52f484f90380e418fbe8720573a6137dd7a3d57d6b973e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e78bdbfe124e11ad24d317f73638043b20d59313f156c0cf0c514d10ac3ea86619f15fd5e91f6cd234cc33cf18432703beaf48da59fbf4153ae327cfa24500a828d16420d84f91e56e739f32e18bc120a8de181c26de0c3a5c8747;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h852d90cfbe56885b2dd42406f9a3d95c12765e49988d25d8da2188aaf8f2b298f58671e0b6e3df0442d30b154f4964ccb0051de50f6e9282c0e1293904add35f278c5f4f1dff0be3abfe08b77d8000c3c00b2718d92d749e4c6246;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17baf39dad2f1c928d5c4bb19786b1e1dc9023fd559caec96f005323e9d52e66c336694a10e84e6e28558052104f6f7ee1591874077c76087c6aacf6363c3474fb91fa7ea16dc0fa25813ccad4bfec27749150ef7dcb9124aa09a4f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ba969e128cb537efcd08e7104e1a982a4ac2f760a02b42fbbc62db76712442f3b060159d4c7eddb1eb2b5c1741d1ad30bd0d7f00e8da2c23540822122437dfb54bd0878cdbec8704fa36bc420e68ceb2ecb1c532407bffb183e57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b394b8133adcfc178a3560a51f564f48cb634cac4ffe74687838cb5048093eeb06b3d91ceac14d653420b255559d438c25f6e1c31f36fcfd8effe5d2005a0eb0e404b154c3e66734bb900ce6115d4daa3ec715fd13549817d3255;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h118a3fc9597dd942a249af4a86f358a5e84b266d634d3994665e5dee57947d6528eda26ab303015bc554501ddfca40c4e4da74fa98280de0744cd578c876e8ee41790e1d81840d9c81fe9896de82a3e010d6ab8e5c87465e0884322;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hccdc36ff39504d61634464838a6ebae2fc8cafb614878257207a6fe5c9c44bed2875638b67d1ca75a9e230adcb547eabca8f3eac6ad5932c83503659c6c2381c4b71543d4d176524dcdaee47059acd4b74fd9b86315671afd5cd14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fd71bf34fb993189745dab40847764858e289434bf88e1981a6db17a7700a82c0c131b60255286aede1508fe12b36ba91ca56a0cdfea4f89899697d53a623a804351619931047873adc8c58fefaedc05e662d3b8478c669ae7132e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c08b572216e53a8cd176adc93ce3c9044a97cf1104d88fc2ac094b3090a173298f2167625acf39185dba61161e3c0a44912c7e855f502b4486863251b1935caf38784c98a2dec3e631a091d4548e20a1e47ff9a64839e8c16ea4a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7d677ed82acbcbafc2c08d4722dae3dcc03de071c42b2fd8dac3fcb581d51efbc3e1fe3484961aa07ceafd1f34165c99ff7336103a2c8029c5cd93d172924ed4334ac925f05f512b6d4e87682f7dd8ff865713fad88073d8656fc3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d2957435c646c2e77c9f514af2f7c4ec878f7bf838db3feb78fbc2546f62bc7dfff42482b077739f337ed644d32911ffa86827d04a4382cf47ff8e7046a2c3a7a5ac5163fb3dd0053675848de68f6cce63c1eccadb3bb49352c67;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h56f7cdb8c231504beee0456d2fa2124e3fcb49e5e4cc5ff8ce73d346df141de83618e57c0826807b40642a5f1f906efd4e2a8bd68fc24809c0ea229d3f5c5b8a541de75f6039c4e6515bff33d43b994d0740fa93619ec5cc72815c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13dd279dc9399da0cb668e9e23b5f33dd760f05b21f7b9b08164787be2b3863584a2d7b28e9776e338500675a92ee7fa38a8b5709c2728508bbf6540a4e94d2bab03038461d2d4633d44c9b0de32c1fa250ae96cbf353f2ee688aac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h87704b267a296f469a8bf618c44919d8e58e430718311d214b9d72fb9fc1f4f1342f3dab3786af75b183b3200d0544efeb22a38965eb3e8022eecc80125eab8290ed3b9c9fd0757b1b6f8e86f3a0c0ed35aadc6df8323be899a81c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd6045230beef238c8c3fe372c938d9e23eb8ecc8606bc19951782ea53ba1fb138570b86178694b07ed4a9715555a5c280a384651273a936f2aa49dea3e46db3584d7509ec4b511c76c528dc4bc6ace57ce788f953dd2e84aed8c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13b69e50af5373a5a811142831feab945cc06a05c6b0ffcc34e18ea122663005de8eb9050c1160baef1d6c50458df33c9e76b8a1ce57672c97dd83adb47ae59708d24e6d67a9ed03546739738a50e49ff9f8dbdd0b9eac80c1a6739;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d9335ad4b80876a0afd92c02de277e9e85e1aff31c4dc9b12c2b483e3cd1b7d7fa63764faafbb29cf4b4dce79d8e8886b0387851700bd3417ac07e7fa9ad1e8f81967e416f73f281037f7ef97c7d09063a7d4ca47d608bcbb64e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbffe7e1a172f9336a8fc8695f349fcc621da9a1693d5f98d87df02afc45fee9725a51836c9adeb5aac06d6fd2254e7c6410f786a96be242095a890809a17d0c8a17708bc407d3f797d1c046bac41762f5e544cdbf051dc4d37c179;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h547143a305541de0c1d306b2be75ad2db63e8c6330bf9348b196209847620c129f42ad73f959b53500fce64c1f07280f13475bc83fa267850badb7aafb88e62f6109071df9813e1b876794ca2e9b244e8693dab77ad2afacc699cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h129f30ec1b568dd447e77f39293e74b1943c1df0b1286798e533428b836e2f577fd09022cb629648cc462d73b434c20cbe7ebba4aeb32347ec54428faf4a99bd1102594a6a03fcfa56512d11070f66276634acf4b2f4e8920ec0f2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h26e44cf375045e98dfc9496429716019774b3758959c7cd5baa47cb27c7dd0feb37455e7ebd69b98278564bb9f2aa61f169d96963d875d05363757486100a7b7f7aff5ceccc5895f6ae23c577d92c2f3814bb3b7c29c919619bb9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd16ed8c320077dff90e636836d198cd7b7eb84d9fc120552878013a4212dc4ed2005285bc55c3d3555fae0b88b2c48fe179a1d650aa71b041dbb7f455b20179b913210a1747a3634864e4f856bac12ea4da727949ad91d6e7d509;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14dff5b0306e891832d34a106ace331c934d5cbcc406d0538be1d54c6232ac1019cea8909fb3c0d8ce092ec5024f19a7c0082782f574a44847a8008b7ef4ba613078f54ccbf032271d4b1702ff6ff5487f3fa82d253688a93353567;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd5bf3b17e56bb0b5a8e9dec3e7c4abc27b3d1f976d45100fe571997b5a78af5ef4766f122d83ec2d73822ff45f774e374e5b437db6804ace936038b1a135ac0865159a10f1125a5c928a47c450e3f451c3585c0dd0f02ee675ac3b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7cedca97c45311adfb5cb9dd58c1d477f20399a29cc350daeaad596f017a6ec9db215d058ed1e9c3e8a17bac84a639c97d7eeda490a4bd4c2b12aadff026fc40f084bc90882f8758f25ef06b629d2cfd58cd65f6096e706e7d0724;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h68147f6c12461841c6a30f2966678339e3ab7f7bda14f7dc763dfefee2d8e5e03916292a5b4fdb82eaf00613808430c4016471f09886310cb8f7f5fe288f1d964c7697f9ba164061ff5975584bbc224a662eb15e5b2b5dc2cb3ccb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha6dfe3038d4fd391557c8f3289875d62b44936252e13fa93fe41c5030ab267d708e3d78a0851b488fcda27652568a6fc23d1395906e6fb11ed8ef1bde16fa71bb4a9723fc5d32744c139b9a27129e163b01b1f271fee6d0a94a728;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17478293bc2087521387247caf645c51e41cb16b10fbf0c9326471d6d1d6cd1736138bcb1e8d72e2c5a9cefaa94dfb1edc876bd86ffef93065eaa1a7cc0173e8f29bf62cf8e87d5d147430870fbc2be642de7fbe163bd14f10e2c78;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c21427d46fbc5bbcbf60d14be172797d3f6810d45ca1c4ebb9193ec882f1a2c86507357b7ef5915e31156a4eb2eeb73640fae3df029275b3ac85bfdf78d52b25c13ab68c2a0ab340b316088c1a84b8fb2b9cde4c36af31e2a38a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha953fff2bc4d47a028b3c00a261919c50120fc7bbffbd1447dadda7e4e2cd41da2488198500608049be4814d1a2a0f967bd9f7570255e2effa9442550c17c70e2698d728cb9ede62d10e6c241ecc2852b6133a5c81b53a77587cf2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b1e4b2f7477541b87c31996ece886d55bcaaf0d9f517b9017072488f2612b5d26014ffe5e3135cc7b1d59e4b90bccbc337c5a86604f5ebc9127c7872c0b9f72aa5e180413212937d3306de67e9c0798564dc73f8d73cd3f72f53f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb3975d5c5bb6551cad0b03d67f3f87496e2f24a5cd3e3ac30dd5a2063638e7e7f56e09a9478edc9050bc398f14f7a41f3bb48ea2d4ef56b962e3c1e73849d0db9fc22b80933ebaac6278be06a90c9a1a9552de7fe2b6284786eb73;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36563d4624fb58cbf0b76f58f961beb84fe6101c13522cf37e441604ea49a269b4b953f8567d6d5561ccf3452345e52b30794edba4a5b85ee9a1b1d8ba0f649328b6353bb03b246a6bcfcdb7a8be0e90f8c8c50e4c84fba91fea81;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2a78050d6f6d0739e6b4af32761de67a3385619e698b2bb9f0978eb3bb6d85e40ed335728bbf1f276f9cbb48f26e1be71ca190c8cd51bd85c84b321f60527ed4723ae6a4ce602f1a71dd062b3bf7138c9cef13a7e4ce14bc26df27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h549279fe30f30ed44103b6f7ace7e08b285bd77678e9a84a240fea78bd03d0bcdce86eb7526db64b20ca4a0e583e130f21fde782f4476610c04f01fb0283e362272351a39c0acaa08e59eda7eb652c00953deaee73758972dc96a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e49238425bfb625dcd5f120d12514c5f56f78e74ad3d5ec7b204e37615252e080cc83fd223ca249893189a99e5b3da3bb41c355ede571400b75c988856886001e0e6d9778c07986b3cccaaccfbc47e6ae4c947ca1a1e73eeb2fa21;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc12ea6d1946368c536b80e2ce488957b2126b52a878cbcf384f7ea803ec885103a5370e72bba9e59a5c6c231838cf9f0e35865f5f24bfc3b80d86cb76aca45412d4bbbacc21cb8f88c7a4b01da4a266453fb75364d5d2d83e49d2c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18f7c05cec314445c884feb9f0561ed22bc6417576bc91b94ea7b753794d6de75a9404aeecde0ba1ca4ce47c3b7f7529fd0b89621b22683b5cac7944e3565cfe7edcfb200198277d8a4f9093362b904bacdf03d8b01592d83987308;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97222fac101f173e6e8f82cb273ca491b90c577a4cbb63f9ee5f738c5b7ee4ac1a9b83b25dc4f6c6d23cfa662de50fe865fefe2b6a1d305e7d9cdf91ce5737303e5c1a367e10b5e46e509036095e109231b1c8e4f5b4d9e2594e8c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf02426aa25c37a26b8b4a11446f450216999334880070a0b6ef0d7f8afdb6e8b685222628e86e465a8d997ba57c743baba918d7f56822dfdf0f24095758e02adf7868a8b8463036f78681876fb9dec66cab910d7c3b88937ce8771;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142a08d785b5bb41971cb75a49c66730c4748d15046a1948c9f3dd8f0e2aad3d2c0392f44fc12395cace875d284cf5c126c3a7587e19928987ee67fabe5542ea0988a0e7543e6b86558031c2c16462b34f1225bec5d18677b2dcad6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h115fece822751fc3bb9c25dc5daf68b69b8eb2a4ef2a9b165a989748052644a756d43d2835f5b4cdca8dc4b027bdabbd309fb239696b91adfb975062ad33376bb79ad3e783c6e9dffdd5af4ce959ec3c3f2a50a9f78b78430afa686;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f5ab1e7969dec8377f17c8ee2f07026c2cca27a58762ecd95d59e9e21dd8834e765c0ef6c239f908e627cbb9a5ca7135ace33792abbb9d4c3c9113c25ef6a20dbde44e86787d10b31272fd2ad98ce9e11ab2822127f38bd5d5262c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha952ddaebb1422173a9dc6ef21d45ffcb19a9cd912bd5fde0167962a720a0fbf7248d911915ae6c0cc1ae6aad674265af9ea5928f102f533a316388647b2ed2345d0d7cd1da20e23deb8cb47b9071470b2f09283a64163ff4e5290;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h72dc54d9f87cc6500ff0898803fc75668044c259b801045a66be4a9a171203f9fc09ccb81aa97fe2fb21fe15b08c9cb504f19ea78f1fcf2aea9dffa95d2a2d6db1b931b40be73e34d6e6980db262bdd7f9100adebc375244d7c2d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c0bcd85a8dc9f86dc07405ce9820b9356fa724d0ee8150f0b2e1c242183701a1ac75555d54d4da20614ee3f3995b986c16c051c1d9a13a8eac3b25bc4788c7720e9ff9197079f163123696ac00d1ebe5b808fac302a9bb8215b3e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h153c1d72948a508b4961f95db369f550308a9429dd658d521584c1be8d29cef56dc0c69b567173c21e1cecd199c4fbff857e45baed6b06c7aca956d5c35c3277e1cd7669a8a2231fbb7d702527ef0c300a3424173709ec617b1c961;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e500298d58d19424047ed28b682b86ca4d055cd1f6f2826579b4a4f4948a266807e4ffe471efe2cbfd1232283b4b072c2184f146e9da99852710553214a6b1c468978cf0ef1e5172bb18ba816a21ae7cf552875af51299fefe8734;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b8d2b6912360b80d514b830b4761f7029aae988d13e551c6d2c7ec7c20d244355179973522ce839e638aac7efcc0c65338194d89d2584fd0032b492e427fa1c92043dfcb1fb920be0dea3c79481c7d5ffdd719fd7dc389eb93600;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc8c5c888bee6afb86b3dee2988cfb71c24968b0bc5db25c68f6363d92b45ac4ba42b2dcd2c34051503edf63b7a94032de223a92ecf9c55caa9c260a861e70278d191c68bf146c5c978b55daf702da95fdda738b1f144897deb4f41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e36e40e23db62f67f33b16dc0b4d4fbbc5c60f3053a434e5fb19ae3745bff6b63474366f1c5ad623e957151e844fe0499ddb0dd9efe21db88623a0a60d806ae33ca86b2fcb4e5c4937d30d878f11b9883d6e56dc6e51b6f7cce1df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af647c3769bc77fd920d783543e014051e4acfe1416584b13ac116ba6fd30a13476d26828ba179f2f10a8a7f6ec2b4767ae8d64ad19b32b6b422608698109c41f400749ed135f111e29ff97be5f97aa628d48cd36b30bbfe77f4c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h349728a48154f1ed12407f74c6a2cdf73747a1ff2b9c6a41760a4967f94414ee674f1679cf0cf14edc74d43fe6a8fbf2a18916a228f2475baf91bad462fee19784b965116fc977f73697d0e020cb6b45deead60c4558ef72c41929;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h46596dbb438e9d8e6e80d900206003281baa789c838298b154fce31b25d1a95e700cad3bb13c34b4e2a67a87d0d06e226490873e0967fbc57f56cbdd394c6407d31507a5262d080e48a6c6733bb968f50cb78a7a79de73f2e27445;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ddf8d074fda76dbc342fda0ac24c8b01b00afb71ca29f2d1bac4f46493a99d8274081a9e4dbc9c3d268768e891508f2473a6d9f20047dea899bbfd50a28873271be61a39359d92ff0c704b9ce285621a6568ce10fd2dbca23f38a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbb63733254ffb8f13d9d15f840681ffec1603d156d24235ff81adef7f174d06c37a0cc3002f5d8423b90dc42a509e2bebed2cf8caf76c0de07fdb33c1c0dc64534920d5c2127f409a1d08da9a0e34b13459633ddc4ab30a1a9c21e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h58ce8f0755c7f6725a3d2e2d6ddc1c59078ec4c244ab376f0cf7e30c6a63f17f8448592638a2c83a3a4ba43222015cb30d5287912c28d3505bf985436f5cb1e469cdda8adcc08e148eea3893221b78a09baebbd0a84938c47ee43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a15c510383a808aafabe27b8e39d0538c57cc5298d4aa778fc8aac59c20942b2daf1bddf206b7c94cea8d5027db64737711f1abed4c3cef28ca7bc47031f6cd49357583387735a921b4da89733b1cd08878d33ce478c4cf42c9db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe17bd2f3222cd20a84ea030a49d87e78c12fe08d9a1b8f94156ca907db0bcc21fd6e01fd02b211f5297b5271c4d95ed820c97fb3b807cc22e75091b1af507aa2521c2b611940feec9420488c180ac5c78f3754b4af69e835f7c4d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hed9bb0abb0f3ced050fd6ec34802c9212ac192ce4e8f377d0d7fa448493334c48a26b26914eec9f17fdaa1e3f02f3abbe44e0ec0b799587e781066edc472cb6ce5da1ca1e4af1d79f3c5c549c7136a6b1cb9fc7e2df1faecd43c99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7177836096279dc05e19ed3d9ed6b7238aa9cd7fe287f3cb9dbaa3d290532f2c21a9e56b687029c74370f0563c4ee1d63b330c4f1be5aeb2f13a24c8b08c667e3cd77ee6f590d1de3c63482e270a1c05d6910a0e5fb63d9742db0a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9363bd990ed555a7ba23af5565cd830d3c15e0201efea4a531ff245706d279eae46303659de7da0a10286c3e976393546c9a65cd0787c5fc5d8d7f4b3fcf8470c44d3f07eb82b9fa7eb6df643001db5ff4c7ffa9070cd5c21241bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b6682240d772fb2610383bd87958fe5615badee0516a5495ed2679cee2a1a2fd0cf48237ba2b54ae5b4b9136dab4dc9d8a51b4d660f08086b99ead4fac517bf50e566649668322f22f33c3f58aa4f0f7d8c45b2c874cf54b608e57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h993eef459ee4abe8efa61be5c102396ae77a0d1efcbff51fe15844da40082be1bfc941ff9b7c0c06719932402ebb5f489fe65b31ef83b7a48b82202e02662490cb371e6e2981fedb03b7d2e7602d5a5a24bcf00647214ec24e0776;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha15e4c0168d49368b718fc6f758cadb80162b8b48f643cdd3545048beb11244db942c013eea75d98c328b0ebed0c2ffa7abbf33d6c1530c5802ec3915d4f658eaf6659160f22999f729412f3d8dbdf7474b009da41135eb7efc44;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8f6093bdfdb9b8eabccdb07fb494182f2968e6d1706475aae1856190d4a3a01ef897d669aadeeaacdc6249b43533e1069e1b2fbf6fcff25f17370e09df7a16bf1d50287f0d54b84ef010bcefd7cba667c7bbecf64e423247215ade;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3960480a8948989458f4406e31267dcdc8e0ee9beb8a0f76826037031653be3a9aae75f1c61c70c3b356b4ceafc0d334c43c107d048f377668b2b820abb6b77c77ef51114bb9a8c02c8ed073a8562b37b123f6e08b094c9ae91f4b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14757b61afa53029bcf2b1f841cf41bb2f1d9ad6d4cca25e15653a6a9cbf01ec87cf39d36d258fa49c9b440efd9e9476bc82215bd77df2ba46a55ac8655896ebc0e1918f26d1d187ee7e66684ce783abeacd470e653f047b858f6e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19250a4ff0229987c845adad08b51543f332312496ca945c71844309335f4d98198833eae75f335e548a27e52ccaff2beca556e3921adfd1bb7f4fa0f9203ef6f8495f721ecac84edfec9086e7f43aad7a1aecb1c944de06b95b9d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h129a5e153c133534b08ecd6a695726b37ba0fcc81fd64ea6a9338f6041d840b95e8c9bbc3beceb438799ac966d24390b8b21d1a5aa8ed110f61ec0024cd311b0d71fbb9655ea077abcdcf07428125f315ed3913ee9721284f23ac6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbab1543a9619d04593db89259f4e6b6fe4acd329919ebbaae04fe1477f542152301c40eac87e651f4582afe935bd944aa4d4162cfafe39b187fef292d6988eecf3d1ab34e5b46b4162cede481a4035d39743577f519b6f44e55c0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h707b7763c47e205ba1a903d0c016aa2b496bf0091d4fd0c6e0537653a0e3e98cda30cd04226ceff0ce444be05cd87575445a3e42dc0dd482d7161d17efa711541cf8aee1227ecb5d2785624a38d711914f2b0c3e5cd716cbf52fd9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e96bc6906d16b2f1aeb36b7ca50fc3ab54c9d2751dbbefd6c6c6474d76768d9cdd1f76e0ea05c7b8c2f8ed9023ffc8f3a616e15145aa1537688e79dc8b9c5c928d272c88f4939fcdeb43a7fadea914e15c8b30bdaa9883390026d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h678524bf53a09d7875709ec8570624ae40d310191e4d29def8727ec95c7923714ff065a0b946dc2ac9e69b21857405087fc5814ec5818e7d67c182d3284c6d1641bc74459df4b6137eee3d3172fb426ae0d19e7c57d56e65a5db18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5ee5091185a0e460f1870ef6f353ebd0f5cc31bcef756eac71620fe544bf375e4044c0f7967ff33a0bc5fcf5d101acc435e05f5a0c3b412a212de47ac42334856a10298e572eb9336bcf934fd936240c64d8a10e4a8ca3c7dd84a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19fcf9a1bb969dced29cf76bd33916ededac22142ee9eaf3fd912048459eddeaf42cb85308a1cc91cc23993cd6b0acd57216a8c542b7a38cad34fb3050da65d9f240d53270dca2c337edc853e14831e7254b3b659a0460b01f3cd28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd4daffb9b8d707533ffdb52be0c86208153a410a259e69db5ab978f97f6f51e23cbcdf0e044429c3e1dc639d8d69a94db3d3643af6975cca443c4e6825dedb132be4448729b6aa8850062eb153c090a28167cf4b072676282b010;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cabf8bb53cea907152dcb27872db6de2a600b71e8a3dc7cf41dbcafffb5a99f463c20644672cf4258e69019a40ef1fb89f8185e7f196f4b9ae9b99f63fce4e76811664469e417fcbdd1188f881bd1b6cd5e13b7c36eb7e70589ab0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de288faf1e087e46c088e09973e17a7186ad61c432e81fff675216787508888c4fd9f19694d6888ea68bc300994603f3a2ff1f798de4a8830776721b5c976c4c6f2551bb3b96090604af80495a48762e445eeb72101787791ac4b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h986e48ea81aefed0ab7e25093a6fa3dd75fe81097b2f36cca50d4fa3787c08d0a76ac0ae40eb26bf0e4c33ec15684a6f99bdee0f996f9d14824006fdfdc5390dc41f15e81f00c4e41d037f563a12e18f55a282f0afd24f3d308aaa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b20cbfab3a65db314f233d805c1529e3f7696eb672cdf806795c3fd8f1e96811a71af1edaed245c86299d5a053eb3b622900d693e3a09fa6cd4f914edf29da48d426770a58cb59572c3c724689ac9b8711c7d291e955af082c42f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10fc1d3a0e2b5a86b7e2f1dd136a6798722019a557dd92cf772b9ef8158828e25c35d8f7c7b51bddb4212e5efc9761cdddf9cf00ae46ea5d203de35179fa9e97f9e2b66d4508bc5653dfebd632abc046f15d7559bc7f80c9bd8b9dc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8626ae386b2944db0cc2fd365e7a3db05d8d60a4cbb62832f3af0e52c5e16445e4feb0af3e70cc8710be10f18dd11e147f1dab86e4da4bbd06c109758672c3116db6f8a7df46160efc02a4660ca0ce8279862b98adc58d7e29802;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17662fd14f909dc8c3560b77a07ff349d6a420f5f9251cbac50d95466084a60cd6aa03f31f9f61dd9724e5676d3fc154b8b0c46a2ac27552d3fbde19db66cb334686c5b8951a47727e49a52c8141f9b0399a63393a301b5e1dbcf26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h144bdd64e9b00745e295b243b75f4e7ca6edb273303ed2f975a5d5392340c6d0a806c9e89759b46666ed68e7be0fb477bd7a8e0880a8f36874711c742857c4e1271ad0ecd65e6eab570a6fe6036865e6e89fb3556301aa7c16909b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8b465d09427906e2dd9e4ee495f96c2061e3235eeaec1b72c60dd23eea3d4240a14c27da3d2995b132109e9bdd0a46c5761019b498caa8a3cf631dc163ec1996235c10816d67be41c182f79bfd9cc33ad957687205dfb1d45824d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h104a01fbbd423066a4ec93ca7df1cf413db84b382dba2bb7ae83f8b5e0ef12632fc44fb48c5e9e0151e279ebaf002ee1791fa2b9805240943de6bba32530a72c9410f115da39555dbf720fa5c91b10308d8630a07128c836433a6f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h110ad460a4cb2cd5250bc0a5d22c8d1707d34b4c23dffaae98f597325ce825d09b7ccb806cb7f642052853b51a4775334ee25d4c1e12e8fe3c14cb426968f4d38c32ac1e171d330abbb217f9dd3b236f2398d2fdbf97c4b93c96812;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hce30033ff94096e148d1154e077b0b9ab9220b0fecff10469881d7a57d90efd98b2322d855953edb7a32f6c9917657e8a6a6132fa16b17bb5631ea542e5a688a521cb5819fbe5d2f8ee068a036a446939fb5d375a0b4cf020cb5fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11cb27bb1cd1238508dfa9083f83720dcb96ad1ed2c7a385794c050edf8cb5d49e63f66d2d7db0b513d2c6f5ed9002f98964729d87626fc3734c6b77610dba8d13308c119bc562fe9ac9b828993ed6bf5e3990b5f9d675c4507537d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e86458048a5b5aca8b4eef199aea0ab7207b57760510fb127ee2ce59dbe07a370e0509c08da241f89640802e6ffe1a9d850c7474c0add7965c0856b8ed6539cf1f6b435c96b9ac13925c50e164a93880a70d70a627cd3e3f6080e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h63d54411ea6fb68be3451f09fa896792af03051882db16ad228c03e60bb54bc736f0f27189a14adfebbf0c0aed1a99eecd5255cada6c1abb960ae68e9270f6ef6a02004cc01222227ef71b2b7ba8b7e83e2e107a73f171f7055962;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hae5c492ceb7a1bf587c767b974085b67d31abdcba5f02aa078d0161fea3701042397f86da6248ac9ae3c025cdbf4faf2269bf50d9b41b802287213f7e72fa51f03ef390fd9b3654d0120e7d87165c4df23a23ea0b8874ab7cdcc06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h109d68c881c735ccbc7710ba8d08db27a77547dd97dca626d27aea9e0bda218555c38175d726690b39eb549d3c91209ac435581d3f36fdf4369896e4b89f42efbce0acd279c3c8c2feb8dcff2747e261ad49c36447443e20aecdb9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec65455ebd95018859a6243b0b2fbe7a8f6d1b1e4987872f4f28c12a7ddb1dce16ef9854c97708d503e3998f398295683c3008d41d563258c4d61f8e9be88576a380606f4177734da38f6aa096069cb725a5d6a827525d06938ad8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ce50040dfa75a3f6332d27ae740a0f7f36e0a9a48d06d2cb4a6a6ce783d8786a016cb2b77d45bb232fba629e82d3196aba4d2f2e4a4f69457f11a4987919242bc666ef3f305b1ae4d96749eaf2ac5d6732559e602d502aa1bcc3b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3246fa6f3d571e1b24065d8458707661eade03b21c1cdf363aef8bdf142b9aaebc4169bebffb92cb1b31fe5651246da53a429328eb31f7353933ae21fe004e742e5824162abdecacf940f1a01814e25b713f519fa2eabbf12876de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ecd8d498c058035ad11500cba168f5b22389f9a4230c601a56c832673d2013a5e8af08b4659c1f4e0e5fd19945494dc1c197564c34db3922bd66f60ec71335a1220d656a18e5210178e7465cc9d5a6749aab0d1e8264b65ed711ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c8e24ce56323cfab246c249bd8d3872a78497011f2a61ae2f38aa29859c2a8fcfad326390795430dee98bd5b905fefe8ac51ce59261fde709522e91b367b71fa9fc2a4f3eb37626a2b8fc432d0ba09ab9f71dcb54f0eadf5229c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4161f5dea6b4ed1185394f315b3876c82c7f32447a45346de4f93cb9df7f014b3bf34f4e83d8724871c84582d69862f94ed2beddf143eb46069ab89b3083e12e007677444df60e3943708bce97bbf262e174f5f48ce3805ba8ccb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h398a7f4accce5738c16eff6fbd32f24b5a31490c66e2ba3b46f50d68ddd0da18e35970255c71d5a3576e83dcbb468c842af42687dea85fa91d690593821833129f87de0525b78266f957070daf56f9f0e4a32f36af36907e6ff463;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18a7bc6e0c281b5375bc65edbad80d0aeed397435ed0358bac2c917b128468ff44b506f204e16dd116a29da15d781d97137efbd9e78de39e5e049171da99770cc0979369de75252eb0e8c966a896d32e79a575341eaac37ee7eeca8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b0560ff0032179e66319f0fbd40a76e3e253b367b849aba5e3de1ecfd1ba9b2a1f7b86c0edc8fbefce562af1b093d3e6c401f8232a61e41af47d0bb4fc7ec228353974c11388e34ff3f534d394c55764340d75715f0531e4635110;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2a4fb5ad8829b26abfd112c5dacc5e5d3d7d4eb9777c8519bacf3675baab74f412e56bec1abd51bef1ea7b24b5b1b5ec93116f5e9123b074827d0794316af3ff1dc615f339853a4800c865d23f29b5fcecdf9404d8cdf66be2a2c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a50b7128104794d0434ac0b7cdf5556db7c4987c27e528cec9d446682c2d9c6748d120b3b7f619aba67e64feed9b717931f1f9760aeb56028ebc3710d202c5d390e9aaec9c8d5d909c4eb63e3edec0197ef73e6d2875803c7c04bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16b582adb4b493ef5f2123e05794e0c09ae35361771c55cfff12aa3eca9df9e30baa4521f9ed7beb87c390b207324e0571c0957a67c16b3cd9ec5f18e29e3b7cc59beb21a45ecce30da0229a23dd74c6e3ce42491e654288edbe038;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb6d576ce0cb1f159d85bbf5314ca719697579f22a884ac4882f90fd14006c37f22223e308a66c7e72c3bb5b3e864cccd2380f98a4c60b09ed5c5cad7f5ad754ceff645456f6145473c7561184e461ea5cbe31770d7d81a122f8e99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e3a1d96108511d199e039d0f7107745e8b5fa6be39699acb476283c086142b966506f443f61710aaac766d4180ae0dd27f83fa6cbab261215004ab29cb08c313c610f10502a10b70086d74618e1f7d59493696171e15aca3a0f41e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8815c23deaa8109144e2578e716fdd4ddc00448ac3e74824481eacb95a56c0b4d05a44e14298078629c28b180ad5a941ebc7a2618aea16443076987f5c86a5249d39e980947ef0d34cf90780d8205764598513c08d2f285bc87040;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb835694b365a05614fe07a9bceb45dee6659546185e0646f02991787fb358f8273a2d78b2383a5ab2b23e1d6c1deff24e39cbf3bf9cece12ae8db7da8e96a0562499fc4491a047886350a97d2aa7dd5c9f3761fd3e778529e81e17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h190987bc6bb0fb484f6d9c228a0e8448acfaf60da205404d3e9c23fae1804bdbc29860dab792b992e9467c98ddb86f1fabe5f51f80f143a8d18adb451fdbe8993a3f32f93d231daace880a699a83947575e54547bfe9b7dae40cdaf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1890f47ffbc34e5219b41bac49f587dec0d5a7e56e5e42519c610c31b44ffe24efd7c8ef80749819667a248dba0064f4ecdd67fb6270937403082c6d5f304f5bdcb964f0fe8a5a05b2f2704e7ddd1751777c5895ff4f029c3566fcc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf68dc3c7159e9a8083e5e86bf54920278e08342fb00cf61562018fa401a63c25e7a9737239288b7a12eddeee051c2b5694331ef641a2c110fe6cf991ad8fc022d304a3c55054715411b6e2a9629a7ad385756176e65320c1b1c9dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d65899a91ef79208d4de5672a4af011af8848cfda6fae161b08d96493008a201bd734554fd8f346f051d9110be304a6006ce3a9583aa4f722bea58e1f1355c51e84d9169af36418f105a83f6f4a4a0101e39eeb1dc019b9893ef0d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98d7232c091803c41ecf1784824a74d8c7d66742440a71b8deff56aadcef8a1106a1822bca9a22b52b4c24266b4495a754a279b8579a8a1877795c341f0ed8b993e616aab53299b281de83f926208f43e8525fff4effcd106f923a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1780eeb4e291e46ed7aa6d01b949d9e10ce226861ee09bca9c9322cb1aa02ed60c307d548bf627667e542d2cac10ca88f7b01df6bf1ba95975e6007402366d528e628cce8c7776755a413f6e7b0c19283a0c24d8bfa171ffc15e0f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha202484f6724ccf23a482cd10922f6a6aec1f106ce29dd4ee02b94fb4ffc63640d2372c1464c6ef16f1334b26e5c679a622dc760753492c4c82d4bd95c325e7d8f4717f07366c4b7d8b6328bd30f187338662411aa2df14f84edf8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e213f9b7cc29460be11711ed9f839395bb1a67d0256bc7c14d0e872a36bbb81b92edd906f65561a62e39e6d552aa4b575f3fa93a7646a8b8261c86dffd53c46b183ecbd189e01a1b1165a814b3b1585fd642040d67c12cd4924c84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h83b2a5e216c573fd1c5a409be5fa99bd57b475bfb72b328a131c1399d83028b779cd5c92ce3988d25d39de64294c3c2af969fb7abad2e2dd8d30f8f1f54c74c7abdc66ff6e4b9c5280e780512d7053b39ba9e012763f9ba728d7c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e768fc336f43b7d6c18e7636e2dbf4bfad2f99a1a9083f5447591deaa371121d47a13b1f929706bc94165ddd5fbde07f2b74e049bdcbdfc9d26ea4b4d430abb4c10903a98fc7b1a9e42d526761b16edb89467da166352b340e84bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdc0cfee589445cbc9c2e99ebdb35dd3cadb58fb10ecca43246a74ae3273dc79ed78c4ff98b4e06a2f3f0a2a7dbb5c0b99301e1778f3bb223e43679e947ace3b2cbec17c77f0518eeb82f48113a35e7beb7e4c1e28c8fce322016e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h761ae243efead213b94b342ded1715670a838bf1b51f426b17635ac82a0942f5c8a23721448fa5a256d09cdf1b97fcdf51b48d2d3367ca4c9f9844af312c3108a6df5d105a88b38f9c72f987e9e29af9acca89b2637d3b8b401df5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43b45be28509fd8c4fe114f3386484cdc2fb0a70fc628e316c8698095a63299762967524f14f2782f7c84588384ee9d2d3c3091fc9308a4fc619966ab804575658ce9f0b1b64d77f8ff9b6b4f0792044dfcba87a5237153cfd601b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19517abb9f35720b6b7663b542467a7ed6623bb95baf847a5f1f2f372dadac4a9fe690e9fee30b4f62319259bf4c41109f99a5df0511574ef47deb8c1a272d06b169c6eb6801e693a246389d592dabe26efc903a4b448d8b12a8b81;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9463d1cc002aaa2bdc4c73efe53ca670f6882bd59742e7e6ce0d254c9a07f9668a029eeee8635bc3568479a3dfed128e012504fe8b6aba00dd8a48131fd22ef2eb95cd098743f51b60d7b3786b162a21f92fc273a5a971bd4716f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h127cdbb5221e0cc6592665685379ef3043e283c2f147c81740179bdd9f953e7a20a4c5eff9252fdb1d2f822393fcc1fad38382f3b542794a5f7df64c9c1b639668b06b1d1a650c96d543cc071ddd7019a07d48ad05150b49098da03;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h98195bb81bb45d844a126433013986be997634867580636f196dfc51e4309d460a61af735967388a69054dfb4815547a2fe045387eb9e8f065e82ef31faf5ba008d81a3f9928a5cbcd2288bac4123db42cb4b37c8e8d9b291c3bd7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h22337889d4b29ba24deb7b049ab07a58820a4c757d398c244c233b0fc7a49e26c435de2a5b102ef2ccea60fd327575b6e8143415ea515482df796b613e78536f528772a14755d6c4f40c2a37d3cf501364f335cab50abb3405fb72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4dba834878431b98c88743c581154f88e8b8524e5c6cf62eaa88112cf52b53ed34714cd4a0189caaaa7e4c01c4ed57daa03b4771d9f64bcd72a585ce73e063c09a54255f950e0b4090c161e85406014863ad052cd9fcf3adc773d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h160a5291f18d6854599dfa1e13f3f079121e422724128df15ed7838bfd164ae36532086f35f56b8f705bbb1a2065db38a8ffd1a2e0fb22aaba9d9d71391400a9c928d13e0619f5f9867af870977eccfc7656ef5464f33d4b4de8cc5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b030f7f25d17015c443d4eab235f7737a3102dfcf8153dcd195b8b483b7f681de188246dd5d61f8de31fd09efedaf7c0099831acbb9f50e3aab7ed9c169aba20b4ff0f547d3dbee3ac001400656974a59fdad7fb57958bd56d8aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2cf34f6b313e1ac7c070241a7c95878ac6a694b4525747042038a0048171900bd2a52eca74575f7d3768166681fd6675d1b1694cace64150c95fea35505adc46646a809fc6744b4efd31104e57c26ce8641a205da40c53481a5c1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d5950aaff85c594247f7bab786f40bba10a61cbc096bd5cda5cd011493cba9137c23790b93ca224dc7e7b8adb6511450b4c289d224287d5bffec685fa461e32b705398c577c694f45bdd90398e9730dac2136aa1064d973f2c6e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he1e1762351932c28b6f4e1217f8977201ded7fc07be3fb82670d01e14f7eafa5646c984bd09bc8a98c86382121a47631ab6f03efd382feff42f2598bd72a0706e75ef838991d2bd9df061aef1617a7b87a5d8d6770906be0e2fa7e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e784059e4e5beec7e41757938ca69a7c0dff3c97f5a73635d2204216e378b8d87c9f546c25a90912d2c79e9e4f0a01370e6496f20f128c7f86201eaa1b52e937ba5b64902a80becc25540eae70c838cc2e68824e85f2d9654219b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h182aaa29eccbe85882cd7213304446dcb5fb2608da80f3a5a7ad7c00a0453268c84384d7540731c0b7bc08f2b1cdf60ba1f99f1a26f4b3d213b3f2adccbeb0c6c09e1fd41009f8e0ac9d4fda291396eb1f6dedede10dbd653f9e2d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b8ee8382917e84835a86c44074442c7f2060361b84c52de0ceb5313339bd3a4c361c39994438b4c566471ea46b3e09adb257eb66659d78662c63399c30cbd344c17d0f745f335ce24f727b1801e9b13c414d9de95baa0fe59de5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19c8fb2ec10d596731647d857806a0ef7e7cc1467ac75a7fbeaa1b087355a5956db9709d7a9e816b3d31708c59d3a7b60ac4fc5f1eebd7ef477bef157f19966cf626a3034dad6dab494c8eebf47e2daeea4ce62fabebbdc625d8da9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h171076fe6a9f1060f59caf705529d6ad1566d87297865d70733c1268fad6ca7f4eb33e27ef764a775b2b49ea07c955c9583492cfdf16979773fcd8a9c0f2b88384b2d1161ef9c43dd93fd217313645a6dfa827929aa8bed5c41a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18077a5c46506a675320402436a5d8306a957168de5e45daaea86659eb72c013142cad9ec51e452e7c06e21dd29a9588a851a0a74397d230b49b67d37f52f86f18a23e02d274523114c73b10ef04a900630dd6b363344ae7ffc05db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h70e3766f1b36470ffaf754a8ec58a734fec1eb09c475ff7e32d670af9149024bf7c8e8644f42bc6d7eba8940ac563ded1f33d5b46fb8eed7effea3f1d9d0f20fd65a68301a0d1d5cda722003c8f94197b845e1e856ce7c5ef89822;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b9d273d0027c81dd78210b18ee55c3c4f1a90e71318018b3ecd3b2159907d612aef27db1f266a5229d0f64898bc3643559cd18258ab68f1119e4a9826759c2f9514c260d68577bec4926da7e5ffbcca99794f77f6a3d1ecce4edd0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf605b221d12f05ebdb04919525c41c7e400643cbe2ca8c85e2f5b7edc69d962d56c75f2db29ea11e24b9c28756c08ca6758e599581b7bf37f28c0dfa585f4df4aa36f8cac662b574eb4cf08747a96fac61b9e652a85255956e1df0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11733da27e599cc7b3ec757fa1467a15994eb58207cc15327c4a55825fb79f3f9849d24f969015863ad7437ca9cc6fbd778e4a3c67e8a80612b9c4a3299d2ea99045552125214e2c6c3b6407411c2b805636854181d65877b7a9a17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d316e9bb34367c81c7eeae8e183c9860a8539fbfbbb69b48bb003e8995bb4812ce82ab139dae8095943cca0979117519d3715f184234eeb409d0c44a3eb04ceef714a45a33ef3c9852fc2c0d97bc5b792b07b54f7a9aa5aba9dbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h29573d81ef62cdce6cabb50693903aad802e9f22ad1f8408e02173b915fdf7936359fffeae8b86509d6802b31af2ac58557c1c90c2384441b313d47931f0c2e8de9ffe92db9822fa05b3804580904324ce0e7852025b399cce4855;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f1b528527c5c8f6143f137e333b0245ccd5caf2073c889baac3b87aacde12c281b55771aee6805d479c4fe16101b2dac16cbebeba403c108550a3e178d801c2b13d80716abede0763bd893c01ba3b78426f03e6d6e369d552d379d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc7fce7b9372eb2007584a0119cd37ff150ce120673f404323345c977889e0f7862b2a22fa54263cc3505a011deef205a06d1313d440ab84e9cb6c775ea73af5bf208d259e2dcd9802a4f48b437749f36b59c4ce61ede438215b91c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11b113c828af843d841a6ed9dfad405198989fffb36d219522daa18a5f7b7b77cf408df3732a6c14d5af2ffbd2f4b3c65f42d38f64e03ef76195028b9b7961ff66a70ff9f9cc9aac6ca7ea4208e9c483401d6effbf0facf75964e08;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb341b48a54cc1250eaef2a1db37dec2729b8268b9d12af286d8242966ec947675572c462b05d3a244b077dfac96666aefbee00627561d4c7adfb5839f35f14c1463e58ed218b481fe0a4bfc8f40c691a37107c78575bc5f8b17003;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h872bc56cda78bb30375c01190769616d12ebdcc2185966ba1ddd2908a61395cf37dc429d0df43248374c8fa1e438e213a40cd91d3d771f357d755dfc10950ee9c0285b835fd69b674b393537add402274bf71b01b10a599f911c8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6dae00fd8827099953ba5e57ab88ff86dfd6fb235f727f76153d31c7f877affc5827f6c014ba3d4f4099bcf96d727340c2ceb61fc81e48724be37df16cf8df8a2a371d733dd444e599f637f5c2deac06f9421f66c9227b6660be44;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17c52accb023e088a535ae592dd8c8c589e934ec4082ead71f5d28c44933f98d77afeb35550a57c74a161ae4eaa8bc1192296792821487739f3fa70ec4df9469ae8bfaa38de390d275279dd6e23a59e90902aefedbf90de23eb814d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b87c8fd9d6fdaf5c762603e22e295cc954a5cf6b10f2d7352a6f7b94532448fe035c3162665327e3347c0d93997a043dbec569ccb859a8c5ae28f710e59b53f0cbb8f2f14ead2753c6d03e7625a7e47c8ada4521da374f6a374c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e7dbfaff85faed0a992d9355ae3a61e735381ff57d3d58917f6f7228eb21354493603ee9d6e27dda139c0dc168f203b4cd06d8aca5019167a8a1288550fa813eab2f7dee0afca688313d8f0cbfd24eb7e90e437855c43883bf900;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17132d5aeabd79368230116e0ef92e0d86e09ba8fe0e4b2b2a9d211fde2db848da6a5b2502987e359f790249a878017c64ebbda0ef850b16050d7076434af5262edb481b3b45d892b567e5e5f42b9f486fa1260e9fd11d944657a36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4efe6237c0dddddcdce6ca52bbca8e2fae0dcb38266646fcde6e2223fe74c1b4bb48fb00be5ca50a63803e2350d2a8a34438b5e37149a45e89d9dc4f1c79e961089eccd7ca13694b437c72648abadec90a7cf349b1ca96d3a46501;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10a8f8a1c86aaf7e9edf4f2bc1d0179348ebbbe8f65de272a69f7b3b4cea132d757960d7688d05d91c9f50d6ab98a10dc8d24b4d668972152ca770de70db7e5d9ebc6d738440f907c7117513d236226f78d3e50823d10deaa2a6bf4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97d089c38c91090ef992373f7dc56b59b86335c0502ae8a638726d40bb3c1b28d16be667999dfdeec85fafb82b7a535c407c5bdd5300b986aab34a52827ed75b086d92f245f8c6e919a9f2176bfdf62baf96ad6723c6c1bbcaa1ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10abab925f204827137e929bc894c876caaefffc8699f3f42d16c863dd598883048f9f98075a008f3a82b391cb77db1df71350aa666bb6bc692c36fe116b90bf9277ab7a81bbc7baab9b16d1901b1653e17327ed1806555d789bc74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b0596c8ca778809be27382408ff54837937dd80f38d105e7df015bc86352c210c3393c94042451c93b040d9149b0e869a5f87987975700197cf43bd9f721a366b64fc31f07f4ee2abebd0e244dc7328cf59315e0dc6e049a54c4c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ddfa224b06af6e2b4b7f522c0db1472a27047f1731674fb3193753c4c465a9d4015d88b2f3312f66540d8e4f72962f07342acc3db6e33a61b744ff73b102e5500e1784f49b278523e3f20dca8c02cf41f155e446e98b7fea01f0d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d7cc19c52f55f2923652f218fbec352b57c5a98b180cb67c2f6c5fbcd3cdd2c8132089f333a14544ccbb23ad870c204233bb313933ce113d1f49ad8688455feb477fe077f256dd13951b82409f485e529d766a14aba46f96dd5aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177391d23c0f271099db4906fc0d650400d0476088bcdf009e07c0ea290195d529a767ff78861379f771618f90ef3b4a181ebfafebdbd15f0699760f4ccd7579290a22efd441f1477d7af5cdaa0a3456f1283ee06bd0b11d99151a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8b0a5fd01d83f60d1182aa58aecaf060cbeb72210b0a4c854a1919fb93bc54e4921b91b62f5c34586f734a252f7c81676ce203a2ba481df4f296e0b4e2d57b59b35bf76c3a97de03f68d9488c40b65e0f40178ffbd0f807d76d9bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d3606ce094f59e036d644cf584d866248686ec4107698353e69a5f2ac33759cd2437e187e003d9ff05716411dd69c5e73d81490f279d00b670b8ab9cbb98b5ec3d9ac71a167aa0ccc5f35cdca79da3c9f889bf276673c745759cd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd57e649ef30210c7378ea38a2355ed7a577f6ffaa54299b087252764742dd4d23b12112374e0fec2813d07814248577460849c54abbbf4b3dab3cf42cdda9745ba1c415f514872a90f36e6dc742965c9722758a34670e4de492408;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h71b7a9c6f59f6f0c0a23ab0d3d74c31dd396a29b69fab428b819623d3989cf7d302cd4f95ce1f426eec79e3266bd65b73c99411d3ec234b32b76e1c7b69e9f0b2f5ae1050ccb5314ca7a64862910f8edbf62e2145c9e813ac8b263;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd21d688930053fbb5b1a3c17831e13d16ce4d0dbc4d1b54eca2d425b3a3e06cb6464c09d1085c76001440d25622bb4bb0613ad9415f07c35bf20b3557a07384f0a2ba900ecd9a356d989debfe328fc5a03c9a2e82fc7ebceca6ca7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9a15c2eae5fbe07bff050cf3083bb3507243cadc806ac21afc48d4b3efb15454fb8785c12495149ea76109e28f0777aff298fafeace4606223d9af4b8e7bf7aa3ee75c4b22d17ee2c7f7e8ce2ef24018b8c42cd754cfc8df0f75a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h86b3fd6235d71f70bb4c27764267ecd6ec2232a2d312003aa2161aece4fbfddb6a239a7c4c6c7d0f661145950d1009157dd0d9e0e95590012ac961d52b197998bc370f31fc52b51741f779dc88f57dfdfb4021a737a20ec6ac75f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136865d51bb7cab5b5cfc2293b734cd3ff3809afb743e352e20c75cad954332c4a8abcad2872729ed14e72bb3756d29a790e03af6b231ecbfad4dd00a1a3a849d4a0c6b574a1f8a6d452cad36a998f4c4af2bdf3c8b89c9ca31c81;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c54c9f4a34b9c6de72bce1687bef3f9883317247a19e5c447efdcffa0e51d5af54ca973fec044e2a8176469a5db1826d68b15b1fcff8e6ffaa9784432ff1d3274b8edeebf764e4aa2c8044f09ddb3b79ece3a42394c5a51771204;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3913002c0b979e77fbbd4a6e53db3f69e94bc6e0e89c319c0f48578a3420e9aa036803f9f53fcd6f99a28e53e3de2aedc0125db6bb5d57a7c79e000be1a8c661ca9043144531cf772c4042ec79e165ea2c0f6d5deef43a9e65c1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h71db3ef27b10fdc7a52a7300da31f10001e67cf2f3d879383e80672fa96f090a61bc8b4f2977c21f6233a92ea551375581ffba904a347b61cddc29ff945dfa4b805a97fa9aa6bdda32efb249f0f98314b661b393d82a1fdf17b002;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1afbf9b0759e1733727feffb67ebd09d43f823195b9b3a457cc193fe6c29064986d44cb0a9371005121d7ce914bab82fcc52bfd1f61eeb8d429ff98eac01bef3d808558605d469225b1814677f15820690904f4331d6d6919b95ae4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4d4d47cd268858d4998ba26ca585f02b519f7ece46081d485ab360d3f6889f9369d3b998af0d5c7f55693521e73aca37badf3e2835b20399f4bc681db0eaf41f61d4df7f029f7b5ffbf1beb9f124ee9d85169d79eaea8d6dcd2f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1963a831c54cbb7ef66356879118dbdc53d20ef9c2fcffb6159688c4cf659c536a5c47bb22756043c80fe360d0c8ba0d2c7281b4d5fc758e7450c8dcb2b2b1cbd4eebdaf26e8bb245c5d649739ed6f4aaf2db84449753b351a4d884;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4092cf2ded7b733e2e2a475e5e81f60ac83e7d6785e18f4248e05b51b879b8ecbd7802461d7237f5ddfe0d684d570190ef84669162b38a1869cf279c8c62428816ba29abf61c7256d7c8c4838f02f607bdb4b2fc36efb36aa87101;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h67b2f44cc866e2c7ac3b65b4911308a00436417a210f8a4122ad2824210f4ace34d2ddf7057b03274317acc058365d80d338b94b4ea41203f2f1dbc47aeb119ee99466a2ed4c91394612e466410b9932e8afa76e92d38dc41b703e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3d55fe8e21842c0cee9c5eda17327b23cc9f0a366ed0b50ae7cc63dde9e856f1dda3e930298d72446c883b28e7be47e2647bca95665f6c94340a3e0009fd8a7c01d61fd24c050cfe6a502595e45581bc2b3093c8cf2681fbf4e6bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h54dcf45c999bd29f1b0cf9f634a6d5814ed0bc3daa2331868e27baf57803f8b905a2d1e439f548857e700062e798861d57826474743289134de4549c9120f227dab2cd6515c0eb826f9f0f103b5a25ec0d88cb324a52f55c7aad96;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5319c8a72f38e62045b5ecb9f2554a9dc8902fcddb95a0ddf55fc841035249f0d1b75a065af8c44567560a0047235773bbba751b55a21f7f95f13da20e6e9b0fc9d5f3e1ec2fee5d3395108a29bac285f2be04387ad0c9e02887ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he46c0f95af745d984eaa4a626858bd71a19a51450110e83be897d718006b4e058676495740cd6f9727dae0e6043919ad7dab013f36094d49127ba319007b98e02479efcd86ed97fae80983de83297c158bac6effdf483a5c3c03ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha2a3b49b1f1b3d226bbe699368e936840b5c1c24682cf8353a06821a5de2f9cd46a6a600bd27d0f77ebc1f30e6ff2ad5409a371a7e73abf165450cd8741d0b7dd63310af48b6bf78f64183181996022d540afdb47cc81abf59f51c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h80e196483a9ba6b2d19f4de85dd02c7355eb8603a83d2d762ee9b88849c61afe6e2fd03be8da061ba8e9889025a50eef53912aafc69a62b0033f2672a101162f625c413c01d424f8d2d49368fe25e7f475f6959b4eacdc5667506e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5a3fa97a40b9d25c5d1a6ab23df1c843734be2381b342f15aa094c952fe7a9738ec67f9b7c8fa23ab4268426b3088279a43290abd520b5cdf37fd53d7c2b0aff2bfefe48d0185df0c32b47ffa66b3f91b0b7679084c3c093e1c422;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h90ce140247ae28d27cacc4f9f0b9a0d418ea09c6a1470d7bc1daa274dd052479c66cb6d2a126358f9df66dfad692a8f4f97212869e7cade538ffd7914f4229c4ac477535ad4feae8bf8089b4f7c9a19fef56e428fd88df1c3878f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18bebba257a3a4d6eb78d7f43b4447fb1c5cc34cf5bcd55aa386abdb9a0229c79b578c79dd6b54e798797afdbc2e19fcc33a5ccff0d1032084a5a0b204b03e38a96f98085271ef44fa4501e8e7c026358b4ca28e040d8bce8f42e17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c7154e2216eb55cd3115780e9523cc5ac2e456aca3295ff92f993da0771e4bfda06c0445695679680c958bc38c8b609e7aacba169025e5660013b5a373bf6e9017e6e36103bfd16302ad1da5104ab659ae90bbb1f9b6e941e23ce0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a972868d050db144e459aad76b4641b522fa79061f7317ca1ef3504c1b08831b541c491a6283487a59512e2e309af239c2c31fb3352e21249bb0adfde8bad8a1b75822679729edfe489182fbe22efa1dc16c753a3c5a3cf93b8211;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19ab6069308569f78d8cb75eca99ec42bfa0fbbb393532859496c001f6a99c6e59539a9d27d49549e47b0051820dd8442d8dead85ca377b22853eeb28dc931dd787fea79d2275a7b6f3d1d7b05b2a0da15f590c5fddedbd96bcb8a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1af4c3e0ff2bd702b173184460dd59428aad41a3c3074dd67a5a0bb63ec49c0bf0f53b747ad833982d29e9b90e37da4ef71446479c2a6992d63447164d0d07053f3462c2eba3edb02209dde364499b353ea6bd5e7f1f3754079497b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2e34d41eb53f7c6d60ba2ae83d2fb182000bfe189c91d93ec6f935aaa411f1e1dcd11aec4cb812c2f70a52013a1277d42b994ef558a13619b114cf14419bee6a09f313edc613fdbfbdcb7d9f684ebb1503e0582b73ee4e7b090d82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a0478b4894b1d6c86bec59ff6b7bd7f9eb433a4c2418f369deb9031c659ebe8f8fc778c0bdc798721f8992637ef4717bb91d2053d458f196bf255c134824221892583405086e9ff50e6ff7a547135be43c9712f8673a1e463a1082;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5b50ab13386e1a480c880809d5edf61cdd334774e9c9d6eaa22730f212ea4fae4961cd6345ab5ff7b764fec6fd932eeb985095fd4a76d5bec0637eb946f3de4fefb1811243b6e508b9eb4106db5f668e28b8d5c66389f22668efc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1258166c7dcd9c2ca3c306326dac1df348ffe4db2a693a983f17830f23226db9a0d905e51ebcfd05a34fae3f6d7e380e3c995a4273129073f2dc758622a773ecdc7a2d543f41f4093709c1e7291569a09087c4194c62bfae462b562;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10c88b2c13bd13dc53215ad7c8fda9620c326857ee1bc8a42f8e6048c130d304bd70d20772f04c577e6d15da81bb3c8002f6119dc350db93a0d6f32a1c049daebc95093aa188716fcb7698a02a5c854dfdc5e0ad1f6a503de88f118;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dc41d09e41f8c4b34152a0ca89b537283e478feba9575e2eee5b88c2c582bb47c76b2bf847157460134be87c07d0a6b9e65beaf526bd291b912a5eb6896003a7b84431a2b5acc49609766d3799e636d687119a5a72adec49f5943f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h85ce0a953cb04c0dd708126e043d8f67165b492c1a0f1f2d71d44cd5c4b30d24b39a37ece4305c85110d3e8dff9341f572258c61acc14b7d231bb728121197baa9ebab0880bd6ac248ff456386b4bcd8a70308a69de2d4d4d36723;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136fc0dc441c3ada5994779c9773c5cd75447129d1eaf0a7e149a6a8bc746c9b2b8d1a379cb183e1f8f4b3bfb8173e01f9340944a65c36976dddc00f99acb46284546dce619913e060cf8931af27ca8bf58af2e942308145b7bca76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h164410b4ee7c6f279a15370047abca263c92c233d951d4a684f23276fdbe65ebdd098d742adcb3018e8b22a3ef630727ccab10d1673b481351c6187fe94b649d27201f54298ca5b98436eb14abb9e5962a219ca5d0235c4ec75168f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h228cb55b07a38cffb71e18487ab535f5b34b91ae531feadee5d4033472aeb98117e33bc4f56dc8195022da54b244b2ab4d8a13431f473e15a8aba7fa867b85d02aa7d652689fed00e281f4092c82318cd18999618fae1fe52579e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h136fa10537be1dc4db447bf88068edfad628485702b36483cf8774cd5496f357e1b3455f855a77d3cc66d9c0ad3bb8db367300880dc594d8adcf2df96ccd070188d19b1860877ed00337632cbaf9b22d7b19defb693c53cbae1e697;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a7f48826638c642c6315bbc2adf3e1847b8054c3a70f9098ef18979227df60d38b2b3cdf2a7b8ff56b08dfd5a03fba0557102a16a4bea2ef6a29ae461eaefe8cba5e2ced1e34a547d5bb35ccc805129a16c777193147030175a1c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11009e4cad29649f5c54f276b51320e657b3e684c4e72ca4ac5aa4eff36b64a0f8b53fa11f09f15583079c71e36c6ef993bcfe552b75b596eb060f77b9e0f3a139e23e2d19e2d7ec843e6db9487eea2160ad9b2579babd8e2db2d39;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1251373bbec9bdbfa86c03f0b7db59819c66cad622ff098de158442be5c74454b909e6797a2d70ef4edddca6d4bd29ee68114b64321586e802828163d2ac1c03024828a1cf2f73c897b34b3bf1ddb4be65ef91b2b19f7caae986bbc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188ef3a8a4133343f158050f02c2305c0f3f2d9d50ec8eb782c3f917bb23543a579555bb82c561e3da5e86090e7bed39245193129068b7661bc21c7c85a98c5010eb53967120a231ad2d09404c8be27065920a4399773f4cd3a339b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1671c4f0e1703dc30e6c1bbdaf185759861863cf450438ea3c35c8ed55c2bdaef715fba288ac98764ae3becbeb02784404631a59cd97324570a62c638c6c8a772caa371d472cfaf669e63ee4d0135fdd69b2a5795cf2ad5f869aca9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h193e7c29452ca9fa72dbcde7637a4e7b191597d7b720514280e0eb7347a54ff2c51bbaf15286639d3d3ba0d8de1941db5b758ae5bb082180800cac4f7a2ce6c02feb25de76c808e5905e0208be360f27952a04b5ecd12000172f3ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h59a599bc6946d8a66cc9fb0870b9f13eafa1bccd6ea690ee02930140353dbee44e436c68589a180909a62895ae3d10610692f5f290eec5205a76fc0b93d7ae4086b54600c63027ad9299926a2592cd1d52e449aec71d75ae6c201f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de95fd89f708eca8099bca4ba2bad5b8a88a207b67b204502fe573e93d2448ae183e6569e7534bb207aa698f1f503df8b90163cbed6577f40bb8eea3ccb7c71e62e76b4d132ac225beb7300055f1ae5aab4850ce70d6fdafd73a74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h171a715e032b4753991c31d5785db563ca9c16af7964474e78a02604c0583e9030da6f473ba2335b3b2155c63c6d8d350d4aac7d0a143db83cf087b44de159b8ff973034c37df4fae54c42264e950929dfda745b3bdc15a21b177ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111a5f51092a624a062228139ef3149d2b5f39708206416afb68749a3af2f2a80d373645433603d6bb7c7b626edf6ca26813a0c9e85b80f4a0157faac4c5d15b6bc506582dab937d104612645e0b3231fc01c8173d4ed7d8e9bbaf3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc1c7a5802d87d6cbd19c4cda19c9034db56d81de512303b19fe21512ad60e5e0f619ca9b07a3faae4a851a9ae4991c4c671b5ccf1b1e0409128f470b4085ea8101e2e423f82e4e5e934d7c127cd23aa09447967671c87e6131c7b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13f865a17eea4795f8a844d7553a678d4c6c25513b66b829cf1c3875cbb8cb18a022c9613e5545aafbea4e58c3d2ffe0aabb45740b2516d4ab915259e198032f1a460bc3fa5fa0841fafdb8ea8c4d49d83c8d388865254e48c38689;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h764b228bfaadbac96080344e22373fbc43bda0cc92c733afaee73702fa49aec5dc914b3a55f942ef6e9596b0ec6af270f174d77f0dd14d97b40e1ef58d00667de34af34d12595e5fa3ba7dcd3694188fc32c77e468bd4b281f4fe1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36fe3ffc4df0a844f7483f7b745fe9dae66c8365cd8be055a08de725eee4d70e3c547c5374475fa159641d65bed286d62e56acac548b09230b9e5baac71744047c39d3f98880cba389f3d9589c278395f4fa15c641d5187e462334;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12e0a1e19ac80e55be905d5172936e8e34371abfd1c9e9dbc0c808e3baf3448372b755e6b42d7c4d52882d1817e3a1d5d913217c9a869682f96f8d707dc4cfd2d546fabcc981c21a9310bc75141617be54211d800161faf4e22c35f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbba52443c25dd94b9578ec1c42ca28f26103763648ebba2e7a2bf8cc5725748cdc74a40f879c8a2b4eba90f868e301aa27adb3ad5d3e06c8df10bea3e86a6e7366be13316de6354ff9a83bc77925c2fd28d7e516e9681c32b94f0c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h73fde6f9e708b61dc0873017cf96153c3f43a2a2f91acfb9553dc121a50f50197bf3b1e7dad645e860e3d2a5885b21c2421b2a93983021b3118159b44cc44cb0d18f957836b502ac890a4e9ea1372c8eec61251003fef44dac30e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab6fdfeb7f916537a5fae9f1a698b13b10566cf6e9084c6e7a5d0a06fa35798c5779d6ed6473ebd63841abaf4e292d68316e240faad721af117e7ad585da8d9ee3bec50f4b4ee9c68caf3981ef069a36df8aee3e7d274428968cc1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8ac767370bd55d78564bad91285fa3602ff7b11c2be39bcbdd3266737070665a497b34ca95ae4aba414b87a4e7db316e698a0405709038166801596dabef7014d80e11a2e864deca46e7d585b499bcd9967399015d7d521ae9b89e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1008366b41167e59d3b15c51376bad115b12968c54b20a7914c486843097922c517f79fa2885a5c01b9bc52ea607219434684ac405983332423f0a8e097226a57f3703c72ca5ecbaf3bd2ca3ff3d27b9f111e6f035351dc27f072e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h878ce52c252b4a289a70e3804d3fd7b23de6d96fdaafade75a5e33174766e102b3b1c9ca6360746bb63e4dd22d54f7c4ef2ed02597cc0bcabef505dd1d43f7b5f34b6c96232738d4002bec5e2029306ab05c1d2506df7cf98b673c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he412d43b70293ec72fff7bfe9d52516bb03c9f3543faae5f8ace056c2ccd2df820c83a083a080dc83d350dcc54746e52b74410414187c9a7518c291f915f0b41933736193b568d95fc99ff78c28a856fcbe90851ff7926cabcb3f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he3afcfda134f2377c5909063b9a97fa42ef52f732cea5fe00af04edc5ad8f03286a01d791c43156eb68b02b80c84344a7ce08e2b0862ad343d1ce69dad6dc202732c148a4e54a6e47ed218dddeb84ef965e07ff47e1d86b6179bcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1024950ea3d12d9b4c404a15c8d054dafa857c94c9be85df84417c9b4022aa36127d2e55221042d6b3f98938b968585f396ceb55b88716f45955a9d331b601bd058cf9dd6895035cc1854e111c005a728345ba0321a18a75275bd64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h110cc732686116b98c5f08bcbcc5b7d24ec0a5bba9c75ff773938c2966dcacdd51def34c6a329bf7075d3f25143afab1372cbef220e1bcd1b11027a28bcfbb0ce362923564962449bb374312aef432d7ca017d5c5a3e7d55350267f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2400a4a0f71445dfa8f78d7d3f2e8061286cc6a7c487c9fcc9da9339505345ebd07e256753265e06267b1a40ed20ce4d118537dee8cf7a3fc277c71c77a364af80fabad8e860643d9b918aab937bde1a4a586bc97838b358edb2cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e04213106e9fddb10715b3d6c9efd81fd76e662e5e754ddbd5de7afc8bda1755b0ed85d801c7b4134ff840163cfebb1dbc9959724549859e737f122d74c78aa2cb9a19ddb3053e6d7286785be0dab9c64f5694d9bea32921a382;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hda66f1d3cef1c3f18598ac014a09f37efca5c3b4e3210f4a01b9c7297d0326849ec67ae4ac55e416c9f2e4d81c710c85446221065a3b0e9167f55c1c2beb4745f10f7957833b718b847f06c0d8321ac77b19a05e03ff6a474189d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7b80063749da18185bf0ea8b0899e5be5d2c9e37e5d158041f3decedd87a2facb0d0b13f4fef5239268af3caf2bb0d6f369e635acc6ce6c20c116cebf102b64f986d251374ab460ec417ac6be211b11ea6fb465fca8a91987ff6a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6a3a1d12ffb98d6b8923484547ce4767f0a3a32f1ca2cd962f01e75355518701e51b12616683292e359c2de0171e40fae91f13da5f05881b280c1032fc7677640fc7021b11459a61be4c6a62718b2583394e87f47e33788e11ec11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h501ad3081bb4eaba05f4c8b4e73d7b6a6fbf545d17ebcc650efefd72a12c77944a64bba9d9c8de05eae361c54024ba3e4bbbf38f8bfdf99f4fc9c8c9f4bd5f4dcb28acadbcd6745f5866c6560cc17c9dbd1f9ed10df1fe1b96c4ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h188a47816a1e91e204466d03744d3ce5f53d607aa81393c4cf5355f2b201ef4bd48cd99e249e2b2317db4a1bf0c076f0764e18508707d887c6b2a5a1cf2d81f538dd2f175dd4bbbf74d2f2d142bcc8499ca7eda8037f74866ce7231;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4dda663502584a5700c11b61eabefca56bb7971e117e02a2c14267bc9cacd8014cf76c89349bb8f1de486bda04ee3ab945b0effb080cd5706bc3604a9c556d32c2c844b7e3d365eb891b3c138830d0d1b99dc36fa64681bdd24cae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc941c39da1c4534a61e5d7386c4dd7b11861380fadfa3a6257591c28d8d0052cdf4f637b38c92bba0c981cfaadeea58d58dab7849ef2a04ad8d5c7e998d44975e7ad922b55a28ba31c978235612d417495fd1e8982a865cbf02ff6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d48d5a6ab6a10e3d8c8a84628502ee3941252d636d7231960377fd7478c9ab6a228bace9a4b14e278c5087e8bdd28126884350e641eef5013223fd5e6df9b9d34832f3017df09d3202ecac0af5b710ff93f8d5fdf2700f9c57e8f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca21cd7b2584afbae5209d993a89264ce8b0c520321dc305c97a383e3940845598045a5518911ece49f0d320c137d2249641043bb4f19a2b4c5f82c6787a875ee0e17b58bf11808705f606e14044ca4338b7f99f7bf4d8edb61e03;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb01f8cd058f5521a8f8ed9c4258c542f4e321659b6ea27d24a0a70ed07635a6cb0c6410e64b9c53efd43e35053c55e5fcd4e96f21ff9d4059dfd342528c60d776361ce4cb1d3bc4cdc5bb1b184d58bb5f7b572cc7fee0ffff42155;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h852f7a40e0742a1e2d9c82fe73ed5da7c9a51b5026d8976173726414098a8f2271714d655e8cd0b11f7a124b25c8e26a47ea2dbc0af6d750f109f722480110d1a01e6a6c4e3e00c170195ca9b3131ecf7f83aa3d19ccb26be7bd02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13a64e88db7176c00fe360057daae678f59bdc54ef82da54c797389e02d0bc9b4d32ed9f572696c0c280e2474a74cd471397d54267e2604a1c5cd1cf93f64261c3cf74120fc25d4f51885b0b5e5bc6a0df49b0c6c308ece95df9f06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14ffbbf4dad1fbb3dbf584d9d79f27526c02925755778120adb9c933d33ee0ddb9769efebd2f730d5ce16fb337cb36c295e7492b38a3dff3c4fe1e6ab3b979bbda4f5295a0ab78ca04772e113b20c7d5e33867dbb0e7e296744d632;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h74b1445f1175d119a920310b615ea56a7dad0abcb0543563f2fa9ec86a3ae408e72444990bf543bfa12224efdee4a73c5488d0a51731a54a32af2850a6c76943c8e32b13be897558d2806372c5cddd5fec249ee9b4cce1dcdb0683;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1373aac4d88b07b99d48315f5d8feb3f668ed3b8aa6ebb5159f8063726831f84f3575be43bdd1656235db87994ed002fafdc135b391192153bd723aa596e92afa1c9b13f2aeafbec96c0ae2107c175366a36140056ca4340261ea76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha4c3ff4b59930b5297f8747e26e62933011d80a9cf94edc9483a16de6a64baf7dfce72448a4585b820473d9aa8df1f58eb262bf39fbda894bc7fbc47df66132624b688258f8c48d71ada71dbbdbeaac727b96f4c0d29f814d1ebb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcfd1f72e692fe228c96aed1173695ef6ac4cd68c3a1a016d803fa82b567eac1e95bacc3a922086db8cadc21f0c05c8dac71dfdeb03593ca225e5398815d771d59810c469683775950194c16a75a7939cf421d114fa6d18597fdc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4b0b0725dcc0447cfc4567a7d158e7928c0e0dcaaf127ca6a868ca370a18d3fe39a0d1685928a4c3fcc352482619f1501e89ba4b534a2b0c3797de0a6d61ba084fe13042386e59fca3ae81a68e7519d8b6d56b29ceebaa17e0767b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d7983efd7fa4fdb51fa70414d90a85c1f37c7f52c37a88c353cd52337a088d16e724ea715a219dfd7a7fd94110e6312091f93343e6e7ed39072e2de69f0707d6b9d8f6c0352c0372014276017ac11d50d9a1ef3126a812c527f4f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h92c7ae92fbbffb7c844320ec4a5238aa405ebca0777fcdc4655e8e72542515624fc925ae638e6c77bf01235f617e6698f94c1004724705ccec01e16736b7d41f8e9ed53aa28337abbfc3854e3d6ffb2ca550e97fb19526611d31d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1619efc64baf2ccac87c413b3ff7d326815a94ad108c84c2ff06fb9304bcb6cd003e8c78e53e81492d840d6a1da7af4f93be97332b23a009ab30466a939f82e46ade3dc6604e728d67ceafee4563006741a0204bd263105ccfc06;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c4cd4ab63fa995fa11569a615a575325c3fb7e927043188239778caf06a3f458874ff84646b1b07a349b66c22802c0d40c3e3926ae51b559e2026e1bbf5585b7840899a93360abd42b6b2cc9f4e172dd98af184e4baa0a16cd51e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h421eec443cda9a49d4e4117f36a9183b945b8cf94a588dcaf174114ab23bbcaf609496a9b67a8bb3c7fadf644c88cdc2b123905a905e49b11339260c4d828efa45c2b8575daa0e6bb666596056668f59c6e1edee4d26337bfe2b2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6b9dbecbd183cbcba4ef1c8c9fd64ccb879071cf991688cc95dfbbbfd75ec4c2b4eada74dcad38e417bd4898a55cb45c5d091ed6945b47cf828e48b8f0d6ada00d71ab71be92c0d4956d79d9f3bfdeb3ab9064c8b5b9d6ee48a055;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1642c070eb8c970ff60865149875aae95359d2dda3215f81e44308bb82f147cfa43d04564ba4cc285e8a8b5074ccdb7f5136d6281524b41c1d4713c7eac2a901b1e86f02329a87da6583d071cdab4e7a2bfcb871b5248d96fad0f45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb8dade9567a38611b2c8033c5a8b6aeb579054a8c0e023393791978b314a362bce2bdd01e65ff19261401393ae4a3ab2ac58817d62204fc182f5670058fae878db5f3667b47c1f35f81e4727ba5f24d06c03af0c670026855138d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d3042647918e11982cd39dc471c0bc4322f3920f0754e982939618c0a1c1a3697855e2bdd3891d4ee46518014fdd4908d4a20d3181efd4925d17da8bacf35fa278ad2eb176cc5df42e6485b280bf4b97630a473901a227e86c669e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbbbe163ee994a1f89b203240a3e156b2d0901aa2eec815c867637aabd8ec02dfb86bbda52dba1aad6400dce5acd506685c227fc0fa315745043dfef7c3da3f62e8663bbdb8ee89771aec0490c24a676d67265194789d3b9eb6eb5f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f41e505337c4c5ba07fae21a2bbcc1a0ccdd867f75c33b6b457f0e085f70e2732803a7050f7a9274fb782eff20b34115b27dfa601ef462f2c8e1832b18334819ec97824424efc3d22f9d44fecb5c331475f15975878e8edb56839;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf39cd7e456020ab7a130af807e91ab06ed23de9c78f4f12a5f24209df41684b6fff540afd9f45bce60f634266757be4b144fe6502d7445e7ea33e3b9bec8b4f4cd4f1d51ec8dae853f9d46399c9a7577825d24f48d075a1905ca53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10456341cf736d279cdf648db6d4842bace2d766c3e701427a130c294d63eeb188040e3dac5796b294bbd8ff27cd19aa22322978a010857e6bebbaa1f57f78b852cb00b901d5e7fcfd30781d04c7dcaedfd154166fefa8e14b6ab7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h122ad10076ea7f24134d5fbd223015c2ef3e7e3d25def53d421909cbcdce0d991fce55ba8bd37c4c44a23dec13757a28410aa03c60a9d5338319f8e2cca45b4cc15a4bdc6e7b5a69f3d9be67b5b2b8fd3bb6eb97a78133afca5ca49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h469f258c83c13ba0f4508778aaf4db4155962d67f12154c49a990095881a8020103f3fbf340d126a6fef46d0fc10a6eea34d399c41dc1c8c0970e8758844dfd726c46bdcd584ee61d65bec91c4a12dff2db55c62368d68bb6e9fb1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114ee16f32d504fd82d23be9e5d2c2695a5c6c2bf1d8a5295c86e63ca803bd7439e159651c23cefc8c7221224e6e4d5faf273440152f201086b772670a0dba20f238235d3a51a8bea61fd7438048165f2a75106023f40c1dba9331a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19b9090a8581b1e4959851f60b7f6801295d1172f411195656246dbdd9438b26a92bd91faa2c79c6c0b97cf0b74e1d09afddc13d05f0eef93aa8ed25d9d50919c001a20ad6cda0c54e4d2aeef8504f1b814bf5aa5272b5e45bddefc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1549dba1d7b1715f9fae842f16d50fcc6eb8c1d05a330ae8b87e4db048d06c7ffe188f1877adeb2759f954e73cd31c51e116780b7dd9609859661a9293323f15dc9960403ac2d23b78c9f7293b15f4edfe67487370626cf65ed1807;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h23dfbc1066479763f86a2353d6bee109191e07d3d467b7286df3d5cc011f86814ee93cde01097d2b18a7e5686cda0849e598b5aa20ed3235b0fca1a282bbad47dc0c00a93910ea359b44ad53d9c27b5dcc7637a19cae81061d197a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12f13d9b5da0581a5e7255c95e77dfa2f75ef38cedff4dbb87353f7c27cd802c17c89b97e0548cc66e0b832b01b64eb139babb0269a9fdd2e371dd495af6da10c6f4c8cf04896d4dd261f389955373636c1d1ebfb88398243cdd069;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17ea8794866c0737ec8ecd66be29c9afe9494e04d7f38d509287bc5fa08fad2f8d44616162924b5da6eac5bcafd128a7027aed7eb7b2582d0e52dde0ddc4ab2e740bf2a3503e9d1d0b5fe46f5376052cd6ed7380afe26bc64dcc2be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1640c52acfbb285983de76e5aca1096ed093adfe12ee5b75150a796d9c9a991308a5a4b98e5ae6568ae9722a42c210889ad5d1b26f44df693d4720afc988223efbeab83709c91bfe107febbe3fcd15854b1fa4ab411d966f553783c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h137503f0c11a27d1cc4d34d2f7d84f4577c3699ed52cf146b7439067395cf91c80eee25f7f2ea2d5d1cb7404853b97b61ad4552346f73ada715a5cc1bd5d09d183d8b62f00704a555b2522e4885ca8b20c66c7b6e27212466bfa929;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de727ba82c88546c61791cc54985a9dd9da498e81116a3674ca92e8e2c576b29450d910b98b45eef25137b1ca3b6b31f7bf7f5dbbfeca20022ff1bff608c274ff2096e0481274febb377652c4cb6ff2aa46af4b24d3b1771818d1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79b85053c5dfc7c291d78473d398f1b9a2f132c21e7aa00f93d793dd67b1edcdb2cdefb113dfa8ecd96d490c89f97fb0856c87bd529595b6531e4cf3b9dbf35bdd88c26ef18f5def48f135bd2aa9fb4f9920581fbfec13cec85ed5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15744f604b57c5258ccdff0c2d7aa2de0b71c58dad8c9f822e1e98efee3e1e6bb63a5b7c4a2f0d7af544a0c727cab87748f3f298f9628cdef0faa7ef0a01ea508d93a06934efbf8388eb3ab053e4b44d5d26403ed1c4f711b5d7856;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5df6bfce70ffb5c69d78ade3cab7d2ba75c95eb8d385bf230f5da492c2fcde5e936408535ea9929968de1ac82b5a95bc3264582b7c3ccc2ebb0ce745474c00e2a31edfd2ebd2187ae7710ba933cb656886f8bdc279dc096fa4c6d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc9600d4c640a00d6c929637787cb54efe25a788bc8f80972167a2633d5673829bf4220f9383623eed243f0cdf6164ab70838096f6cf93e192137084ec7c012b9e60805d982cd28819c82043f85770d75db38b43aea95623b522a48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15aab86f2bf1ecbaa42fee2d51721d77951288a64760262f18d2329bf93ad941daa8b1c3c23654af164c70c6d4950f85ca783468caadd94e6b715888e74894e118e44d8cc9407cd13579d74d43c9e3aadfe26a1e80009df4b7eafb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17edaea5eaebce42834b32d78569bdccead128e3e54d15f09a64c5c380a3945f46c35dad0fcf9ed49d56711434d320ca96b7a899bb2c948ab301bdcafb386ed8cfabf0acf3ef477f74a0cb21f4022df2311615c111019180a9f1354;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd8326c5e2733c277ecae740f85efaf6a8b4d2f27314bae123158c1923d0119f10180801bcb2a721be710f0f5319e5048c236471ea0d2cda4d3968837fd1742f06f8bb70e3ebb0372e5d315210e33027a120e05317330672980dfa5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6bc4429e92e276f09b39ed6a17a4b441a7b35038eaa72e74d8d9ee3b058add4c2eb29d97193340d620a8be7fd74dc8476960c97cacf197bcc322151785c413f89f4bfc637688349f3743df61d9c949f8ee97089f6da199b9b9c2de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18bb6b70ae8c28066fd4b2cba2684c370148e6c62236e397885ab230f2b87c5699eb9231bdd300d8341a25d57f6add0cdfbae03bf9ef10a262c93ab3a39cc060bd646c4cb8fde76271d326a70a686e8578e90d64f821aef9fff5bf3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1324d3e6f8f12580cd340c1b0ea324d507a55bafde0c26717f0dd55b058fc18b32395a75acf268659b93b315210e5193dec0ee76566c7d0606c232224a1bb83e283e049efd15acb77a740c9172db15c3f18393a928faade38b97685;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6174e39a4630ebfd2196222c0241868dd6cddc389317381ea7804096abe6faa11b402371f849b4d291c2f393f3cb3862720a9a4576f1de111baa2af01e536196b045f32244014362e04ca3a656334ea1f298fdd9a56015b554c01b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd582f7aea134fb9369dfddf1d2ca3f9b48dd74346fbeb0f45ca936c50eda3f09b7b4ae02773052d30b1a322c0c1bfd616e0dc6cc3740a96655fcc1d5091069ce28e1f048dd619e8654ad77a1df662dc1584955f1c7899447e622f3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb2a42ec803d1e0517598fa3d6857daec347f979ecdab95037817d628b4933254111c7e22228f08e967f48a2a95e3f1b7c8f905c59361c22a355e8df6bd6d64dc43a66510e258cf05c67f60b3dee5f1fb89ab4c972de463fcad7ddf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a06eb1b2b5d8f7452da9f3ebf2a18fcd7a9b361573ad60e3fbfb8a7b98b1b07d2ad81ec5004e87fbac2b61f348074b98df955362388a050a9c2a92d9217929da43d6b9b379b33b7a1d897460056babde1b641360d00df300cf72b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h464c0f52c0955dae4425524a41c370d54d5a1d17e6a1050f1706e70f0a56662aa29289a071e105fd2edb61781af1a215f0a87ae14e8ceb5ca012fcf51246b607e371d8c3b69e84cae6b33831c86b1ba743882d58d5fb8187d2de84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1eb2e574d6257b1a66889253809054ad200977efdc01928e3accfed40cca7857d17c669fa4b721255051cb486242e6152a3105f27ca3d5aef52ee4fb4cfa314d47065f1ea2212d309203af5c270903d95ca8599b95659cca81ca0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c5734ddf5941265cbb1deefcafd2fc4a85443748d81b4d381382f19bc6ecc4987518b697dc4dfbe844254f2c0eef96adbda1383caefd88587c9959ede04084ba8055c41d52820998c01f4b82762b7bc199917cd42fe7f247814bfe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4552c8b70c9f451c287e21caf0173275bd8e37f269a24d727efbf01c68b3b331302047805f339a8a642f4388ddfab710f4abb5c9e17795d1fb14d53d258e333cb86346dd132448b588ebe21cac87cfe350ba8bc92f417f228bffd6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12b480be3b8f3b03226c0926f4b7d873463e59583991e500962a50373f83b50ef1d76d14fb65bb2a9f4efe1c8c473256a0127546d7bbcd58971360d725ed289afe834feffcd69f2fae8c6e94c24e9201bc884f55878e5044dcf67cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179957ee14f0bfc9c9c72985d618f57226967c06142a5ae0b71e4b1a9b412ceb743dedb65605551291ede4823039f01b7eb1c0442c036bf11a72554931508331db6a64b175f2f11b64f59efe13ca9c9026832f7b30f65b498867d18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1678967300e345d217736db87d6b8ab04b0787a7a83efcbfe2be760fc4b93820359370a12bf6cf6ea420eda4568fbbb0a47223fd38f9bd0a83ea06a00d2a1eeeb4ec5cdda7256f0e26c0ec673a09ae93afe12583fdfbbf927ca762d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5c7a8adf5f9487cc29607e5d1904373d2cf3c1f673e2f07e6ca23545964cd045a9ec547de7ec439c67d44b693a17e878a6928b4a7d43a56a5ce4ecd157a0111dc7a7afb97f97c0fca50cbc1b57fa2519dda76c966601ed2044a9d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h99d0fca6c6b7100118c24a80f07c7d0f2c6b1e1ec0e0bec7167f441727fdf7640b9b52130c1a82d24ce72fed8f37cfd84fb2264539349b6beee58e8f0ea8225360add46bd631565063cb379a5f84466fe03b9e0117890516004cf3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a299944d15876b4b16059978cc729aba7f4ee3ac9ff28d7340520dce77fc45b9ee9de5a89260510b41c9416070e3de1e1e6a2dbdef14153bae4f8d80d42b2e0493fdaef5030f2f8f0b032afeb90c495f46b05d4306318a6b01cbb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h619558a7c529b37f3703e0348eaadc506cf0f1c7878fc46fa5de6554dff9e5c48179a58f1840f7d5905d840069764f973a0cd8d67d7175d2660234d3581e2359aee50f007aa5ea413b7c24d2f15e3c0ac9cbe658930a6bb3d2bec8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h163f5721161ddc3122bfb8ef57f9a06309a5d7988d5d8a03c2569fe3df1400c7daf349201b50729172544d041d6fe1c201dd001897ff3ce0ca34c64fdc624e6ff499986913fb877c0bb04a368fa607df9a9d76d26c9533653362dc4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10798451482e80327ef49d3ea4cfdb2b399c92fa33f8dd40938cb37c7e186feae157afe89e4b7eeba883b992225489af4f6a887252fa9cee39d889e71538132d02500c38d8868d1da6c37d3fca99aaa78aa80208a830c3f9dab0f38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12a72b023bcfa44dc67bfea5d76f4773241cd90238ea6604e02cb504069b07e484866064a884fba6913dd36f484c584176f8402a124f407d35a4ccd986f8e64f992c4e6376d400d622e05c77e3ae9ab1ed332670a6346bf3627338d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10467feb0167c4c1ce99dcd28e44c031e79566d0d690388d51b1a2cb735970a7c6234291a36afb272d62170807245ed91cab3ef40e78de226a3e3ac1c6b5eb8ca0635a23af42d5f9194cc10a2bcdf175e0af51b579f7aa132a0a132;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c3265b9ed429d69def34245cb0a712f521d4ebaa8626ca2298061e08ce3c95cd9626e337c2070bb3c1e9e1d4a5de5b4c719fd1a9d88cdcbe27f303306e7c8e1f756ef63375863d16b337e10078cc929c4bf77445107cbf90f3bc3c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c89be3a13c42b2bb46e8b0eeb900974b6ad4574173563735f8d24cff6d9c83fec4a62efaf0490f8a024a39df345000eec3da580bfbec6635f2eead2aa7a1ec93574e5ea5671c5707eeb025bd73ecbb33fdc3be04a07414df57972;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d2fbb1e4bb93f270e80a100e886dd2b4c90a00b85cf8a4fea79cd87b18ae8ac150efda9cb6f086b07a8c1bd22e13ac671e2ef363e74cbb97d300be5297ee6bdf4b429e1a79fd137de0dae97ed765ec29df627c2f88c00db58f664e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1313e6d22d8510fbcaf95af8d17454b6ac152fe8134e532479e3b233067f494a2f65e709da89057f5d3d3e203b425a70dab790af301c3921a34b7054f43d498ab71d0e07a0fe2c6d8b927b3799e938b10dc97bcb881c5af2ba9dfb3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15bdcb316f53544295f92851b909a548657642258a84cf863f7233ad668f1374904a5b8b2824f57dd93d9c8655c67c3db589b7b9ac01b74c78e1974bb075238b19db5bb06b99f2668b7bb5a6e6aca2b132548d702882df34f0e8021;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c0a1cac66e540e55398d761a2173757f7b58ff91cee6dcadc3d0b81bd44d62b69df5cbe66f9c231716861e806a430fdcc5d1280cf37f79e46582ce1d63295323dff1b660f08a00ab6c2e3bd7321b5d6bf2d2ebfa9ba0ffa0a1e1fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h240007d18ce6a3fc17c84af514062f0bc41caba6906ac3ec7a46432c673b1d2c69fc9000f9fcfd442c42e9fcddc1f7b30b6fcb1b153823c3ab68991adbc4d7279cb960a428a93ec136694a70a4544fcb4c13ac5befe22cb4b2d5f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16f3f6a69c017a4a2cf9dec5a7ee784308bf27c05476e9101ae7cae01941e5c48965281370be47ac403b1a8b604b669c4c99cbca6a6b0f070bd9ee9e0e27d89eb651aca20fccce12883591ecd222a5bf51256cae5b1d55dce41a6aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19e8556eca6413def32b2cb17f3d61f58cde53c790f4d04454e862e5eaac672b2b518fd5d56344dc983041157a409b3cb8e9912efc739c47eefd3d89e587f4b0ba47b3b01b3305eb475f634f68bd5885d90bbb0a1f489601e70f45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h582b792c19ff6cfc0937b51e60d43494170e0f4a3aa233183f77a5fde5a8cedb916f89d063de1888ed8f9a7722e0de330eb1bbbd32ed38954f9a89fb659a460355985e6cb31b3c9e0c26272611f04208cbd93a5a476ff90cbb6734;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2427f4ccc2d10c850c79e8de64d99a8c90a945768569c5aa866fb4ead7e81a4ea00272be17d1109ca5ef57aeec16b8e0e5c905c24960e2c25a15eae31cf3decaf0e8b8fe6ee11eb091c295c02e843e3ba8d98283a0a7e9f5ef0d55;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7c799718e2873718cdfa1670d318e66da7df680ace8393402009ed29590246668ad924f1ee638b360322e5a058f84d4a155184dea61c5ec1cb79c2b39533768284d547173c6c3686d90259a3be78cb12e02e4e0d1289ba94817806;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6f481f91a77e5bdf3a38045d33cd93ff7a3b416f4e448c710917455382ea13c2521fdeec0d8a5443bd50f87bd8b7ad7a481bfb6920bfa4e046bee7e1e2c29529fef35924ea6890ed59ff1b8ce668f4ea10825a77619b55637c1467;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb414be85c80794e07772de8e1074902c65636c9d22a7529471701c7858ed1091341e7389a1699bcdbd579a5c727956259b2bac24a6d632256c08a8bddf628ccfb08634add5af6d31ae63a94a49c1e87495a959e6399ac3635dcb10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1babef24aeb9ee08302c4051076cf4991031ec1181a8d52746545b906fe31a1e8727c38fb4e4d9506bd1e40123dac10376c82e874bb0628a4007603ecbcb4d3e4bdfb1b3786c8d8273102148ee014247fae76da9cb1d64e7f5d8f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h141589279598794803684fc21b8eccb860cbaffe39835ac7e3965bb87bef931f6c83d6b945ada331de8f1edb6da512e8f59aa4b8793c9b176ee8a7db265229e44b21ae138d8acb0b6889460e3c0c2565ad3b34356d52930a215061;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8b2b78ec27e4683bd43a8bd790f4428bb8eb8ef50f8672f1c16c79db97a5394d41e1fc0e353ae8c0e435b097144fca66ce29e361b83853f483093fcdd2ea71b016015a2afabdcd1957e9b6f29159d465b50be8560ec7801e1124ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha59d0aab04441ebc2e159bb1e72be30aedef83e2d81ae619f0090f537d7a43801b65235886e64e60bb8aa9970ec093f394d7f78ffd0c18c2f151b424ca0688d0ae3ee1f1b52d2e1f750498c1942e6d6c241574bb56c1ed86f0181a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf6016f16686cb26e8893547ce007d646bf87be9f889677cfbdee8c42c67815cb04b3c8e71ffdc3d62dd4ee929eb146a9b25ff967172ea7980136b56d0ef16e8611fc5a5d70607bc1b8bc454dac88a5c622b41a159819926db4303c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1547cb94199dc6fe9ae295b96ca76518db384ec8cd416183bf8e870aaedc8f25d2e86ae7384eab0826751d4be160f7f795ab5a98637a130d977cbc8525c3d0c7622ba4e4d22b3af84afccf3b1e7fbe7290f05891a4fbc749a60502f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h79455b5e0968c6de5c159c0831815d833e3c9163e62fa5763dbc0463383610beefdab5b17581632b3c393e039afff9cdc8c319f0a5f7c6894fb92b0ce5a78d4ea17bd4e0eb5e86025b5f408c892cf92f31928ddeeddedb9bf5cff8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h99def18a141d7dcd192a9e59ea92a9448ea726e5c82c98edb0aa16507b17b7129c19b043e0dc663908a591490799d3001d7445cde90f69ff54aee139f44092021e5da87b2090d6231f86c3d05f1fd643385f126fdd59325ec58590;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12deb7f27949cd1e08455a9f5167b7c6c9b8865e95491ffe595fd9073b412209086a8a92da5e3fef06636b3b5e9949ffe8fde0d687740a93c702e34a5810b1a408bc35f5f466f2d3f6cb1b16def1cfdf3a3189b238efc2c81af9182;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he0d476ef1076214aa15dff051912d1ae5d2a4e190e477de82755ae0dd6f2a4cb216c684fcca81612a5e5afe637031fefa8792c1b0e3b0cc59e17e18ce76e7d85a075167b99626f2c03cf9367394de6bd8379fdda576da6676d7970;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14e87552d1719dbd1e0b7967652c115b20134715ed0e60cb459ec6eda00f472c79134047378d158c6a40985775646cdc13c4e24c452154d3fe6661906c853d1e446a04e432eb85e0565da430b88c898921f17b58b50deac2ef7e6f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1721760e92f7063177351d27373ac35b574e78d36648659afebd46b4fd94aaa785e177f33689a91c6c321ddac60b0952425ad354950ccb814b91a95e1079d7e6ad9e5b91f03932385880642dcb4f62388396f7de4db6dba0c486411;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14330151e919fe7a74f78c2fb696bae423cb0f1dcdc7ad10f95e2cda04a5f70754c2b43a5327fdad5fbcc8022cf97a88b3cdd79a36cd627eb340a35289640309a466909b3999ae0b871576b883d5bac1c8bf0503be474d22a7541e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17d8a18909bbe63e90dd79929ac3836e233215ba9262a3cc4ade63a3418a67a92a09239bb549849d4e9d6a27b072f9eb8a3233dee6091a92e5424d8193ac7031524aa88381aa8feccde274bc796134956eeb9cebce36300fbdb359f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11c1e5006f43edd6042ce26e42afa7d794210688b13cc8cbd9de1ef9a7c9b463aac3a7ed901caf86ed96dc2b3bf04bf4cb995414a4932ceec2c423f6f77ee9a58740cfee09b6cf2e63fb1355034cc32419df95978cb2f626b7237a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2d9070b3cd31ce9ae4d3a3c155b35ce1f82e6799bf77a6cd5d18289b684ee5fb5e9e5c039b0d44daf2cf4122550b9f12fae492024e20110eff16a6ba74d30490350c0c599b6aa4b506b1de49842e36c2c9e165ae818f8864e70433;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d40174b49300061535eaf8f824dde06985867af113a6cdf64edbe6c630e9b78d4e69adbdf640e03ac3e79fc56315d842e57c79958cc2b74e90bca6604a3205cae632645e8e6049efbf041e604af7b6a5260d80dca2594462c55078;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1586dd39b9ae814ce7f51203721f9ca616cd9d197515547968b028734942bc12f047ff55d0cc4d72faa1a29fc3e0ab059fb2e148cfbc4a5fc5b9998d30aa587bf330f24deed68dda02a9c1daccf2208b9f161e058d99b657bd09dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11adf9020143f48dde8e7590d05704a3bbbb4b0320004c7330407eb5f822a0a01c475419c45eb66459df464febf41ecf844224742208d4cc320ccda233fbb3e322562760533c8ec86c47c6dc65de8ce30c9836a40c7ba1194e12944;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h211816d2b33b55aab94fbee7961cd6aeb8d2fcdf55bf29c38b1b1ae1e8407f6a74d2dd6f1dcd0354b60edb3fa1ab07df1de6720c280b76e8beaaf14e72920aaff012eee213ceef090f597d9ad30d47a24ba6a42ffdc1ea15d6e0c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f8c67d2764c60738d41170d4b6354759f1b992550d0e7cf546815414872d11125e126de50c10e9abed873b6762ccab259b508197460dcf8ae4b5014ca5112355c516cbb8d48c1bf53e4212bba4633114d1de22c428cf79c305a058;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b097c8ea5537c1aa30f4f25ec4446a6c7b247dd59718769211abfb545c0ffd546094c1e7df1b1dbd09daa219f2369d099c532f4bcb4e901b8bc0195a4254802993f7d18b506aaef23f5bf51967059ecf879b2d23998153cb233d41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h179552e6333781bf0ead35a751f705a757852a40dba3710d44ba7a9378181d87a0586ae383ddcc4810a404268c877a7d3b782c51ebaae5e970ad1e262a2b137659fbb09e6c9a2e4d5013fbc1fd1eb4674418200d4256f11e43eb9c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he8a45ac1e81fc07fea78f721a62eac7ab4aa55d22c05e456dc033c60fc88be8c485c7a42aad3adca29c333af13b8f9437b0ce4bb3c267a18864a07d8834489cf9490721739cdaa709d2a25f7a1a587f62797238e8df92f0fa3565e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfba42a9536dd39a372fa08cee1e82e35c5b056b0dee16d713d91e80c50041051a1cb59cd6ccf61e7bca121e0d01bb440ffee1e71ac0a1e0cb35bdba935d8d355d9fd804a2dbbed9ce0b1cf01aaac0781c01711b6f911173b69d80f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a1edb6de691e5ac580921798f5e277640dadd13fedf50dac635f13eb364853ca28f5e3eb3535f6e21fcc4851cd38b0e3c83118757b9ef5ed07bb4d04ff257fe17c856dd1485f9a0083dbdae9bb710bf3b4184b7d6e5c73fe4cc0eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d7443d4b362daed55cf435e929d5e1e964ca9af0df9a48ba4f6de4cca2eeb89a0b56e23e74a1d7ccf10727f67fa0ccb0ba7737033a9685d8ded36f9d8e22e140fc5ff639b07cf109e0f85ebae67c0c504462ce894bf604e8d8074a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h30ba4e8f2ac47ff392761cee55af82aceb8d11230f9f3673d133272d997682c1cbeb12af7bfe57a75b061323eb386c76caada166c9a583d2210ddd2214d521f08abd31efc100bc2866dd0a125b6510359bfde3268b42669d88c041;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2e001665ccd58b97b0ec181b1cb9d6fe0f70b71bce604a42187015a1469285ec0316406e6db7fc901398aeee1715f656661500f6f5ccae2c57a45c378ece6349a0f88d80b301f5217d04c66fc0d1ecb14e2a286701b7ba5865320;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1d120009992373652c312c2ed58bd9e8ff571faac1103a76df18685742483b9d708da0db1eb68454084af87b36c5c801c874a548bfd63ae4cf9e9f33e7f73d11b9b02fef332b762fc45c91ba59191ba56e3e9af929c6a46b0f2b2da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5f9cd8d39647bc7f0ea65318d66436b3848b522b69d12743ddb61eb3cf6f4d95bf3aa8ca17e5dc6115b3e51d27c6dfa9b6ed655f17379aeaf1d5f4a2ec84441a1e37e643479b3dfc9767a7847129358858d96e28ec1798948f39a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9d3ff4a2f440f2e590c143c7f444c14960454ba1a9a7f8c9a4a67a47bb98433f5954703ce2e84aef9142c60edeaf0a9004223082599985b07ef7d8a753f30a078929df9076c97b85dcafb1c8ad22f076d98b2748ec3a16717501f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9fec950c156ddd157b755b810e9078982bdfe3235b1a73d6f340ab633f5f1376fa4c790a065082ca462712c10fb07a1b86f9f3e240386a5be4bcfa0df74929b84336ea0c02d012aa54f262fb49fa4930fdb65bf0d98882bde365e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6f9d85ee16e57f0f2cd6220a5d167abb90a99ee6eb45f5f20ba36ca26d89b02cacc24597fd5d3460fa00d2a5632eeb32a6ac98c0299369943d104b26263bef93afab0da9bd030a573309c3d6b6e8013599cc3e57d69afde857e25c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h362779e5b622157a70c7b96d12073a236ff20f9b19f1fc16d811b84be1e413e1e155926c0df21e97620254883ee2c5ef9dcbde5bd568c610ff97bfdb7ce3280ecc48ee18c48cdd903559746f09a1dae4d00efe0160471054d73de2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h186a9682a00703cf6d0d43930c2a9001f94df151ec11501cee7abae836d84f1476546f1bd36c7b9567820cd256d54fc667f656c503b14346c852eb4da37dbe7f536e6a5f5fddc5bba4bd49409657bb5b49d49e2e598cca2f0649a24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h196aa9d5449245228471a0c60dc190983103845c303cf1f4099ed214adbaee36cdeef0e46622679b138df6b4a7ec85bf0b13de9e0a4a359a0bfd5af10f06cb36a076b0b41f830fb566020cb6f2ae31475fbcc5de235abd81d2da2ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb5c9f54ace69db48999a6a326161a6d2680817b115cfd9b7f7bcef84b19e27aa8f5a172f0e960b213e1caf8a4fd4e7172ca060f917b2673ac05aacb01bfc9148ebfc44698bc363c039902134fd53da6015684fa81ee18bc535eb20;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177f30e2a53fef1087d123b07e029096989c14381d155a1cb16a5f12f72259936362f2488a88b89595072252c28e7fc0d7f2d52819d0641623ac26543747774693f089bc7e9e4f0a87e012e10aafa59891a7d77b534adf0d9328a1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf58281fcaf69916965708237e5fcc6f49020f73ecb1da9c102911da32ad07d96ed9f566d0b3967c3f4ed1ffc61d1679ff2b6ddd1fb2b40874dd76073457046b1f6805763f1fcfb7472d6782f4150d4a586ce1c355cbdef654d948a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12c7d97de390c3772715ef2fc0ec763b355a9d963ed9bb65236b17f6b754c2617dc636389d57f44a24bb04da2d9aa4079dbb7f456b62d8aa625b7aa8c9fb98b6da9eb219bb5b7604568a7c4553b41b8cdabb382944695d0d2af2874;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19d9f13fb97c01ff5adb25cb6939579f48415096b1e236ee69f8a9f5084e5c0af2203b390f1d5e2e4ad847863fa0e3bc590830ee0d834026ad613e49ef44b9e7af1560fdfd9eda96dbe478c15ad4bcd34dd47709eb89c237ae10a4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h99d6f530dcaca1844941b60ef9b8d86c1985ff20d6700d5659ec3763b5a028e1c6a295b913d43977d4ea4922de4000493e17796b738f2cdb6644ff42666a9c5a1e4503a1f824be09a8ad0da2ac5f4909cf3ec1724ec0fe80a8640b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16c1051ae0b0a86d5ae569d696b3519cb949cbad346161a619e2dd2cf8e8e29753f44f0c3f8caf71464fb6d23d62e68239b0113891d0654384430880491aef383147ead8f7d7a3ff3e76c30c710e15c1f2d10c0d70e4d9ddb4d7b9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19802d3f21752897319a0dd71866ee61e732d056e86673efedeb8971a66d1e79a74a4f81b623393f91cb1ce9335727091f8ee1be20b90a5ba345b6ae4ae3e0d0b6e4d13bec40fbcd0636af757a502678160ac5be9e97f37a36b9934;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d963c895b0b18873f1d06f5108a54bf68f1fb1a164f0f7dc8d9cafae58cbf06ec92b08863d780a162965f5aeb30fb5ec37689d78330543ac6b7475c3461254668dc5237157acdff73d5954d53fa841bdf4814912407f624e4bd24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2919b5a11434519fcaa94585ff76a57e37a363a2e6339835e8dd1229726d60181bc6e023ae8acd85f1099ea0ef9bc31468e64e9251a7ddde575844fbfd1a84d29e418055ff1a23f314bbd44aff647d3b9faf715ee6856978651b7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2e9b34a8e3638c9309e9567f2541e1601e08819cd282368773fb39894db147129e31244f542639f0bebe1b786836f53af0336c7d11bde2c61b3f946db4455adbaf32aba1949fdd1a69ca5c266aec6b0a70fc1a824a631f57e86eb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc711fb5f13bd885a671d7666b4de1f414035949d73a96df0a5cf23d465fab0297534c0c1f7c58d4f1e66b840150637d89fccb2707acf7e36d93af9097cc262ae179f630c98e418ac8d90339bb590b7c4080e4ae1614eefb4ddb7c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2eed672691f6402a3e1aff1e386099519b641bc1c6ec8fe1ad28db6d3a6370255385a774a867d40691eaf4e990382e668537fd37e7c2184016bb55d0488d5498a41a4242f9c9f2c08a9e56cdd4dd08c2e9b8b74fc27b6c0802a54c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf2e533c1f99e282f5b6cd12cc39606d1e63529cc9f334f072aa0089d5f1712a18404f98c35614ca52d8312c3c759d530ea031fac7a7d5ca2cf31083855dc3a63cc0d76593fe160baa7d245f2130758728f55645b7a96570f8d1fdb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbbb0e7b768a3b975593557d23f292014a33104abd2abf2d956cd66356d0fffb7b97785a4de75ad4b599975b609ed13e1088756e7a7bc3cf72332480658aac4077e36dad2e49695d59db32f865b4dc1f3d98af9b39232340e95cd45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd945c7e0b45ded1040af30af21dc23b1c9f409da5f32d9643483f4c0ffb603ead7a615361c90f7b01e5268608fe67e3075f2f46bce95c9e631d142613d3fd8cf493432b0e45e08c35e835dd1277c05ffda16d6f97e8ea2d27e4378;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3d809afe7a0bd677f0976c68f2f179b16f170993c2922ab8e62b08350ba6f388c259ac5790be320355d4eb0a8d587b170adb13b564fd13e27b5aba3007891f828f56eb53380d12b0e3309052b810134e242a66ed8f796501a8616e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4bcd444e6db41f15b7219315c2bc07725f44850e2b95e6ac9f5d8a19b9e7c0e18a9fd5e55b21137e37e60c5dab8d5b177bdbc23a3c9b47638ddc514199ee3c8f9c295626b951c5bddc9ec1fb599a266a34f2877075b00222cb879;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5a36589cd67954ce7f9bc6584eb9d3db70263b271d4f1965f9f95d7893519181dd32553a398d03d6be593ae7855b1cb0c2dc55c3a09d596d2635a615552315293f23277aa4a62507340a0ce485b15b6e6fcff477fba866ac04fc1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7f763dac99d63c53abb6da2fbc51f8984bf83634e78f9d4ab26eb246c68975cefd8678f180febf56e87b27d5dd6ac8b599c5ef8731ae667d5722bb274bcc5be7783ac6e2b42c4814085b9ca3e3ec220d77317ab2e572c5f3fcb38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf4d7cc294d49661d52121768e12ae158783af27fba98369573618a26b752ddd605be68d9af5b1fd3a02a7a2c4b3332bc6264c28ab0895841e57abdf793d023c1ec1912458f4a450bfd7a19e8e3d1f5e1f9c95d20932746ee543cf8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8d9a8b8ef21ca8ae6f47520d0ccea1d0fb2986962b7c6a5ef5138e6170d83632f1ae2e676fb89c83bc2c78b7661343119057047d7cd0095627536bf6fe13774a6dc564972b0799079ea1bd917e7073573c574d1133a7a4bb8f91df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h62cc1f8b1ff70c59f0801b6649d4319a138a6bc1335cc2ca47b90a9e8cd132096f41b31b0338aaf39b36272736e321fca0eca7db2b92fd94b2e9b386307cb97f2bd08478a84513e9009ce072471ad627ea94198815b90473e9b105;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b5e6b9b05cec4c43a8873c0b7b06deb70e19e2888df57d0fede8e64bcf45bcea18c8ed8c6086fb11d0d05f4e1bf69cdf8f6b765b39a5c78b49bd690ade3b0b9f9207ed0a936da9bfc04de9432b72f42fa63f33b38e8c1f138a55b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h76ceb80aa8fc5672df41a178897d9da9c990bd1cb972dd4e0e99bd9a9d236d8a74227353c521455a41175b7dbfd91c159b304a24d3b3af18f8a36ca676561b5f7e05268c0b27148c2c523224e361ebfb5ce1f2f97762d88f360534;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a09ba41835190a66f278ac65fcc402a6cc66786c2de9cca91f49b0d3374651653759f0d2bc382f146a50785171e9d3b3c90af02351a6fe457a7fc867d0fb6db08fe9a5a2b2ace34ae562e07799dd49834c1d4fe3b239fbadf00d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb623ec4f00c002d849f1aadce96e096b5ed3552756e5e24b30c95429a3f2fab38372f4b1c3ed956ff3dced4276552cf558605913b62e1ae90f2eb89c414f1f51b7e89264d2412902e3d8f0ca0958603741a57fe783a06bc8248b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa648df6bc7cd2a5d4a171f0448690bac6e9f1551f1b5363871b2191c7cf6cf07ebd30769b931eaf9f97a3140485f5aef4832e9a53ee0d67dfda27ab1c7445c7cfa3428e722937f1fc8d280749b8cce1d6d4293454a10f14ba445b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1845f777df75ca7e853893822301136454107d03f3c8404f98fe3e54374f36f55f749bd37849ee217f76e372b30304dbf00a0606ef9f30b0beaf05c274481d72531522132119e45febe21e2af61725f9b872e103a2745dc458542ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h83af5adbbb3111252de58b32bc0f492a0d2e74965adf3d189e1416fa0ca562f6d94a9695a1646cc185342974784b31b5a2937fd4d2779185760887aec5054c4bc8f5092379278f2cfc420c40f781aad1b55c4eab5b68e0b6dd0d64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1674fb8e469a2245e23954a39a1c9ea3bacd671314653ac3a165f76d4c5c116c0ce8118ed869a3e2d7e82db788bd5b6895b19c3502ff65ac13a897ece3088392e83b529368b1aac7a34e0485f9f492a115d53aaa0980e45f5051c34;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h43707383a861436f687e6eafb5e515590dfb472d8dae9e0a03b43f919369860b63e9a6c8688e162826527ba40e47cd84db6bf98d5f8bb89012da490d70b4353f32231351b87b500dc1eded179411d107b3220d13fb54c235165503;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h29cc74ecd4883b3c23a6818fff8244661d0bb820041a894b40d5a29b6e53f3998e27300a730e735a51c4f5ee76e3b169e39b0e9889891bccbf490880e8879d2f969a6e2fd9004b7e5acbcb3d349cd87bd0cf3cfbfd8e01fa5318de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b9858cc5fb9f1764ff993904c48fc676079a2bf47b6238903641a905564f36a8ce465357e430b58c32c668dec4c03bc64abeccf9934564b21c5d7c536d3d1050326047f7a2ea5974f361297597640fb146e0563059605b3547198;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1dce9335185ea4cd44b77aab5a942c3a28c32905a79eb54c1b62e1b48789878a9b635f9ea0e270609c4de511d319cf59f97307cdd69fd04837a8824c1094a0b00284c42a1c823a1360fa00708bb1167ed38a77ff36c969d25610d1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1665c029e52e8aff9d8d16bc662ad96b296ea5e412ab0dd878bc610dfc93e281b1d22dd3077fc9061880ed6720772d767ab98b0aa4c6e5c576906fb2cdf3aa28a98f645cf0401419ad08fc895cfb29df87969d9fd3c0d6abec381a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9eae13e0f570b19045cbc5d967d5d9575253127d14e29f0244c4692347c247a04b137f743542508b2299d2ca451a0bcc249a13f4b5376cfae8cac02fa2bfedb28285f36f32a9c133d6cb3db9d36f8d6038df72a51e44eb4f5b9b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f7542a1525d68db91095e0b1536955d6740a67f99ea10c15070b1940702f71d2fab9086127e13dfcaa47d0582556077a4bc2ec0cd86b61b94c4a383c19c0bb7cf92bf5f9802453e6d7e46102bfea2dc54fefe06f4b9659b45a3f9d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4e9b12516935345cf9329f3d66e78ce657fcb91b29c883c4bfba490801c296f168aa6679486ef591c680c3779cce4ced491f6861cffc2831ed80518935fb3e3407f97c7ff12ffa04de45c2cd5ba36b0c1b7c0106f24589289dd106;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h953e8945041a52c619a696c50fa25b419e6c5d38f260dc11e16bf8a93cf485f4bb747ad31d64153dc1bdcb1f0363bb75e16734a5cd136af69fefb6ba38d85de758c5387fcd52f4253e5e83e716a3efd32fa058a381a0d4f89558bd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f8d4a49273f1feea567884bcdcebb7f598ea59651a3cbcc306e4449b76a855275fe4657703a0fdecf321cb3cc0728a6e52d6f55ff726addde1da9d66f57aedfd77362fd3c8afe70959e182a13dd85d48a306cb4674bd1eccb4fc93;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha198e75be3f0abad8740c8f4b136c29a10f3e20915d3991ccd52026bd90bb013c9d3c7529c864b4cfdaad6cab85c1b24b7fcf858990fc2ab8950faf5e7026c24fb0152ffcf764fbd991ac874010528ec3dc9d01b4c192e044f41cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8a860910e76caa52bf5849b3ec624880d1082d67f8e5f844666084e51a108f28fda62d44db0ed8fd614e898dda7eb300eddbb48e151e5ae3035c06374088d48fcddb140aff15ce574a2b7ffdc95f44279f1068096e337adfba7bc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1657076d73dbbb03d94891524397f87e603ee4bc1fa77dad75014c5d350c8b0a3577f24c4098904beae58d2126752356c7f22390b736ceec23fbef07fcaa043098760a3ab6d789fad084d733cbcc150b248e3b5806fc4af3b47180e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16adb77bd557c1d10bf007c7765522b0ba5f5187fdae426d82076e29e40bdba6b733165115b89d7109f7016b604760ae3ea063b664e9ed5c47d345201558b393d301919bd22a478fc442fd242f094968536f9a16cccba714f0003e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h142bd0495d8c0a10578bf76dde26060f64fdcf0dba10625de8b059a0e4ce01e9df298eca761234e5bb7805556c1e738eb89fee3eb6347393a0862fc042ab3d8d54d50241900d8db38d8e0019efb3eaf29b311875bf8a50143f2e242;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1900022bfa6610b62dc116b65fa643be9dba05259b87df8dc1d1e3f33ee14c66af88a852effbb9f8b6ed1f825d6a2258d8f1b5f0737ba011e9bae3cd59598701061334d186beacff3b01aa57ae07da65be1f35ed608e950d7a108b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h111f33b2f6e73d714528c96459c55627a0787ed8185bb32ca8c8ce601b5c8820d0e27d0a1643f4a41f9997bf02ad682ee44aab8115e91700051b54abf035fe984faf87a02759ca2a37a95f5eda5648ef2feaaae46f04252a75213a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cc9e25710307494f3a79307aa91d3165258be28f0ffb2f0e134daf54d42575fffb572f48f6c15c94df0d31ae07f84f6abfc5e991cdb8a135bce7ead6bbf800bff1377a7b449bdd0d824c21118ec630118d14df84ef267699cf6945;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f130cece81ab8cc0553c8101d2cef66973f6c1f5756adc5534addb16d50a93044eadb4e384e02eda0fad02644d15ecf8593bc6247b4748da11ab5207211cc3474b68102532c3e0137e75a00eafe3a5e0d6079e072c9e961edcf175;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e2dd2e64b592b29e18167d26ac09281076d1d24f52dc8b7aa5131fdce90a0c1ac308d7e9c51bf0c7ba31be91eebb34b5391e681bf46c7eb54f53a92b01674c7bb61406782378e6b36558f866938e3b6b46a63673760972ed12e9be;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf6d8967c676f48a457d752fa77768724d8aa33a8e89df582461c4312273a0559e997e32ab8ce622bc59aa54f7e7abb4df7a34de01ddaf92b8ff25e7242b34575a425763260c5d00cbcd00ad725131c3a621d7642513ac4f708ee61;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105146c7f05425cec0f7bf58e6ec14809c1e8ace819a5680fe06883ca8bc404113eaa3bd15bb3d90ca266170526114de63624f4121a3b68604ca197768cddab77cac7d53a6ba5794f9ee258a1342cd8d8ed740bea58ecb45785da67;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1042a6ed177d84cce5a6e526bfae1347aa2cffef8872237d2d469607131140bf44214488ca2baab41aa5498704d76596a180cdce0f333c416741b55677750c7033ea4eaad0153c8f8e7fd7140b766b5475e5eabc6e4baa711aba9cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a9b8a7b75db5f42e943e8b205043dd0ad2ded8ad6d085901b1848b38bce0a0aab21082b915b0dae413f2c1d808e4192e75bf583caee278ab75b5788b02cc3b2c4d687b11024bd19ceb14d29cc97d58008c975701daa6e78d93c17b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb29dd0cae515a824dc062fabb05ac7460b8c5e816924ae4ec3e230edbe47fe98e6b4ed2bf806e89c4b7456abdd37ea40fd98e79cf156db552701102dfaaea0607caddaacd37b9575fddf4e9dce0fcc3860dc48da71056d77ccc576;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc3c42eec3fb3ac6417238b224beb3a7ab4cb80c7a47dcf478b0bf9226a46ef304d360aaaeb89894a1d74ebc48b1dcab2f99f32366ab4aa832652c7e297ae00059f1aa965fad2eea91b185e38484fd286f1bbb63ef79659916039b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h191639af41c903b0e3853aa707ee42d87f412a2b0d8594b2359828ff0e7d9fdc6f9a319d1177a7ef49f1f61c6ccc2b117a73f06fe087ac78606d8ed2d8466782b14cc59ff21d9f8c2c465478f1797458be5be6dcd362f67d4e09b30;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97b2a4877659ef3bda37ec5c5cb484736824d750c7268c3f6328f221bf6676ed5a86a311ed279d5c4ae44c325c0c94c90603d9659534cd05c25e77b9097316e90b9f23ed0cf31b3b2f86e479acc9bc7a92c04d0bbccde1599d1cf3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h97ab4e6a5a7b7c2b2f11acb8f5fcf339fc0909a3e2cf1f4c085082f36ff806d308ed6740d64700d55910494c6a06a3c0b132540583e85b66974dc785e5443a4929fc9aac92d98a80f3c68ef971d7748fca02790dfdf655e664455f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h151372dcc791708a87a0ec2abae1a33b29230ed182556014830a11f6827e7cfdff1b042e76ee8c9f23ef3893946cd94c991922eb6169c77131c4e2366a5dec9fef1213ccbc2b825e0bc11c1318d30e9f4828169b5d53ab6b58c08d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha39589ab28a66e1b07a8fa770b51243a213756b2d2694c05d197f789360d2d9ce84ce1605fa92aede33b8f15478de63e6e67560f01ddc3738109ae03db28c7a80d21c4d23e9dc1692c3f51d0ca7cc798621332890f2dbec32514c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4f74c54fb31c2babfd3347cccbb152a44bbb6fabce2722fb337e39228200ecf21022c41f950b229dd0875e288f6a68ab02b0939397d3416060e2dbdce11df59640dad0a789c887840d96f8c280c20f58ad46ce262b613a18b05e2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19a094b64a646623e78b5bf090988b557125a913b01ce18f06973e9cf3415c2c706ea5048720526c2c3343e68a2a32f5307aacc043f28cc7580ef89e96762e9cdc2f85f74af9e98504260e8f63c05f3be8588fc5aa42d1a31941dc7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdfffe459a1b14b9df417ef2d77eca396828c666b6d60486b74cb35110ed15df67ab44e1c89a90ebc5afc5f5e43b9ca190ada0ce591abc48be3d06902c9d618058a85304a7af304fbaf70be13e530548985317ef7c0394da9ab5e7a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa211d55718f35c137aea3565e950c192c59f75db98651230178b4f996fb64c883a99877440b675267f6f2b9a1856359f12d43e253179f8bf74f2391331842d84ae30d817420bc2e95b67beaec24348403e10e039f05bc15a70724;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9b67bc797cae4b1e4e87cd07d78159300953e7ede64e1fc9c69a82eee61e4fd9708b7b4af4487a31fc0b3c83c6c6c0f94aaa5f73713771d1355a38c7cc749c74ee6ff19a677b3e04145e84ce98c3ee74eab78778315be16791390d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1198ef35113c97f2f5458686112297e001343b5df25cc05480129d5deb47cd130cec27d326017154eb1f3e9436753cb78a27e7b6cd806a1f7f2f04fe0fb457523c346fcea40ff123b7a0c8eb399bd21dbb4d4b50025f7475181dd0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a28a3bab063c599ef45ec24b126760c7d1fa7f180f93cfa2e3b32938a9e71aa0dbc37a256957fe07df488496ba967d81d38e365d7245fb3b8ac2e13cb664d10defbb465fb6669c84c2503bf7915bdd435d48d5871a99b911695ae1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h51a51fd78af1f039e6cee21f579172808892927ad0b39d4c4fabbd9f939e107f5122b81ed9648a8d868ee3bb5f5302798f92141bfc24fc09e7c56865eb556569ee921c997e41ec810bec43f96e5e97b0f39e51414ad5f05149ed43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdcb063701660a2dfc2adac20edb8b2688612daa85c544f501d46999b201ee0b529abe9b23ea9e897e6733f12099243446e816b81a85d443fdff552a4ae8710b8a2e4d68d028285ad81a22bd00763c21ea41416a3e28e13deb3f9fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e1ad0bb569be55706c410553d16dee36ad3b56b356e67a7feb1a242db583c86028963f89966f99ce1a79f9f85815c1d10c95ec18c542cbe573eb018477a156bbd9cc58aa9fb36652e877f7d1b9fcccf34926720efad997eeeddaab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haf11e66b35590e7352b6020ac2e650ccba05c0d9cdd329ecc304b4e94eda83582937cecc624ea8a6969bbde0fe0785235754e5b5555fbe7519d0f621c8b9aca1a79588013120f4407cdb815e8f1a575da267e160fcdf3fd08880a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2059265f51698b87ce7aa2af1c8d1cccc2a7118d7951125b1e811a1f42afacf9d1eb48dda1571341248094022acb762e0be6d5a57cbea664776f5f7329f35354e3d3a9bae4e8e0fa1a40fc2f1749c039027b4bf5397c4104681cba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16848aef9a51c3e6ee67b1dc7f2305c20585443371a05710039d342affffe4759aacc53e4990996e9abfa19c22640f3d316e7e4421b393878e66ec314f9372d0477e95a04cec80d21ad2001954a4ed4f0c6893ed85587310f41a468;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c23956372c579a3c261f778867e80291312c1c4272f31a311018cdcb434c859884fb1fec87692bf02df01db4390983b7e8a879a3330caec2408229b5b0534081a824c00850f72df3d8d0564c50a4de88eb34c7090231100df9d661;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h53cc8ce3b8927cd1230e6441bf5849ff8aea6e4c609d61646d3993f108567b080edd38860eb4e3e3698e39d552d98c273ee678b59bcedde6531a1855806f16d353684b793baff62b967cf95fae3a95ab68b3b3116881edad10513e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc4c83ae84e3e25e5876403ab34f3ffd741750c197a69eea328d21b5dd0e001bcdab832f8abdd50123c48a30c416edb7035509cfa34a5d1de195879d453c2b1af87710e83102fb0bbc2fc6bc37a14865ba9b21121e1ce539c20b0cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e4ce0508ad1e7088b295d12a03092654ae7500777f21cc59c34af9636af60c4bb78a7a66419b2257e54a1f01456d2de51a9ea5a385c00ef002680bcadd911554961cc9222d099b2a297f3a54ffb51d496ec64ccddca1a1160ba3f9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c8febc32cb8fb86c9278821022f5221596954d8f8fc6810038a18e21ae9ebe615a2a5b5186b08e75742e6b67b8b741d90e319db0822cfe622ce035954c225ee0372542def38c0156156f3b7df59c37f1212c8d7676a36643a153f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5bad059e6851994e119894c29ad3e22caedb8d8e24eebdd0016d913352d6452f8030a97bd08eee15c3eb125c860536e95a20048730d6d4690e158336a1f2d29f75662f7b36f720242b737cd61ad3d364e184e8875053b3a1733f79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h50ef122e0f1a9d47ee762ea4d3051c83535cd4f60904d159f2ffe80130d43a4aaca8b628bca77a89849f4e9816129dbebc0f67bc33975c8f19ffe4cada85913cc7ddc9d1bd014fc3e78220237cebf15439c8eefe561dbf391f090d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f759ea7d299a46f4c43b5b65c66de67cf3d0ea23ee7c4d2d9f73da49b030e9a5c8b48fb7b921343c84a0436ed486349644e11f7ada34987672da4e990088bee077e6a56ab31b7d874ddc32e7ab7a6413e0c642a891a34fd82d11e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11921adf4010fdf6054c1c444ce3ebf65b8811afa587b274d3eb5887f7aee375f358819aeecf8245c252eb05e790a5881aa7ec6ae730b24ada6d50681cbeac827304cd8378824b58983153d662e1ae72ff9a0b643bb0821ebc6fc5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h184fbeb24f8a2d61bd0825ec83b5b69ee85d08cabbd69abba6e82d6c0b68615f2aa0518b51b9c0eb44f2d87bf8a2da2af1c32fbcbc92acd11d1b5aad2d8da9ca1818d256d471127a18c574823906b7b98d418cf21b5fd9a5ea62de3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h183a2bcf44c2f7997956976b46d3949eb6e4fdbfe9c6571404e034a921d2abe8e75df45df915445ae8442d29febcd4d3a07fa90108478d9d35e877640299ba5d88ea1b11e8349c0b43addeb79513d5cbe6e2c77f337675dcc7868b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17a3068a94897fa435cc2d1b3dc519ebe89b383162647ce54e06b9687c88ff1154a3122f6b3054fe7423efc0a4e89b2b1d39ea8b0a02e81ca076efe36e975ab8fd2c1ea9c5600a3aabd783a11c8eceab5481735ab5e0cbd3e89c5cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haaf3b34029ea42a3fa1e6c074eab819a8d6056a921feea5331d97bb99a9ec435ee7efce29fbf8d51cce8fe30992d2b0b773d92f72b9a2a43af16aee002d2555dcead75ce5a5cdf18104723e7a39489d1d37b47557e69099a9d7103;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcdb5fd5dba89925246bc5cdcbe2b5a1af3371dd570fa36171c22223c8dd7720ff07ae1ccf7da1c61332ba9dfd17d37807330171d04204f325f7cd15b8337a224a3bdb4a69e5ddbd9ddb37d8caa962b02c9664bb1fabfcd8a1c00d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h155b17eb35a7a9fc352473284a5a63f69ae1dbffdb027e7dbee29b3853cf5d6e0c5e64ae7b27ab8faef12ec223f3c18ccee27151e2e82f1e8a41b927258bc44f79fa7e070e2f71cd9d127e9450893ab8cab15fd1da4b250663b4368;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11d38f28c2865e7618e3aa334028297049cc82977fc83b98722daee4d27f5189c359adde12c9aa4aa37e35c78ae4ffc84a1d3768665523873da19e8b429e9f64649cffba80a5ac03e2a757bbc422cb8fa3410338b45fc622a27ac68;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha1485e7cce1f946a2bb5ae7c78304b07cbc27603be678accc0c4ba03c12ca156cd7ca743e37fc3c179cc479d443f7d7eae3967cbb296b1df29f38016dcc63039a2a82b168d1c0640988d205ed56b9e74c9c4007c46c16edb36d80f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h940932fb128c31e29aed93d5dcbe95da456361809c38b92adde6c5dad58063d72fa274e55f1b549189bf175ce7818b73a016597c76fdd2f4816d0291e06523fb25404539639ee97bb9e7ab4117a0c1ff7005fd611bacab6ee27954;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfe2f0e27080bdd0a90f93f917bb54a41f69ac2d7a74354c47194fa611d7908604d7863c3a6f4507b22d6e962208f878c5fd1e256a1cfeb17795bacf62660e565204c5769029b467e63d31a78b2fb247df790a596378f4af2ea4ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19871d623e1eac8a650563ae63d9e2121eb83d0151fa374e07cb901e47a10a37aad224dbf941e6e82b26f1e32fdfd21c40670969f12878b415bf11038832374b087460d1bc0afa7f02d98d03002c97e3fe2d2e727f35ff313c2214d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1148db33c36557cf208b8c6d8e63613a0eea6b9ac0778cd6b2b91fcb2a33c9a4c272d112e371d129a463e61e19e39cdddf5e0e729ffa41a7362970ce7eb2ede63f3b3e41d8a82315dcded464c568cf9707d451e61e34f486ee751c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'had9077dec14f4a3b13c1c93609aba9433f0bc783d27e03e2fb33541551b5800c4fb68f2cd3cf9491b33473b9603774ee267fa5178439914e87b825ef8fc67b2918f9c09f03ade4696358046d98c606e4412714972bb45b411fe572;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1423f76e32c6851ee509a4311d5ca8b22a2abafbe9137af2b8a1c6de0306f521e637a861767af9558f846fdca06cbd776742c53d3bc0de325f0319029e937f1848a7cc035993bfa31f9d7bbae2943380f2fd28deb9af73984019921;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15e967029f02085a4d1f5d80b1baf5d27c00e75a8cae5922b4a988173924f9849416bc6e777cad9502e3b0aac20a5f9dfd2fe91e83345de9c958e3743827d005db6464162992bf12ea078b3f4ceaac542c8d7d0a03997952224a7de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1658ac108e28656d00ffc502d1059791afdd01d1e6bc2adab3fb293d9efd166c22bf26c3fb5ed1f05bef47e7281978864a22c428956d3dfc5cdb1d47855c00c0dc2470fda2273a40d540fd3811fe2be25545352adb286a2b0dd51bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf5be554b0e0ac16a6a467f27f3b9f5726ef4b261bc7c26a92255f3fabb60786d95b0830972c516067e05b9c816d7bff02197c2b0e3ad537af4711425e92d37aa930a96ee1fae92ebcdbdd51fb4dc12b348001d06ea3b3fe36ba5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cbc3b166d981f441860a8231977a15ecd4af842971ab27684e0dee53f079cab605a6bc48a28740d6fe8565cf2f36da985a189e522f7c16e58c80c9ae0b1189b2d27d0c743d5fddd7b4e6d42d9ec850f6007be03df57208db6f7f0a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fb34b13035964e6286ce0cf13da8c5c4f0fd1a0daba203b732964e60cf9cc63f0269ac08de51b27a5ced60fb59112cfa6bb2be630943ccfba693ea6fa3fe3e5716967cf74b21760800cc58bfb7783ddc29b1e9215c3660fc597ce6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15d89f0ecc6e14063a7421574027864e28d1f3eb818011e7045031e25167e570b031975bb015d6d889b3915c34b0cb6928ff6e5f0867d8f409aeb8cb3b1910f757bd209cc5dbc0e10656bcb3ec66d61b70b380c5e0d612ec4a75678;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb147125fdb2c74715332af3ec8d18991740a9596da21f9cc4c50a7f70d15d18f6c44d662402a9028c766416ff9185987beec887b560e7cb8028bd54d44b032936a81ccb593bb78da51150f28e27c712161295f2ccdb6b7ae08a0ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5e27d4d11d2e0fd5b5e99c56ecc2bd73fef89bfbb0dc93bc260e34dde58726a0e193ceb8d19e6d98c66d6bab76403104186df54f72436c895d5305a8f55a565c1888acb56806fd8e73f2e585a3c2ea87f1e53a6ceaba040bff94e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he9f318b1593df58dc305058b4f5d1e9c97fcef148da37c6c834fa997b987e6c95c81c2a1cd2fa4d7ce043023d8d42d3383b20fbccebecbcdb5548677601420ba0cc7cebe41f603eced6b8957b3b20626dcd86885f1f27105315482;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8034e94e0acac0935c17f3b2feabfd7b536241bc539a870d2ddb97505037264cfc7a0becb71f18d4a0ae1f98ec7a0bd5edd93976075b83e6d95c36e8e38d20b9770824429151e7c625b34562ff76fe3ff26c7188d9045cc0f11cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc373276e5c5295c76c6a2cb0955953aacb7a2d66662154db4386564296a859877874944d81468892ef8f4c5e5ff91d371c85b5732b993bbf9ce7788efd6758c74675156de87de7bc636f9b54b8e26b26ddb30c81304a5ea15261b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hce335450ff79f531141aa13e25542561433f3b2e23b1efeb2a10e0dc9ca914dee069f4185d54fa071f488fa9576ad067a0f096bd2259c79ea32b7c7d1a26b358d2ef0fa825238bd2a6f2e2e453a8b89f54d5ee6a760b3e119984cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ec31af693bc595e9437128fb60d8bf08c3d30b9d64e74925925140380391093329b87fa1e3ac15e164cc1a5b11c4270c5091854f7b2bc3d940abb1e31ce4f133a991a1798f97bd1579462430666a39554b8b38ab99d7043b8fd8a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a68c4436ee149d64074644aee768878061f7b6e88965975b137e9220349413a298d05cd88715a8ae6f02c32f5fab6166cb3650e615f7e46924f5736f60355fe8f21d9382b929c5427719f596f67ffa38dcb6d569529102e7b8bef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cc0138b421911b0f812e32ba9c9b3f77d50c17e5c101212e43511336958fe61f0c6ebd1cf9f46248203c061ae9b1ab134653be98d5606307f0220dd04942ffbcadd88d2969d270db0eabc375f90643518d2c0e9a1565ba4acf9992;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h88871cb8126712d9d83396594f7990912ad2d926862b248992872aff25fd4d9359e7f7f888e512a67d749a1aeb181534a90f601ff77e8ad761f9360ff79363ce02b7fdb7ac074af33663b93f822cc3d83b2154133a3caab82338da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h143696418a14d92603d884b648a04f2f39433b09050e86b046fe12365d2eee37324f13ab1334dc896b576e696b8da0f135d8ba27f36898fbdcf111b26bbeda02126b7b76991fef75083ee891ee1a985d83faac51490eaad6946e27d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a2efe36daf40a78024b3ce6016e78673f0bd5483800eb8d39d6f5dd354fd4cec5e7cc89861a20314873004939c2d056113f2c5150bb63dbfd41b3ccfe3d86756d324b34d0c6ae20fadae987286e24e679c5f604a9f7cc5d6b2c630;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdb94c362a0bc61427d503873acaebd17d36d902a0dec410b061383b4f642a01056a8feeb65f0234e09aafc5d2dd1094540b380f49e848e3e54dd3bb006af50395c3c877ffc099f317908c97dc14e61ce7c0d228e611a4319dd28b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4db0de2d87e6c3304d4fb352dceeff4d9cc0db6911c7f2a823c1d528cac3b95a801d31406f10e26f9ac6da89428ea0b8d3b683a6f7c3fb9035e91112d8fdb1f33df658575b750b896a27e695ab9f46989b51fdc6f9c6a564b87632;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h524325ea356f7b6f9ecd07b0b33fde3e5e6871c1892169af720a7921c88432d849574861b7a305bea8857ca06bb61eddb1eca9caf7654300f341f6c73803d8844b094d5e90a8487a7f6411b02811a482725e2864260edf7860e142;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h24cc813766e17861fd47c1571655c3d62c806ac2073a3e800fa25d4160348922f4a4380f90a61a5e09d53df02610d943d1a5531bb7c67af11c34513ac0f33149b22f82a2ee564ff652fcea56d772f0ae146ea32b20371074d467eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdf4e38482830ca4fca78678301169a18e1491ceafe3ab0c747c86212f0247ef2b21ae817de7431d408bfa64bf7a599c2b44741b723cf2bb936f992caf2349e2ff93f99560b15c9bcaf1fbac5b8408ffad3535d2fc455fbc5414849;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ad6165c4f8e49d69435ca6cc2cc2c484fd5d19882af2006f1e548bbbee1b531ab341ec83cdfb8a7c285044fc0d0ae13f5be80e7cd7a9bed6a314f0a9994816654f2ae941be2860f40fb330ef3aa08c99ec9024eeec63b8dcfc48a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1403b13103afd7ed9e15447a3c82833587651bbf0b9ae8a67e02a738a88f27cdd8977bce399a9969f5ffda2e8730571c4c5dafd02837029a76f80cd56a52517c5e55fe6f6ab8e8a8574303c52e456e8c43d5ffc7dfc1547ebb5dc5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h9bb277941d31fe26c4f4f5412a140b92397b9a10797736180a88267c41dd181ce0a4f62ee7c06104e17f037901aeb115b1e71fb4758521189001cf557ea2201d95136664c556a44811b2b788566c6d9c311a6ba3305fee6ee4c394;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7266aa6a94cca0e23e3b2b7e2f167756e39226af1ce63bec3fdde71e164b1ff92df289e8f8d24e3c967a85ac7dc60393b464a9c710b7939d16126695ccb851f165ff0f7dd687f6d3f1e785bc65036a8c3861c8389a7c4d2f2eba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha18e0cb9c9763988f3fe1e17abb0464c5bcc5bf5f005330c2e7323d0860295f9b0b1e9cc35d48f6216390d72495d43e6973e61138cceb150d8e4598a6ce1cd2ee5e73788a632f5dc88b47b3f0d450478961f85e0f7efc65d0baf57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ca10a5a8aefc9e1d30c95e35231a465c04761fc073e95d25d399f4c63527ecad94ae9ae3aa09ff63e71b6a8f6064b5eb5d87c89a7190adfa57bba6113696591775c23fa2792e2a7ec747e3518d9f2dd419dd5496757e44c8b45dcf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbdbc143a32a1da18a7d8433fa0b85631bde7b8297c48b203ad3921839eacc42c6819aa6a61bdfd7fb999ebc74e6e7be455e137883c9ff7c7814ee3a4fa8f07db35fd528343c7e2c248d2572c6a8971585290c8956eb4bcc2771803;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h46a80f4b21f17a3a8b92dede157c457da505fe3fbd6384ce54c94ff9b9e665281a55d11351d444ddf436d9836af3463e1809af9e4077d4dfad66beea8206e911d953a00bafceea9716d2088fc969905c8fcbdc49b5c11980f5ad13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h88a9aa3bc566afb8cfd07ce719ad94b9ccd34c0fb1653ae4b6df7a20863dcdd882b89807664cb653aef01e15817c576dd85d1249779c9f7190ccb85d47963d2e1185b5cf121322ac3c41cd5ac9ca4f6ffc8e7fea5ad15fba241a5e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3c6c38ed382a08a8cd2e33289b14534a3cc13986d9af2120dc29a0947aeebf560809468c5ce18608f065244db0eac78f9c8adab1aae0d31a2d03d3f760122c248107baedacc52dc7f5cafc270a154b07c6a233d54a2a5a8da66d91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he155e2543267f28099f8571a1766ae3a99af020f375cac02b8446be547e8839c92e59ee42b32a82ab99a9b47f9a8116405d516653df3365a54a7467cc3f5e2190f48135361607e438d294624422c521d9d12123843aebca88dc47b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1681148add2b51d3ff6dff442c6d020d6b03a82305e6397495db2269d77b8504af411f95ebd86a0ef38966efd4425c748587994395469c2bd657ea8da29650b0e58c63129787d44eb5701cd7618230a259d7956c6d7480be1e6cde8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1832a080e3b862bf5160a821d35bbea454bcc7973080e33d23ec43d4ee28da8a15451e73ae8c82f481f52eab68133106e217b9f8c580cf9757e7db78b43df6d2435a1766300860d99f4c0a41b775948b89396fcb7a460080ae9e0d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hca8907d9be0ec6fe71f17cecb25f204b855389e2951a86141842901951074a4a040bcbb8c8be947cb0d664c32f993f5c73577ac29e342be83e621a881592415df4344a433d7a1d96c55ac0a0548ea6488aeb30893579848df612db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c0e5945e64ab25e620a56a0e0af77c1b9280c35a007b998dd3efe6933e2aaa404104f75523609543750526ddde995e15a63c128f5bfa7201557cbc118b2bf5df50a4e90a829af7ad8f1af3b89246d98b1f1cf5dee924c3c8dbd8c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h114ca0e937a29039b39075d1bf839bcbef85514d5649122e30deb4f4e9a935d21015a4ca4c7d101287da6ab37c22542f8d2ec34fee1408bab1fc74a2f05182ea2b13e68ffcbf1c7d7d7e824d03403e5c27ad889255a077fc7804280;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14b1fffdc8c9c934a4d1a85f726354c823ef7a2471d808b152cd2161f834e159e6bd6594e650281d61bba52ace4f5be355f72164cefa156f9028c18b01748d3f5d8761a12bf6dc2d92c91bee2404c124a242992ef25b7e12a1a816b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb533067f48f2ed859e2765751367bef1428bfe9b5f55c8f2e09eaf06b8b33e36da306cf24fb6c75b630aaf110c1ff169d0ee6819f63c7e9d87a0c5b2901d63e15738a4efd81dcd62acec3c8614f8ccc0f3593f089f87a9bf927dac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f0651861dc7dd1d6f180299dd3eba60d8d682371980f0ce6c41110b557206e0896d26ab54890bec3aa8a61ea3f8b7cc2dd6d00fc86479f73573decb30ce0bf7d19e059e0de6501c9fb483fcc03b9c1d028add3b14d93af5055f49f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1cf55c236ff33edd4d66fca5a22e7aa5d0e90528e374e5a3700e016f9ba99bfb43ec99e6c8f1f1c5a28283f7a115719c3ac4d605a66d35fd30f837505b2dba1ceea7c441f699aa1dd8145bc939ae649a48879dd858a3000a5380e9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h5ea2dc687cd95e4bbcd31b79a7d1fae393224cf02cb83310f31f1ef6e9dd2bffbb12cebf092c8a001a028f0be79e70ed879daa1dabf8a7a957a868706cd89a17642d0a739aafd31d4526bd76622812edf379a10c58a471992414c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h177439db2eb1e8f9e0bf1728ba4000bc80cb0f03763dae2ebdc54710f3df02da6c7875d646538c7f94891cdc4eb6394b1642e8a16cfaeb0487758d4d7fc2bd2b1326c1adfe657059fc2d6670a56a51dff0756494e69a0e09531875;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h12095b42f5452296843156cfc50cac87e6b2605bb132019f7b213472c9a564afe28c2e476091b9dfb6a82674d72a8c515539d4602e8c8df01797db98e96d60fe9dffd2eaae1074e25a0ef8e9952c61628650a31b4ff549a22cb4b04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfcc033bfeceacfc55d0aee1816b68da589665bda038664a2088c7fe1401565ab6bbc83a7927804068353d710cd1b216ffa97f3006ed719d9e839d5f97464ee2ef6564cbf5ad6fe208e5780749780c8e573ccfb3845e20fde65a17a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1695dd70eb61c58cbd919f810c31f2fdbea681511c84db27438681f428ab84bfe72fd66f99f648720e5984ebd02ec352749f0f5e3cf3384db9c534c6e666838b53182b6de4f705deb531bc4594397200cb074b46e44a98d423b7241;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8bac2fc8a271bc3f0d3db2762a3739b4115da811e03c9a178da01172dddbbd315fcfababffb1b0390cf4036afa6ee8e28ec0387f6b5737ec8f7a066a7f838fcd869054a13ef46d37b041d7033b97a13dfd6e0872d9cbe52dda805;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he1d08cc53cd5994f7fcfb329c84c01d2cc95859358291231bf25d9a31c89171074a092aab28403304ca06954d04aa83bf6bf07f59eb60cdf79b49d65ef433426a812c04f7f6fdc2223ab2ceadd603cd77fc0939101200490ff8b57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1192bdf90eb9a70870116ba4b1457a3d1c575cd9d44c6f53d895bc4728c9b66059f056d0ea99663ce9581e37786802bfec3234a5f8db1939ea21058e9e968b5f97c0646ba745f375e3fe5bac900dc1c7c158a3bd760b201dddb930;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hbb4b586a85858d6d71433afa7f452e84c9d0ff67bc76ca3c127d6568ca2e072f62baaa8ce891cfb3d37c7b98a99e8eb47d8406d6fc7b4caebd08ba336175dbbea7464c1dedd584f4436820304e518ac590b8b70ad128b913bb06ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h36fdddd62b066bd34b644a9c5af864dce186c7e28aab1a1f12086840018f1356f2c3ea9ef8e21a660a9ef0c7d54f24a057066e2da2103c575d43b4074ab202fa65961021c01b3b8e50782f22f72342bb03eecc534c92fb54d5c9ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha8d649689da0f2dc9ebb7c09d3302bb7f62e185a330296b4f6ba8c1dcaab229248e59e74ebec12d7937e168fdef0d2fca899165ccb2932bde97640f3f1a6c0fc276c579e804262c2e38efc761fc5caaa25bd82e0a7648c361f42e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fddd1a77572a469755ee136d0eb64200cdaa1348fb53c9ca49a1bdf6976db16c82c7f109b912e569d4c9485426f3ab07bd5c880eb421b77b271ccf382173b43c2d8482f6118bf0d608c3c04e7f6b3a24348e999e7dd38c39bcf04a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcf3d4b47ab41ca20516cc3b4990fe0ca9e10da51b89fffa2e7ec04d84e0f498f3f82551b67004e9b922b32c867c1a6d0dd1cd3fce7d2f09aaf57b7f7e4a5bd868c68896eb573e8f7a134068ca808b8a6b9da4e7241e2e31f30015b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h50910bc9731aef48a95ee4d92a581e17d2c4675381370b1f4f99b5fcb92d04a9bf76a45efd4d98891884a3a506e40ccebdbbd669440c0d6dd2d3b167e354bf4c5cebcf5d50845bb8a568d3aa0bcda13f957385a3c407e0ea250f5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h3b872c71c27e3989db5593929716c123422a09b92febcd9ffe8a177585daea9a40dd3c91cd1b9b525b4099cc7d3b0d491376bfd563d13efa9a2dc8758031e28d8deb7fc769cdce1d32ef378c523d42512d062cbffc566fdf7e94d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14528fdca58dcff8275045a3ff00f733814059b891467d03b654bc72f20f3c9ba63d511428b11c998164b9785173d821112e7a16d4684c45a2ec642b2c598aeeee4e2adfd220a64c5fbfe717928968575aa8742a4c6a71e1198a9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h175383dad86d39c7858ab5785d92a18b87a08de1a17d2322b9caa806e41613292ab433d240018f892aa36f9d07d581fb7914f693b7b2375de1b1c4211733ec2f11466a179adc9f0543ae5f935667087e01431c2b1c7e8b228029b2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c9f65850d274204eab2daf5a134852cde54e19b823a609eec513e43a9400993a0220749a4942727a259d08b0938800c607fed1b55cc4406e7e00004e5d199d3d2d99f423059058871c886a955ab4be2af6f222031201357ea17fa3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14bd4bf96dbad853a4bad518145373f8ee4d13b8aaac82d41ceb6abf44946969f5e67244c384e25d09ca7967853b92a49a7eebc786d7a6fd9f2d0772852b6e0a62fe267efe643baabfa36254a70b3665e6c4d63c6d32d61a165d129;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h165a483592b52a0e7acbf8eb1d8e8430eaffa8f52aaecfbb392582f1c01bb4b11c9c4ceaf8d2ad8e21179cde40101d516402622bef97dce2e4367f321377c9251fd5c7020b87dadcfc9db21f71291171538ace078d723200a55b0ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17349ec4640dc7f05db787707e1297e051d585d2bb53700b728ad80d7c29664b881b7ca67d70c22a889d85576f4c44f85838c89dfe98f23750a9b7be18e0eb8717cac4196f6fe74b3a7687b3b8d29ed649bbc1fc10c0c8caedf92e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h185bfe21a615afc32d660f29da79a443e57bb87516f846bf934fcfc7a3f6adcb8d4f450d2703019b5d0a51b938128b0921a45f7ca6594426a55714c7152f0b8e8b14a6f42efb444df71c18952b5edb3a20ad889a15ee4dcb20dd6ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4f0fa8d5f4ec076dad54232a7d229c36f294f354a6da8da0fff02738e0f886376bcf660a1db55501b32a2dad3f38ce0b8dd762bf86e5ceb312089cd3edb023e04bbc9eca628482ffc44b147dac1af65ed00099ce7618f82f89ba56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10b53b7bbecfe61b537c8f15e002956f912d6aaa68acb6c142c2c755feca572d50efc7e0607d3afd6cab22188d43592a42c3a002cf4b7a12c227f2f10b355f998df6cb8b6af71b034df8eb4fd0b2f3819fd6106307e5f8178bc9cc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h121ed25cd5b3cddd53b24b899a05af231c61fd290a73b13492b1f42c52dbdb1882dd11810caaaa459ad7d7fe4e3a566920a8255fa3dc05c06d64ef751886aaed6f4314b901c6ac8854fcf199fb649df90ebc9b08513dcddba4b6889;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1115620478414b28396bcadde545986b9e7b815ff9e00cbc21c7bad88af2ea503bd76cbbee5a1eb0b27390c2ee4e24eef0776600a535b2597e4459e535f1029bae7e78fd6adb748afe4161483c932a270b30350d7b102be99e4d975;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11acd1eee39e00f5af6d9efeba350c91f01bd3d09a7e9edda5ef495d4ab77d67953820788b52066b6c771e8ad496afab3faf8e63dd6b7d61444e294a61ccc1ac246b1801bb7310978b5186833963c829048dc63164a8c2a7bb945fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11cdca9ab9e0cb922642eb0a29cb40c7f7abce780a5f261def2b4d8be607d50b6540f41c4fc1a5d6ca0c6083d481b5b433996e88db8fcf182cc2d45ae33ff006eb7c269c5967f6329b6ddb0f66513dadb0de22f6a2265a034ba6fc9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hcf0bf177ebb907fb1e4d6e1cb18f739205133f588a0cb04b4dacc054fa5e5f38e10f82aa9a8f0e892026732c5eac54e6fb1479b527f3a15a04b1d6baf642119f9c6d6ca03b0f425632ab8187c9801d35832a1247820ffa30a23712;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h4c47ebd48d963c6a3f5b080865b3920019673d0a238d428e03bfaa88aa3962f0b93f0a7c726b1ec65ac36cc80470471403e3a90c1e32d85de842a069706149571ec8df458768c2d0e251cf7de2b9816e5f2d6418b9a5648d97f7f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7fd6313931798bc0f699ad0e980ba10bcf8793c7f9ed031d2e5a5fafefc92f42994568773843614a810d20a5a912b6c812e13d5267bf29cf53266add044b449f478b7f30cea8bb38c012b4769923d139b68f8cbf9dc3a6c6969e09;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f00fa9af7dbf8d1c7a3e3784f648a6d47b93056d9d0d5ca117dc9b495b466e7b6c57f16befd2e7ecb0117158ab1c4511dc325664b7a22854a01e593abce3ac4d5595a969accb7c9f8c54367fc619c8a33b53730838812e9aceb43a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19351799a2078f1ec0116068af6bb019e156328210c2c9a65291c479460ec51732e2a9b124088e7658f98b92b0567259cec4100c32f10b3e174e9e2c4ea8e6a66f49015d83df97b140e628b83e279c46b40a25dc1ef37a36c4fdb2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e744fc878e7a7be2c4581f534c0815da034c86c13828ade1060748129c7ca4bd7d42d350d67576e5bbb74851946d659e539109eba16695c3c016741a8d25002251f753a953f6c04ba7d3928d06b6b2209c01e9cf01efb9a3d2d604;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e8bb1e8834b39e65f688895095fb78e90bf4453e7315bb62b3281c139fb597302f2b7f365ad6dd0db481946d580a96fe6eaa3592e74c7c148b1acccd2ecf14e783c655f35a054adb02c059506baf8703aaad1f60b5e33af086b77a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd4ff1801e2c6d2fcd4dd6efcf64e6a7b1b0112d027ee58fe97c1b665c2832e7b6ba9b5f0288a1e50b3124664b073fe57fb8a7e15d4fa2b5d885d78cbf0a7ddedbb7a357c1fd8a40b76908f362600dae03811dadbecadb0f35efb41;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h33f0c5655c2f950c711945caffaf7fc1b154667d364c20cf7573da70ea3ed8eda7c257f7b8bb55f22f98f4c7465aff98890fac6666087f47ae15cc75f82da9173249d9e6c9c2dc55242a400bc7c19aa827094c425ad234bd235df2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1fa914f75399b070a46a099ab057b120d731603f7df816dcc664c60072bde571864863280842cab0590b3926dbec5794d1c2de9690ee9103d544347b3751d33a698972d55e1e37c4b09f018b286155bf301f5c38780cbb15ea38b9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1bed8a5779a5243e3d3fbd83abeb0cff56faed92c193f6496e9986c88212b9418f1d13cee9514ec719d1fbda932e35a43c632b48b88bd37b6ddddb1d46ba0eb3b69100c7083bf37d9fa8f1155e03e0d8699c661a7c3e170af730a29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h2eaf85c18393913cd901ae9ef56d13f121f4a5731c7ab4f9ee2599e5ec102ea233a644e146ae895927583cb1d2e93a142e885ad7e17f8b24f5ecac6532a2b3da8f1ab47c168e70467fbc3f92dc0250ebf5215aad0deeedd804a55d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de30888d04486ab39321c8a639457b043c305ae6a464390d074299b46a950b2f3b734a0c36586864ea8865431921c38a787f78c96766bb5f10c5cb5608cfe62ace5c904f26241dcded5b08523553483e7b948c8f52ec49b4c93a16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1db4abf229398c1fad22fb88732fa17d5ee78ab2ef626529a64e688cac12ed62f3c4a28ce9f4512721aedf19e9fa969cb1bcaaf1ff4e09a7a8ea96925472ef6c6a359cb41e271a0451e9d37e6458d49242f221c9d4ed463b0aa51d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h383703a1d0a11aefe6d3931083f667d498b3456297ab370ae2f18f20297ac20be5298088f40db8df2cc165b874cb227c8361d310a040d9a93914782645866d8aef2a4f3d95bdb98fa06d7f8d0b3bb1d4fcaef7e8e2239c8e7417a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h197b613dcbd4f6a70b0c091cfb6b9f1375eee7842756348594f25f9a65ebd5273dfef511c68a396f45a7faaac0826647a33eff24eb3cfedfeed0549fe0040f68063ea80f62e2fdc08fc0ec02b8d20a08723af3075c3c2e5cc222590;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h41dc0b33268905eaac114a15063980d2c8bde6d9176be22f1aba3b95cd9546131d96bce998ad46e1a7c4fc0d4398c1b5238cb81e0dd3087f814146532b13573acd0fb57f6198d1223ed23ab158807277a8231de8eca3677670b32d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16e16920219412c2f86b68c9c092188b6d1ccfd2ff5aeedc161e8c200e98580100e28fc9ec66b20a6a9b2a52c23d4402e85a8a07ec70017e9b60cbde96e17c2be57a5eeb1b2be08c996a63e6063fd2b2911ec21bd004342bfe0858a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19160973294803c69aa8b6e0082ccfd3b5abf02561b31a21137bba13c4a6eaa01d6e339420dfe2755ba23cb1c043fb6a7a66aa235c2b8d4179273cfb9ec0b0704c999d84fd90723e1af04d0c6eb83420791931ee1e790575107b388;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b85e4424cb8a0f8763abe83b814397e3d549786c3d65763ad50e55b474fd4656eb68446d81e64f239c83a633d3c8b20f78214343de97e929a6c512f35cb933a194102df06fc14811b5fbde4af24d0fb85e858e525af449ab00e13e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19bfe5469b8316c4519acc8cea7f6dd4ec2ac517363351fea98c7c9fe5817471613d732fd430395a013451128f6ad78b08cf3f0caffcfb9d28b2800d03d250fce98f1da0e5f5c3f5de6c58382acdfb30d177cc7172f218399ca7312;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1628cc4f3a64f1f7a35d9f6a484756dc7a43668e1b4f81110bc8cbcbaf58d730fd46bfaf508a7211a65991b980846dab5b1bba2407c8bb20e7ba0db018aef1fa913bf3187aa0d21153d0f5efdcd27978edea7d1ed1090507c93261b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfa20d4986a65a5cd5eec1594edc0a2d531621c07a4c8420ace6c194963fd867182a3f12409b7074cba081f2e4bc2f182083ae244720569698223f3bc79c744970a1886a25f2cd57cc75ba72eda7b7043bb0270f29c704dbc894862;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7d28a0aaa4365f546c218a9f08b8271dcb78a2eb13c2ad24c43beb7f4e1154750e42531cd8122de0bdd98854011ad5fc2bdf71ee05037d5250e64484a4e41712716163d2eb85599d3c784077d33157947358ff74b25dcc9f2436c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1635c1b55d421034437639aa31faf1d56aba697c5844b471df72ea77d5ede58029de8008a1e575455687bafb6112f65d90c817f39401062669a03142f067ee0b077aefb8185406ce9849961df3da1accfa61db39c18e91e7bdab5d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfccffa8d6536fb2151aa4f4853c85fdf9d2f12c11fbacbabc6c51165b07578057d02a3c2fd2bab60532beae9b61359e3de84ecae7a04274111ede72384d453e63243abe414f3c4e53a5a1bc4f288d29d7367ea298c22a3eacbada4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h27fe5f144728473265dc68192fdcad8a46c9d100b99569673ce608e76a9180eebe58da0db8b35e3e4e0a82cca683bfe362fc6de0f5201d299fdd72f49397438a85327249ec935162a0ec83849712df6ab77eee896c013972d8c2a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8b7b10579fec015d62c07ee94a7d86053009e1bfcf474fd173970c35922436b45b52e1509b39a3fc6e476cb5624c70fb9c6c2ee417b71561567bb3cc6bea469435ea3377a4aac93d5722c6bd24fa2dcfc5b44ef0e50a5614bc0db7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13dfa2fc2fb6be166335ff16849bc56a176141ea1bedbf23892b743347785abffb06fdbd7fe811af92c0802d7827a494cf60a7d71d49722dde67cd330e2940f3c79596113a217d6f19fd5476f422b779ccbe3e651429790b98a2c3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e0ff06f3b64ce5542396fe2e38293af3dc0d3fd7e4b234d8729172844791bcc75765b0fad09ee629ccb2cd49c3105234b5fe2d0950aa2f62a90e01d78c211b125faff6231d4d677b22bc1b7b2e8583f7b306f901f2d5ef6168035b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1340aa3ae82c54498fdb22e5a509534876c520b7a057d4be989190446e9e07c356cd2c4fb33ff09bb7632b9b0af453784c3b5ec854de2f9abbf22e4b28985323604ecd1a14d6519e6ae50ed080311fcf675089b0a084c43bb7480db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hab3b00fc122c801fa3d024e3fd9c914fee945686a281ae85b830327ed3f423e80b6e278cb58fbf32b09a366f6e1ec275ab4a9595a2f6022d18b4e4e62d430ac5dfc39ff04ed6137daaf8ba8204f87debcd1174b5c114529f076cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h420b5d9e09c358898486106abdb1d079d6686fa69307238cf14577c071e55109be45cce55467641fafc50ee1b91fecd0f16d609d1c7151e586cd6c06317d279a01fa9a6a6bb3319f10978bdc3ace2d9466f657815ef43d6ef05ccd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h121698cb23c1373339a5467e799dcd52474c7821b10e0dedc7751d790886d90744194858b2d4a898f6184c0788d4a82227a1c990b4e3e64932909d0635ed27b3f5425ca97ac0e7ad0f322f11b41956c473cf3aefaa1e818ca4b827d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18d9a7161ad442ef307a62a65d6756ec48992f93966b0923f0a97a9aad3573e6be951bf3d3c2b19e869a3f3c65dd69da18c3b69d01d05e9fc18dfe1909b9f71683b5d1d76029bec685712c0a3302a84d7080e2816ecdd170981f7af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h156423cf5edc2e5372c6d80679cdcf812622f84569e70a44892f4b674db749d6f0a021741e1102476933563f1b3f86675860dff67eec730169046707927cc3d81bea1061c93f1d4696062bc72e8a386487bb7b34f9d140b571fdf1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hc5c36471d866974fb217789ac4cd562ac5dc74f3a7ec74fcb2c4f6e163ada2fd532e05021847c364edf55efd60ac9adcff618fb7cfc8e297a306f67648a265686a5f1c0235e10e6048afa2d7ce7c8b15026c7ecee3bd02e2ffda91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1028b08b68c585c6f1429ca107a64ee3c5389e8245775bd895db2b297f04ead6eb241189dc133c8be55fd9bd67225454a715592fbe5e5c9688fe9fa210bbb216c9abb6b442d01d28ac7143d2ec768c2cb1defe980ee7e4091abc373;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16632eb45c9b308cc01e796de26b15c0952a8519b9acbfdc9981c25243d4464da6414b1e41aa5b82dec4ca0570c86a1ae00e5cf4a19b53a40780269b5ded67894833d53c2307979b73ac93bb390bd50657f971f4671237c7778d43a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h51f0253ad1e69217bb5245946d44bae4763f9f3ffef98b49e7c94610c277bfda5c22a6b9743dde9d84b96031872ff00b0066b37a50d65c26ee8ca89c15de33f3be112db2336480b1db376124cf6a01cbda57fc2a060711f7f05280;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e29133c79560e3793b0cc9b5347955efc47c81eeb4f71d8855e8dd74a61337fcd9d07bb70ff4995c38ac1d7b57838700a9f6af3c0199a39f4740bb97153df4f149f42d438fe176ab4099814ea4c62f8dba1e49ff9a27e9e38e80ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1df04a665b1b1e224810de6bdabc238857f8f8d757690cb49e38aa848b9c45108f9f0d7f7e4390a8221f031708f935266791d9c38aacb7a6c27b45db9262651904b153574792dfebcf3fed418fa0eab7143a93eb91281cbfec15b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb1d1997726433047cce6ffb9cc45ce77155ac9f994dc7aa9092a06289f14aad1c17e5d1901a35bf2e45b21b7a51a2e2b6cef27863b1410a239662bf00198e33646961236d78d361193cd75ca866c62517ea9f4a2e7eb43cad2fd00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1de44dd004045f02190f9e679c6f68579a24b55bbdad829476e40cdc19ca7d0b9f8e703331a867b5fca5a87ed64c60f92512ffe7c13752cd9fa89c1e4316f771121d40fcf4b8d4a370499843359fd906c8cfca286f5b1d558ddd82e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1ff83df2564ddcc577aac24c9e792fd174cab011be2ddd736e2d281fec70636b8b2e287a93dee21c05243af608eb7d2aad17153474ee96da1f0bd2383d6128010ad4cb74d0beb11647b7f3fffc310a4cced3bdd84d5575ac70436cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c052fb764e1e887a0f85edc62be3b395fa2580e812cc54afa859e6b91f6c96e7dccb45afa8241dc159137c37b9d8943b97f280a0f88826803307d74f2c4e3e19c7d9aac51acd1d36e416d98a101e761ac85cb700480a4d206ea5fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f386a3e2337906a60865c6d4f7d920245c3f9415609fa9d6b95ac4816636034158d37292ad229a9eb84e82cd4b5da2c50082c761d661f5b44cf460368c74380fbdfedf855487154c4e5bfc41b32001cab6c915faede19094105592;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h824b98a1d01b6b360fb1ebfef71bfa2d4d28ad5745c23ddc90382795c372307c421207c238bed2a140fe1d95fa62ff531c3f5e13ce0626ccba0690bbee711287b732c24c8e2188f82ee6143e1154e19c180134ee7afd976763411a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h99b43ae8e07053fd491c6f27afe39f8018095d925df966053110c617e61784d04139b164d6b5efc2a42585f98042a2162ffead6277d693f3543ea12523c7752e513ab225c65dc0d7dd7a97cca73f7595a9034ebd6d7d923c7f4dcf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h18ca7fda7124e0eefdb8bec5576440520bcf12082a750da5cc4298aea3d06653f1ffb73b6081c696e26df1c16fb60ee8820510bcd299be8c9902be8c2749c33b98aa2618d5f738ad22a8322b2f0f3feae61f305c4656b12e6e585ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h7d733174e3d749b4df8b8b1be076bc7a866373751d99c29c1e426a98e3b1719740e29041a43053588773f93a28cd79627c8269b9f084f6127b4df2f575427f7ba241b0618d3a4c8e9300a6f1b901d88a84cebff391e990d81d536f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6593466d6f97a649981807b26a582379bde8191dfffb30c22ee1d03e095c293e4249bfbd3ec47d37989e16726eed5cf4343892732ab4aeb016604e16cb2896e98ce27855b07c45e5ef9fe172061634774fedfcc9868ae9c5220d12;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'haa010380234008430cb6e6629ae44fbf5f9f7f2ff1c5e87b73931c06bdd9110e7b7ba42fc8bd8fd21df26ce57f93efa6e1714fb1dfc14e57fa37dd5c8873a1683a505fac859b439431ac622934339cc9e9d3d54af0b271763f6862;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hfde05b9af3028a2d72d89434ac3b89e452884b3a53638db16ac6de2c5b09aee7ede9dca49ac96cc62ef9523fe07fdadf853965fc58dff99b82c2fe3d4bb4b8b7941e17c1f6eb5bd2eef0afbba1201cce9d207f93f058267f6a9ee4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16cf29e41a0b8f5842220ad3fe1ab6c3e26fdfe21e41bedb14a09cf2ca2f988d66ebd42fab6edfd958b7559648f5f263251eb832db1c8470b157a1b121fd49c5e80e89a04056a940785a7c8594eacadebb7e37bc1d296730c8984d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h15688b2246a101e82cc4f270c0eb14dfd920c50f7537572ed7683dc2c54cb938f0fbc7957867deb366c0d9be0221f0ee63a8deb8d664f1c7e35392570cd4a2c260aeaccd0133161cb9c9eb6ed480db1d375c981cde1d8de79f57185;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11e7364904547dacd42320fa59098b8d67fef32a72a5d600b2a969a06d3ed40d9ca0e7718809c5c48ed961ee6cc34cd7d2f8f9221113dd77da3a258f16f7940203b08515d6d75748c69fb383758785ce2e3a5251c23437b49667356;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h8b98941bab413305ee08f7b98d38c6db1757aa605132fa7228e996c5c44ef432ba8163c691b205f278816ee7a5a395af3d6ad036e7e3b5025dc26fec9e305d2f6eebacbf106c82359bfbb3120662254ba4117319d911fa20ddd157;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a838ffba2db5ff28d3edac4a40b902158c1c59b814c9b3bfa6d7db2f780d25bf00014f0ec0e7d527206a2a972513693aaa279304100383aa165efd2445f4c4bba431b6ccc9914b7f9e3e1f4b8d4d7c466d5fd55c4081cb1214763e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha72cb3bd42a176469cc9b9750276aeee2d5f06ebfdf383e5c8a45bd8c1a526222d556be7855321da8c3fd142cb8c38f4b73c27b0ba631bafb92687a69186337faf7fdb09783cf4c868b9bddc8b72e8c5c76e5a24fba15a21d283ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h13b005fd757c98da59373d9a1e1862b8c0891ffad4b7859ed851e96cdff7445cea014e56154dfeb250fea302c99e6ab051514332c9030012137bcc4e0fa4db564d15bc0981cd29c361bab54ed7fda01971354d9c059190ff1088668;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1becda3265e7c197bb78aeddd242d421836101033cd80a712d0372203195125ac6baf3068b12042d6d90d91d5c02e48905587c2bfd0aaa3124b06305b36684c3ce1cd0ef671eda06d201348e176f481d3fee14017eead731a82c8d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1c903d8812e902dd2dc605eaa5640c9a2f53e2148233b3d453e40c0f10432aecad8f19f68bae42a591cbcfb6f630ea01212ef0f8d6a37dcfa84d99ec78729405106a0dec44478b1f58b4861519eefb57d89b39c96c08c6b2bda80e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h471457ee8e328b635cc13fcc869c13b478c194a47998c2fc5ae9e7e49b1b7f789a4b12ac95f32e746099427ed6ffc1594b6df6d9f29872aa61a909e5b93f5f287b588349ee00531edaad37320e2787b22de52f671f31541413d9ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1b7203b24dfd04a6e5fff174d5f74fa0d6bba06874359411f05f03e178812ab1e0be13031f7a7c917f0c9b782d63a12f442f0097951e8552eb5f02d5b30863f82bc68e63c368b481fbb3898b44a97f1ed91001a45c94741fea646fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h19555ad37302679e72daabf550cc1840a8b768e19b66699d94a49cea59d6b7b5b5a007399e776bf90e597a22e3f70e00e4bf67180a0d798088e4f6e0f80a99b2de8727e86a65fe04c4e47a7f6ec538e3af00b60029e4e8d75f64c23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14018758f8251dae2f9e8853d6e24ffda6f1f15bcdcfaf42b7db389d4b8c2ff456c4846ce005215cc22d4d0d4c46330b30c78b0ecfa8dd671342752a85aa77ade28d0b55818c25cd7bbe0c15bcd9ddf8132eec5191df7e6e13670d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hf34487799484bff3174cf3c25d301d7f7e5f5a4367a1a9c1e1e2c5545ed78f41f1eb8cafcb93a5e92f12bcaeefc17f956d8ce431a29e53a567188addd3689bf32b0ec252a52a428fd476108616463424266dfa047ad73d72a7ba96;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h6424eb182be931b4df3d8a7727cbd925b75e6dcf25f412076f46e2c8885bdfd53e6fc1347380d20480ff55d476be2007759e07681b5811dd81b7b2bbb4cd9edcbc7db08cadfaffb44fa0acc0312921419c5308b761deec39df312b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h11b3908ca42df2746ed703f4873d9d6b4bcf8e9ace810b72606d1482894422864357c785a7a073a35fda2b0649211247a4a957fdc82913d7dd521892429a769fd8bedc440697ba6d1fcc1a99ff8dcf9369c9e01b42e1e2040dbd2c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1827a234c28e5119f37c52fd902d3cd9b06f178f2105f5865803d04162ac1e0d385a8f947af220b5800d6e54c1e8e7864dab880f977ad7bc5fc40e455222bc31bf4fd939bc85f2e6fb52f86304ac044936e50666d58147517851eb5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14168b3112b09e392aface005ef7a7fd59ecb6dbf6338cba97ee44a198172705716e086a8c48a2adc9a49e62345d3cf5fc42894b6c4afca1d0f44955333250a0061a4484279ef6eb91bb745e8f9213fc796a16af6cc529d54ddeda4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hd6e04faba71a2439c16d39de8f32e5f0920cf2452e741882c356a02f47fb4d532f891e580266e700a09274660d6c7e732c59f2d87ce18b9ffc9a77eee54c47c38d39c5f873aec73fd3148aab51759f5b24eb0eabaecd856ad8128b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1131d4405bdb4a5522470011df98f4095d1dc485e2f5d9d67c8344f47f39bbdac53f68dc2d3f2a3598517e2fe78d3c9f67b5289a45a1f923ecd7c807e7980752c9d1d5e6b1652a4d9f48a72fef4316c8a3fc1cb6e4204a14f543af7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1df1f9a3054667aab0542f8e96d6ba75f08ca75ef5873249b5a9398aa2b5371a4af118f1541f770083afc352361845a0d32c5ba951c59d4ef9f9333dd368a3004cbd71b653ebad6aeff9ba8d237064fb1b2b772770645bff50f6efb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'he61c3e14493c91c48c6e4963daaf71126039a0c5c1998d9a084bdf1ff012458126034f7b1790321c3f74138fb64ba52166f553cc8d86cd82e7ed799679d3f50a9a6e37b71745e3588b1417806f49545d90ba97fbc747c57c92dff4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e7b5139b0c642866c41a250e84f25cfe600b3158123ad028f9517b4e7ede9f65df4844bc220b329add15e06e94a5511c3a98fde8c4b60e63dea4f44d94d9ca4f0448389480f16d81bb16361fff0e0d43a7a2b5e10af896c826d8b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'ha20fefc3120d7056b1211e8499924273818e5c34871e4d56577749b5bad17d1aede00c828aeec1c2dec1b0a73de29d55a9354c0affeaf29b1a2a7c3bc49f959893a4b092e718fad3f0ced0167b4978cc369108d1f0f947603cb60e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1181bf390d5c87ee7f0130926e147f4f1f80386cabd0213c62f387a706a3d3a628d9c969bf67d6c8b865c8f06a92c5c8b42dc64fc6b056422d18b2a879ce879d5eb4f47df5da34126d2b6e64c0c4736697801b1bf37597b71a4afb9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h64753c578f62428115fa531ed8ff89ec6228edca6ff8be62a79a075f228367a72ae070e24011bee5eb64be5edb116f7b8b4135aa597fac602ce038db4effef70df3dc1e3220e4a10698e878a3db32f1e45f313e7bc09622650f993;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e410624e909e0bc083a54c8e66fa403cd4b931025ffbf3f2495c4e0572a5875f60f7617adcb79d109a66e7d1edd5ecc4d3e8259f813d01745108deb5b7df033b07bc7589092091243c888a24989f6b5fa6d7a9317a35a1f5535560;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14a9ab79058fb51cf5dc2ee30cd0e11e95c656e81d39a702ada2766419d171a17f9b37b4b60cb27820d185e94f8a9495672e170c7d98be384a72ae75e83e204801d1eda94cecd3b45f10c73405ae09c35f855b96302ceed6685ea3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb9a07076a6705772a546e36d431e41ed2a9e28957b7f92ef9e480a5aa45e67b83e3608c1b68cdbcf2d3067c3416ec2398d773457352cb660c26ad31cf9f620261740b2bb78cfbc19f0d824f10e2508c83a37990983e5eeb7e5a43a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h84897c1d840d7afd015d9b8599fca36d3489266b1361f9f6173277a7440b7f7008b5bcb73ea64e5c404e739e6294b1cb42b8b5ce886a5c4320960ebcec9d0e3d00de1fad17420111c38c3dfb3e9cd9f739bbacdaac6f23affc1d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hb83c9d64983a861fe664f7720457c2bad62427e5582476df40372ec9cdddb228054887b8977936afd5ac764937b6054fbd6dbc92ffc56ddd997e19c5d256caeed519b6d7de336086697a7b3b78f4f4630c326d220cd59f118d8522;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e5818f026b9dc8495406c5fe843c932597df994283ccdf05328cd3d174c48100ac00bd2274aba04373f57bc9723bbd819138fb31680d1ceab3c7cd99704d5366ae5dff220ce90402da0c2621e46c1aa9d27562a8c6d094e61245d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'hdd76870d6629f6ef2f629818b0d2efdeb958efcdaa5c4059349c1238cccb5a95009c564762d787a1c23e758922abbf124e568a1d9696f14a6982700c11a5c9bf9aa44db02e617b2138b39493e40719caa9d18e0d160aba803fddf1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h51e6cc0d30003b5552c0cdba2fb203bb1ac1eb187889a19513303a8aab1c8767bb0e71df1c029e6d93b8fe4f064c34067e80d68b573b9bad2d0df8e63a5722a28b17fb8d81b78d265bed77a96525c3cec9c0717dae484cefe059b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h14fdcc3053921284ebb2a949f78a1d6d3cb73229b9b4bc26da1e8d49a26f0b876a6c63141909c4f0f3f78ef1b87b837101c7a26e8e58bf0c17f443ec692cbeb187dd2e376ff5f833b596a5ca9d4add17fa5e6107a728f1d5f988b8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1f91eb377463dae4d4f364ee9b1e804a711317d86c790f960d9a949a681c773221592cd807938bef06d5c3ad75e5be375a7cca55ca31438dbfb72ed59eabdb4875ad62dffc6c76dfe3904afd032bd0aad327c49ce48a7bcfa4d390c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h23e23c5bf233926b3da716287774cb01f3c94365b1c45d0f55d7b9d0da50cd312698ff3994a30a04302ae0bd61b3f28e75a2a22b8a2075031ece6ade476ad0cd20e3ad4a4e072f6a297113f91cc9260f12a01b358a987e38ae95c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h10519fa04519f5516b7c67101441e4ec3f0c1ab4c9f70f5d4e262c3671c44466b46a8c0d865b402a719ee801f4b59a96602418410c6fe7c86a048ee307a489a2bf8322b69129181a12f66d6c8543f5996a279cbdacd406e5c3e3124;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1308ff5fd50134b2939e11090c66c441a6fa55f7daf1f9271d33d955a6ce48b225a1178abad673434cdd9e1dd881642dd75152073e3d5ab96d7384314072ddbcfbc86fd2bc808822a6c3fc453bcab890d9a3ebbf4dd4b0af0a83c33;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h105ca0099cbf1e77fa24cb0d250044fc638e28466046d79d3d635717b95f4128cfd160bcc3d1bae6739fed770e5ea3c269ae9156ac442a2ec81b26cb225655322d98202c7a3ef7fcc2d6b0814feb001bbf6585f3790905ac72e427b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1513e81a2f4019988e700a4d38de2f6ee1635032b70529cb2cb8a29c25fb632f2ff40fe2530f7492e12b2ba4d418470ed21aa5e4b12b011d7eb2f18ea8554236dd8091120b9fc8e78ed24a00c6a7fd17ad872fad0c278f0f35b4096;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h473f0183ee35ecfd9322fcf92116b370bf6427e968fd581e646d98a00e4374c7b0412413a2e910a603674b4636b814c72a845c3cd169667930d172226a8ffd5268400daf1d627942e6af5ff1dcb68448d72a3d843587d52ba8e6e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h17746db26ac8bd1aa7249f66cce4fd3a68077b968801f3f746e72532be9962801ca68103ba04eb923cbc70f4aac7b65da83cd152d059473e8d3287b59a20aaf148600d60f927bc539630cd0caf7dce79b426296341f4deb29a37e5c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h16d0b64e468776ba7ea809aa31304a4a9bebd579d59676f2ab4cc15301b0080bcae1fd8bbc127f4a45df6d9bb6f33e926c98501aa69e0933357340c300fc9b987af8ac0b5db7ab3df8f1a1770805011a79a45a7e76c52206e81492f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1691b78657c38192350391ff14341761387ecc1f42f14c1782a7a904972f31fe263355c38c08d87627b202148404b74d1a985842436576c44d8bc76d3fa7d25037b2694ade2dcd40a0063c1c12195fb9050aa0bc3cc64d9a3c0ffe2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h106cb4e67f75097de18f5d536926b6b31cb7799975e6b4ada46c574580839bd51969d89a4fa9c020d4b953e41e0dea900d9dbb8d9ab12f703e624818a050519ddfd42a2b3a4ffd9788309b5103364d74dfa348246b144925ce0ffd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1a5644f2349c9f5a8ed70c7da2c7f32dad9a583f452cfe6c6782c34eb50f226a576b015ddfc0dbe30a98278863b9faa96be883b30ffcaf54620bf91f6dea808869b792e7bbebe0f57e106853f4b271288ff9de74925611a7be911a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 729'h1e6ef153b0405f7ac8ff973e4ee8222c8ae79f9f08f392bf549b4ca27b6127e8f7ad59c2d632793927e9de9c1599451f93d10357015b46ac0bcd8c57df9db6b1faf9a7c6d90c6d6f0d79504de16ee67d47c7e0b3959fd1190b579b9;
        #1
        $finish();
    end
endmodule
