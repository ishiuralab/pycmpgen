module testbench();
    reg [7:0] src0;
    reg [7:0] src1;
    reg [7:0] src2;
    reg [7:0] src3;
    reg [7:0] src4;
    reg [7:0] src5;
    reg [7:0] src6;
    reg [7:0] src7;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [10:0] srcsum;
    wire [10:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffffffffffffffff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59648161d2c0f1f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b1cf55263c8d2ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6baee08939627e81;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86f95685e31a8775;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef1fd8f48f9919ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec56e0f19ed30a8c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he97670ec7758063f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4a86b2c19f6f483;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e1e0f6f5be859a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd4bba99a318ab0ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc23538b51c45e10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18928d4678c6f212;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14d9294afb5ecb2e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79f49346ce1ee478;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h96e7236ce9ec9f81;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8013bb8e7c2d43c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a5c5f3125f58568;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he94897c0b1029fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h860b63fd61d119e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c84eefae6a629cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he32b59f5617a1cb0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h181058610095db6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56d5a1a948e5512f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h736dda7040bb053f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64c00cd980d00882;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69f5011b92dc5603;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4250cbd3dda58a08;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda9be72aa669653a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hada1e291006b5a1f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8514a657c7ca4c71;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72661da07c733fe4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9c644b49b6e19fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2fbb18892c1a4849;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54d20eea963e176a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h716e583a9e4fbf5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fc4d632bf9b5073;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd413bc34819563d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1746b44592cc6eca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f2c97146c47b25e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27f9b11dcf2ead25;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7836f811d1fed921;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff3f7cf67f7ebc9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd77e173129402a84;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h897317a297ffe31c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35d40be2ed570183;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fa627d10bd092e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h141de691f4de95d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba6cfd978caa746b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c71b94ceb63ecf8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2f42883f598079c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7596ddc0e4b7f96e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h893f8c2948af742d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf22e8711137b9375;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8d6635f24cd717b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9991c4a34f8fb37e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h278db813118fc928;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34399aa9ac1d1d3a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26ed20858ad67b2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha365cc952f03baab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a7369696fbdb9c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfebfbf3de010d87c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9de77f7569bf3466;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5b3f16e70e56d7b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38f4e291a770f9d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34ede00a97cf980a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h37f36c3381024d78;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71b7531ebd6418d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6cf60300af600f27;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha49dffdacf726a05;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb06f6d81c863840a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2251facef566920;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae3babb52c4eb9ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7dc6704066eb163a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26ea446401a1d0ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8051c530a86b060;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9f46bb4c2f19e4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb54d90d3f3b0e94;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5814dba0bdfab08;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1a5562a2e98565a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd513f4e14983cd99;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fbbabfbc29123b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he49f62563270fdae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd2d1d9c149dfaab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76bd76e77a0cef71;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h619e1a560b520478;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6d6d3cff36db183;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a598e45fc117994;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8038680f1818acd3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc88fa25c6d688ce6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc853c6b8105190c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d3903411be9dad9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9f42d1a24fa699b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd612837f4e5758a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf188cf3b3e6057d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7482882596dc9266;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h482a6486a3bf2d7f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa22d17f0b26fc45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6155f133fd84b83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f53ccdb05683208;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3451068debf7f03f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1a1957d8cd5407f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58b39ded98b16c05;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4b996cdd91e0862;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45c48c7ba7791d65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h283662b7f2088181;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74f603e00152c5c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd495ac6275e5bc12;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7664dcdf4b36191;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb78376d2c0825b54;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd72f5929412803e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2dd8bc9f51fa231;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59df58feaa6f617;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf061f6980770f201;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cc107c02c5d4c91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba58aa73b96d8a08;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h575ffc513d8cbdf8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc1447c85f39b473;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3eaeeed6f2d02e50;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3855ad0355806b49;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9d7e97ce8577887;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed81289b093c75a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcac1451e30c18754;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6be512e3fb377016;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f9dacd14805d9bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he1950467a668eb5e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc8c156ccdb8ce4f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h594e512b70e00b4a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb81d2835037252e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h220a470a2b5f0b87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcebe7cfa11229ec3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h971bdb3546d8e8bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c8f06fa75e33fb5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d398ad5d6b077fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63b5c81eb797d30;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45c8faa3ba4fd74b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f496c90aab26c81;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8993ea87e60dd574;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfdb558a9363ab55a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc44d4d7724c9128c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29a255f0c21d1f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he38cbf0d3b92e982;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16446d5aa5687bd0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75dfee2233243dc2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5191f15e948ac738;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h127970e7f8798d4c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22d6c49201653d3d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc76f1f1a53c08dcf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa06d88c422e6ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9dabbe096d7dd69c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf769cb0c5ba3fd22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a8d97669ed71c7f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6731d1d7d9f6a1ec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45e70da578eeb485;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48f97b9aab8a1e22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27a76bab98947f59;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5407b04546bf15;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f0f96256842216;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21ac7c446cb2ed3d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb728f51553cf8bee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0b7ea525a7fa580;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc2de7ba7985ca9a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h873e8271c94b4c46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc06b63be399c07bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd93ce9115b0dc333;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6f05ea148b061e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87a821843aead93a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b598d657b612ac5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h410f8552051ec040;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h525d73e050c367d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5a8570bcbc4cadb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73aa21ed8d25f22b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cb60447f39da570;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6808910529a91a61;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3d3fc271bd0dbcf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7511b464477e53e7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0de1aa0ca9160b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h953948670dd6d7f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2585fd08dff7b824;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7ff485440e01b6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66116b879c694b3e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h376524e4e5dc79d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34c5c5acf089890d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7aa8f8800a2ebfff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h307966b9f51c13c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf72ea884a65ac827;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he44e8d0b0ca61c6c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33623e4f435fe8f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6c425e897e6156;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44d048243cf1bb83;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83e416cbcc15da66;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb2d6e9aebc36e65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbeba94e5a252a800;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h555371a5acd68a8d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29ccb81c06f54069;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc59760fe855c51dc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha79adc70e02f589b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4016afd3f4217a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a8c57fcc7a1ebd7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h430c4c227e9e6f4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ce8c91210d8691b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9ee6cd89d885a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29957d5275041fd4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h179b139b9bbefd14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59c5162af0a993a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h893e45fa721eac13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7528d9425057a059;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8776b22409dc359c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23359a0ae1cfc696;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb79cf3e4c97d5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73ad489558b2b726;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1836111f4e811e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c92d6323aef79ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c43ee61700fff2a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h325216513b6b8733;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b7f53644e4a2b6c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52885a19e06a71a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c755240ca2684e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1961034068b4856b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf53e383b0404dd91;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d788376511a7c17;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2fb5b664a97be59a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5c3285a5b1daaae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d1233759d20cc2f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec2b36fa76b20cff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he234fa5758da6d56;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b531259ea60edb7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5be3076b00b86968;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h24a1af0632e9baed;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h453c00740e8335bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29bddf3baa482ec2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he649fc7f03d85982;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd854d61c97dfa94d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he703ce916d7e63a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h634ebade57c69589;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a12e943a33d2a4d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65a4266cc411c107;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ff3f0fd581148cb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6992a99043965ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a3ce848a0f06f92;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a7aa6b9d550126;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he17c3affca0f8c2a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97721d215115777f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc69a0a7f16f51649;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4a657750f05c02a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc70d4bb03134a494;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha41fdf76fe43fa4b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b8a97c4c0cdcaf6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h404328dc0db3e461;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha64607f294c3a6e7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf74425e85beb404d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe0d1cc00d5c3d6d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf77b9725471e8cce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f7dee02eaaad1e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78beedc37553f776;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61e3c1bff1b21bf6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d500dc59420dcc1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he5fcefcaabe4afbc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7665e9eecdae2811;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8101a0509874697c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h823b75835b6ab263;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ef53703d77a80aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3e3b15716092050;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7484e85fd279f1f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b4180f2e0e15b34;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3799b550f3e8179;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f2b4fb3ae431044;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5067ae50de45b46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46eb12dbaea6dd67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha97be550a9502975;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3130b926b7b1a92;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he24085b6cddf7a3f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb74bf110e4e88bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40561ed595ed11f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d30bdaf588defcd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9abf95e9e6fecc5f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f77a8366b935287;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61df6f269d2b9f13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc03586599eeafe36;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h629c9b30ebc7cb8f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf7f27f0108525ff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h215c1e9a76c85151;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he704670228b6238f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h424ffb34ad3ff7d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h69325b2c77c7661;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5be79ddef094d5f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5dae72964b9b2563;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73490599719bb8c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacfc882179b70914;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had0ccd12d86ad756;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a6ca332612affe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f93825f4253b3a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2eaea9b6b762e73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h14e7b53b8cec7158;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ef80807eaaa4203;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ba4cf76c9deb786;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h902f632033656039;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4358d4fd66a56ddd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41a9d6085e9e9935;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec8aa56fc46ac9cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h680442a99eb1678b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8f253005afa9467;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46e71df5e72f33f3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7421968ea8cc55c1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd17d414786c0bcbb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c830300a7220fe7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d94e085ca0d8377;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb73c7a3f39c685a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heeed9cc8f1842eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haabcabfca9f246b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2755bb6c50050a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdb64c0fc34de126;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d6b7d62ce67a579;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89b183e1b69df535;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h636d475ca72e777c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9939df0f012fe80;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b950dab14303e24;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd3bf25c78aef8d5e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61c8c4fc70a167fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34e70779629c3749;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he338e9931e8fa6bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc143606639ef8b9b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb62c21fb45d9385c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25f5d9c8ac2fde9f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d98f32301e2fd47;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4bea968953a8d17;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcc66345132b4f19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cab94cd1bbc834c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha12c9399bed09241;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7d883d2d9e6d332;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51c0fb4dc5d04462;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a414a1cd29f8d7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf72afd349e48b57;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h678b71ae9c1df505;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95b7ab0ad5f04ff8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h867f5cfd500fe52e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56933531e37ca1d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbecd27ca95e398ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha73c36543e5e594f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b7a535313fc208e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa917ab13f0353db;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h735c1656e37c9d10;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0f132ddc19d7cf2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha34eda39982da9e6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he6453f7e20427af2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d7a2b0868cd6013;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b730d2637347450;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45701e21b0a203e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0e10e40a677d6c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3279796d0617d40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef7e883ab0e272d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6ff0308ea5c25e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h114de05a0fb26aeb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha62816977fefdd98;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha405ce3a27bb6ade;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha17c0c9d66140c62;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h510dff07592b8b22;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdba22ecedfb8cee5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e2f3b0b138b8dba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3cf0239425f868b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4e20f080903de64;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h673ac15ab5ad6f34;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfdb241aae5c2552;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1073d1f817516e1f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb428f3babfee4c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc60992b578ceb40f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1207f0e623aa80c7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdaf02224a32738d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1b71372a4f20dff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb064b1c7769916b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb55ed89403e235cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc524ff93458e3a7d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd810888cffe96cca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha53484f04e72bc70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a9c166712ce325d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac6e8bc385c77c87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he553218fef9685f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a1b1b1aa9f2a181;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef9ce8f8918899a0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27f8087cb84a55e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7edbbd717e0aa1bc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52a934b9ceafb833;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9c5d09f2a2462a75;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38beef0118b957cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c1910f9d963facd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa2280a6bb98314f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10613dfdfdb35faf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he74deb242714d59e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h653a4de797344c7c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h143d675d058c6d6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61073dac74eb4abb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fcc6c0ed6a2e409;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33d08c8422d7a635;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f93f52cf2589635;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb019c62dcc529be8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ba8d83c2d7ad12b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf702e7cf7e01f90c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27e531f74576350a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70c2999446a23184;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e5477d7efb53b9d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cf42472e7893c42;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha84b328edd35b0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a449c8a0918b109;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ddacfce7c38f825;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h137951aff3ee4aa1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63666ecc3cf7d26c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e6c8881804352c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb17819aa672fe9f8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5e3709746a2e950;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4072aa020a7150c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bdcf86242f76d88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6cd7caef5c41cd4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hafd4716ed901b038;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd869e7c5c4acd18;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac067b865c7060af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h939f6db4255211d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfef5b9206ce160c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb4c66173fab532a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77965d349dfbca43;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6c320f84f586136;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15e1f5e40665b5f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd16197e9af90fbfc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7343992e10863a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdef89079bc50da46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30105af66a0ae96f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b0d2720e9b5f7f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b91333ab7d56aff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha30da1f27d46460e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ff00b11c7f15e1e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbea1ba32102f644e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3914d3dfbb293cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc8513b4b7b0fc87;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51aa3dc648d2bf2d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66bcfc796a12335f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde21522d5a3fd19d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4bac62ae8aa7848;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4bb0ee1eeb703284;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95bc89c20125112e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h568ff4e004682a53;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e63dce751cf9b9c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5860ec9126d69457;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92ba6367e5193852;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4cdf0597aebb1cdf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb22cf0f2a80d41c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heebf257850a4f9d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca93cacf38a70853;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h247305e881c1c3a6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff4bd8c5501941a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc004f456a880975a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70a85cddda06be17;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ff3a2e3563bd26d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d32481369eadb6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8249e45aafd2348d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h557d63a073edd1a7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40fbeaa43ca37e45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b4d381c98504669;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9dbc955f9eba3af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc143da74b5097b75;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f0f61f9fd3aa6ae;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d449520ee561d9a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba376c39ffd5bd85;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8559cc10df44b7a2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce46733eeb76af21;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3afa147a77238e01;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha466866a3c576ba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7310ac9d0936876b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5c7d45111037efa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9e465d266959f8d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h786dbaf15ca88e89;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73f45630317efbe3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a1ac8c7079eb8fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc118d2a4938601c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65a991aa6d7fc960;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62ce68ee0a1904ee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h370dc8a2740d7dcc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h127c90f417e62759;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h613bb217045b758e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h378964fb67bbb363;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42dd59e068894a12;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9d51e186a1ed8c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hafbccdcf98cba575;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27c5dca3d26de4d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d60bd7fe3bfa47d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33f349b470a7de02;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h621be57784f7fc6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h232eb77bddddef00;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacbc1c00e4530936;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9f49ffdeb98bb68;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc66c23c204db20b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb21723007ac5a429;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h896d67db317fe9ca;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd37961e40d3bf503;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha12f400820ea2495;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfea68056a094c37;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfee9edb29c8cf578;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc175c19fc84c78e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d98c9ff1159e6ef;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h944f9d662455ca98;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h410c82ab75b108d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1bb0bbb70f896e6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2ff6ef100e39efc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41d004c8572c92cd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h10430cf2194cbe4c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0b60524062b73f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ef3e8629625fb80;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e0ed90961e1c7c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb59318a5a30ce19;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef1e28ccb4eac4a9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf77e453e701725eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb13796cb50eb9df9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h759eaf59059816f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f483b1d506c9726;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h764219d577c45f62;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60516ed07963bf0c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93b8c57a06a3b3d8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1cac3d69c90808b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6eaedfbb65457c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e1fd1051b88c230;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1f1c1fff3efc96f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haaf743390d805127;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf55c153e91c189;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ff2d5f0286c8506;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6cd5458b7c45e4b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a90170f8f022cb1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffde546f64a103f4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18e297fb6052b1e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35fcf77d154508c6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23cebb4677111cff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf01264b80482782d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c14c7d1e801875b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc8454fb1f928b5b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9aa98eaeb9177c96;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc358ec1aad252b3b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1442eb5f1e562df;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h636b3ca0d567c3f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h83aa8c8256fcd274;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb0bb7946d51a259;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8ff74b3e54a9a6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1dfd763e222ae08a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa16e7704fb24c86;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd21dd1b37b0eb090;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he38b64e1dc3f4a4a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a42df268c32dc27;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9eea57f3b47cf00d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59e93af25c034eee;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4da92a1b857a2d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c7cfee229695c2e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf469355fe5f8bfe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he1ffc4a9a950ea99;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf98c20b1e575ba8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc42e1e519b1f23;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0c23c73c9b6882b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb15a242d285fbb6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a4b5ab220432466;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20bf893247124f27;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbd8c37883c313f2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5f150a9fad45c26;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7466ba817104e68b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ed60fe891f4c714;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha59f91bc125d999b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha47cc3844024e71e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a5db0281aa6b420;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9025ccd21fcab46c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8aa47e5a7e429136;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he65f944ad0ecdcda;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9010380da142275;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d42b24f111cc340;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h506498113931944f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54a244002c537311;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1584d32e143b9f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e3a4129a76bb194;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e31f82eb3a22782;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2c93471d23e6f4a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87f5f5339ecf3ad8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he625b5344a2cb806;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9db3b244b3c4f8a7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb838d1a6e0442fba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba2c30a3c7df43e4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e65fe0dab9bcb71;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfcae0d209359b3e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d2a96e8a5256eff;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5967c6fb01e93658;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbca4034dac64103;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6701d3d60d8fbe1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72cf732184b05337;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2be87d7ddd0edd5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9cfb0bce38d9f836;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd442b498b3088e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hceacb15f1cebbb3e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73aa512043cf6402;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd377d66890b4d99f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6663d820b0e45761;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f5ac08a725f1909;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee251075042b3667;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h118d9a0e870b9cbc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcb111200ccdf245a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca60a5656fa0f7fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d7b1a3ab4a64865;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23198b5d05d26d74;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h693ad68e6fc92ffa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc7496159b4dedfd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h952c923718cf8da6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb524470d07e26e14;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1730f34b87e3e36d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8840ccaecda6544;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44a9991c80a84bd8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he598c2771b01b20f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c60296e50bb7cdd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ef863c3c5b51960;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8dac31be2a891914;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h376b5e81f9b2e404;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5e62c823541c40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92f335d4b1264fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hac4406cc86cf7e7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1abee21b132101fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcdc0eb92aa64bf98;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5856ca0e398997f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he1a294980e3dfc93;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab3ae92bd7a01e44;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e9d295a16877f9a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb197ccd5bcec36c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h697f43b745f51790;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h13d8e89868c3e89d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1a375d4bf0c05a27;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ce193d8e0698a40;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8342e939e8b25b5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he06b588ac1062abe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h209f356079df19d2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h302b6681019a80fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84d45dfb171372da;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34415f658c516033;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha566d4a4a20984c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hced0b09447b82eb2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef681bae9728383;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf1e7633dde68081;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae76d0831fd548fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb786155d7085221e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76f0c169cc456665;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59c2a950562bc54d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8306719ec3b515a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e4bf6b48b5300d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1755e21e09cea1ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f5a02bbe0efd01f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2c5117fe76b4ad4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e424cef1b48802c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3fa156a9c31e3d9d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f13655cd66b612c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadceb4a123cfcc57;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e23a621cf8e9ef2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91d2b6b71c0c276f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e3a41fd288bd2f3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8de4663696f02a0b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86c920aa8a19fdbf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9a6c6b9e171f419;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61a6f989a570d501;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23775f78b746b199;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd693b625f3da4cf5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6a4a7bfcdc62bd7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a0cb23ff552d121;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0385ac03bda88a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb94a7a00c3518690;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h972ab87f9fc745;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha6540bc7fff3b85b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf25b5c336d69f665;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a9b42d56f8cdd45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e8802958d45a49b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h554c9754135feb9e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h884f2dc7b5f8d320;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h287004a775589694;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf738533a3a84bffe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57be65128fb80542;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc03af7c9a68eb868;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc294bab2d8783690;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h145408ca814c4cb4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha744899de9dd694f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85319684f45f15c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf6a9f3c65ac71a7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43894119a931960d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0f247c71b3d37aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc0e05cb9f16a913b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h234f734d6c4d5e94;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b48098c95e87f33;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79d751de2c359d70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec162bf737ec0eb1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e71f995d991537e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf4d34c4655ef427;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbfc2187d363f026;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f890aba9a04b1f5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75adaf7eab6436f0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef5eb2db6ea023c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5812535edee89485;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c299a5a568ea54a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b42ef4db4a9936d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7bf7a9fb54256d6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9cdf81915299fd0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha98b55a66023bdfd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc8b09902300f575;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h959f91893f9ef286;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b2abf67cd5e4fa3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2363db3f73512f1b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16852a9d1d3cadec;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63ae47fcbce266ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd389bfa7dc34d32c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h424c29b8d6026b61;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94ac4c1baf9ec345;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb19cb9150459cab0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc75672843fd62c2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2bc1694f8007ab;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95dfe906b88fa7e8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72900f8cf7886d52;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb86e6842714bacf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e211227f10c3e36;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb435de1bf094b4f7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb06580fd374c40cf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h840925b78d368994;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66b23cbd6bfdf5ce;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3aacaeed5063b71d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f687ddd75d840fd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6515a2daf55b1a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h283a468888798fe5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hba322eb74e6f1788;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e3e54e6f17ba293;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h885f5adb7b3e8abe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8acbba7362492337;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6992e9217cfed4ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6a61c23ca0c26f3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19c8a27e8f133c15;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86d8c9964ad96760;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70c656630ed1a24d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d5ddeaa0d1348b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11846ba3178fd229;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf63e3d6dfc61f13;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h731e8a6eb3a92068;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h396666742a685ba5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38dce88f5f02ef18;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28866f8f87a8954;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc6d6c725c330f23;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f536d4648a46af7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3399a1d0369536a7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he03a9b6654c552e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97f5c07014ef2acd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7e82f7a64585b89;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0bc2e0f8bb4f98e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32e7101835816ad7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha436b6c169009cf3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h837d898aeaba6d7c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7607727208ee0c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ea31c326aad7786;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha113acdc002ec8c8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9cebc017e2923dd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa2862de70b79374;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1719dfa8167128e1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0722a1df66d66de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb69c03ba20b99b02;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21b8d9b91763267d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe6a7ebfad285613;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76d36b1828ab7f6e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed9514997eeeb647;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe07ee32b728b252;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12c318eae767f05c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacd0cb702507d94c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc90e95a0b73d4034;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81a79ff2bac64b45;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbbd0e03e07b59fa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67246172d874858a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ac1a71b26386663;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haae5cf2809b115a1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a5f89ebb2674fe1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h242e4102aa2010b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb47bc18ff11dc359;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf65e1219f2bfaf2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd2311fcdc13f8a90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4461bcc9ad8ab77;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64877e7c0d1ee88d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe8bca71a8c7ae73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5529449f13f25b8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44347b9ff67276b1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2da470f5efadc2de;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2c0fbaee53f21d4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h593af77adb08e468;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbea4196dae25420;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h730d010e6f9550b3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha38685234a3bac7e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ac8cd867ac5bf2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbba7a1ffa0ebe7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7aad2be083d4715;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d258d7edaaf38b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4126bb60fbf32dcb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b6a780906be589;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e6db0236b2e8514;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90a3a33fdb7a7dd6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc10a0c7890153ca6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f958f303647b93c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dc36154ed6336c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54e68e673291108c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1bd6a90eb077534d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3eb1784a75ab165b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf35497478148a74b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha71a30b36d86dc41;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha13524afbe8a9014;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hacaec0769fc034e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7991d08cc42c6bb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee1e0b14c6441c58;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf08e4dbe955baac1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd79c20d2208aee4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde771260857db7c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdee24005f34fc8ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5daa23b3a9c14757;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc19d2cf7f0e71dfb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f10b004686997e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc50dbd3fd2bad9a8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab7eceb793930d46;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e0adf67ffac2e8e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51be32db52b69a5d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf7b869d5b9f5f88;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4da851e24ef5b73d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h12db0f0d323f1a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb59f6f4b9cb2bd2c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51468f8fa4c3c5f6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c0951b03c326085;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha05c4b7b8fb37e4b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59648a7dd81e73e5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h686411b7af615a3a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34f9bedba6373f12;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e6df1f6a46c2d72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h316b671e0cbf85b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35cb8730b79f2a4f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5545233164a31c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h13d535aaec74167b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h114522e1ebabcbc4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11e170ad00e038e7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h693d4e3b61a4f616;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdeb3e767575c5b1d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha77cbf53a8228256;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf68db14fd362032f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h691cf1e514bfe23e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef59f94f8aad2c6b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fdbef9ab3844bb1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h19f02f01fff0cd70;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hed14a571ccc9f44a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9537e81fe2224649;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h97f498606dcd36a5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53b3b5f9b00da79f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a7918c43bb1453;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74e7d7254619119f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h170f72994702a3eb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47e327d50a4a9f26;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f9e6bfdee1199ba;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8da3c87a5b7c644a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68fdae465d3d2d0a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae6a6933798fd1c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55a9c8a3586a430;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94ef7725a802ffd0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h645a9bb805eadd4c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c2b30b1863666c9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c83d118efd6b93;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdba17e308b358ca7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b724a44ca78bc50;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7eda310b173be532;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h635bef8f629db085;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46dec05a10ecaa9e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h788c633e867a8a6c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7f2c854974fa4fb;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf23df9fb44a66ecd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf31b14e18075084;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92800dff5ce1bccc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heccb8184cf5ac5bf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84f9b8cacf0f1df8;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd76b660e6b6714af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fcac0b6047c5108;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ae144986846e410;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4abd73f5e52eaf2b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h174802aa7fc928a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4152fc05e8b98ab6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fd2d40ed37d9313;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8ffd6b2d5bb9105;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80bb2ad754380de5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h900931d19e066237;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4264c9241c07ae72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcacde22ed9b69f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb673bef91ade2748;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2f62720a5cd49f3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd7df14d323f759a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4344e012744528be;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8a6023c090817f1c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4f9cead5263f163;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde6d3da9be7031a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4732ae36e1993fd1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f30bc7a3a50321f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44c05b1f7461ecb4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6594e3ff35e065aa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49df53dfa94e21b2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe3cb3def393eeaa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d355d06bfe3e2a7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd09b62c27c26c437;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1582c5a7efdfdac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc54a6ec814dbe07c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5011f778bf8060bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfee2b6b32092d009;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ed32f7db3bde099;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h923bf8f110da6027;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c559c86ab6ca4d1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f26fbbe2b1b2bdd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9903824e2d5994fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73d41d411a545e5e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he21ab85ffdee9bf2;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h863ffc468ef4048c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc684560c0583391;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h764a59fe2aa7960;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11f7c147bd871bfa;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98be0d921aec8192;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h315d4130bbf7fbd0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5414915b50ec0cfd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a55d48cf7dfd1c0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h726db6994b40f871;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb053a9396eb9136e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3a60f8085ea109a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15f3bc1dc2b2a7ea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0a05683b233bc50;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbfa09ba9294907;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbbd2de9aef8a853c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72d3e3612e2e3676;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf50341dd69462d5e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88801011222563bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3116feaf9831abe4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42cb159880c1126f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf284ceb96ebcfe9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63a52d8558803811;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h393359a28122d1c5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heab548bb27c35544;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f161a619ae3a2a4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15b8a0989b6613a3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62cd8972875c1f31;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3b2f37b21806895;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e7eae31b1f1ba6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf40c1a5de169a05c;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cabb3fef67b46fc;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd608fb894d6e147;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec76077de5cbd374;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87ef8d56b4d2ef38;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5e1c838553992b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdbb27743b559f0d6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27f0181e660bb46f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcdd5fe7e47a5858;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68d97f55d2fc66e9;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h226553c8cb706df3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a3a118d2134b08a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h703f4d4662a4a552;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h13d6b8c1d601d6b6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd077d4cd0d1c9e90;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef995e3725527b5e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fe067535ab4ddf3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2897688db4d62747;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b4700e173490082;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h917446e502fe9893;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h153233d8bcb1199d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20a209e7f42cd902;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3bc92abe549181f1;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3899d38a8ed61a6a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h765b7181decb3afd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf73893356e29fd72;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb56ef68f188220e0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fc1b2641489ac57;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1dd5b797274ad7e3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha57d2036b2affdea;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbfc3f70d7e4b1af6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50c95d0d2082f0c3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ad7108edf34a2d3;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c053ef3e9145086;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0e7c4a0cf95896e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99bf50ff17cdacd6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a7afee24d6f4943;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ab040b3e258ef4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f8ff7c2416fdf4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h274ea67377ad1e60;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28e998b21f8792ac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15dcedcf11b188c4;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddea1afca5317f2e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7858f0823f2b8f47;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2fbb6ca67b602a51;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63f790383e9f2a93;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58290782e2321e17;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80a2cfa0b8f07a60;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4cf2d907e76cb51a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4375a8a0695020a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e8732556c25e859;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h528892ed65058a97;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47f81c897fa0e354;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf61f593bd924b6d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h871d518b23769f60;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha7f8bd29ba42b7ad;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a62da5da48638d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3becc16f7154f89b;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a76c5b8db2a8e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9aef8014ac57f67;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7078950d59d4a371;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8aedf47ec5b48566;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h663309b9de19bf7e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0006bc6a46373fe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f3eeebbf3007eac;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc0917d61d8362bd;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66cc235d723b0615;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h607f02cf171580af;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33837306e293a016;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e18cb33f7b18063;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72f6c5696f349bdf;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdf6d67309e4e3c65;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94761b2d0a29932d;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h713f1e4b4770ff4e;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ba1ccba1a44eafe;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6f0bef4bba67ac6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d2598b902fe8c12;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4573741249dfbae6;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35f06ae00ba04f6f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h462858ad18f23a1f;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he8d10a9ab78303b7;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ad6edf46e8f07d5;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77a395b43b4df1b0;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb48c7e90cb4a9081;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h11ddf956ed855b73;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d5b8db04046190;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ee3ed9d2fbc343a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc852ba668234f95;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9054346bfcf8434a;
        #1
        {src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb871e1b5c8e3bbc4;
        #1
        $finish();
    end
endmodule
