module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    compressor_CLA16_32 compressor_CLA16_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35));
    initial begin
        src0 <= 16'h0;
        src1 <= 16'h0;
        src2 <= 16'h0;
        src3 <= 16'h0;
        src4 <= 16'h0;
        src5 <= 16'h0;
        src6 <= 16'h0;
        src7 <= 16'h0;
        src8 <= 16'h0;
        src9 <= 16'h0;
        src10 <= 16'h0;
        src11 <= 16'h0;
        src12 <= 16'h0;
        src13 <= 16'h0;
        src14 <= 16'h0;
        src15 <= 16'h0;
        src16 <= 16'h0;
        src17 <= 16'h0;
        src18 <= 16'h0;
        src19 <= 16'h0;
        src20 <= 16'h0;
        src21 <= 16'h0;
        src22 <= 16'h0;
        src23 <= 16'h0;
        src24 <= 16'h0;
        src25 <= 16'h0;
        src26 <= 16'h0;
        src27 <= 16'h0;
        src28 <= 16'h0;
        src29 <= 16'h0;
        src30 <= 16'h0;
        src31 <= 16'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA16_32(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    input [15:0]src16,
    input [15:0]src17,
    input [15:0]src18,
    input [15:0]src19,
    input [15:0]src20,
    input [15:0]src21,
    input [15:0]src22,
    input [15:0]src23,
    input [15:0]src24,
    input [15:0]src25,
    input [15:0]src26,
    input [15:0]src27,
    input [15:0]src28,
    input [15:0]src29,
    input [15:0]src30,
    input [15:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [0:0] comp_out3;
    wire [0:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [0:0] comp_out34;
    wire [1:0] comp_out35;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out35[1], 1'h0, comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], 1'h0, 1'h0, 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [15:0] src0,
      input wire [15:0] src1,
      input wire [15:0] src2,
      input wire [15:0] src3,
      input wire [15:0] src4,
      input wire [15:0] src5,
      input wire [15:0] src6,
      input wire [15:0] src7,
      input wire [15:0] src8,
      input wire [15:0] src9,
      input wire [15:0] src10,
      input wire [15:0] src11,
      input wire [15:0] src12,
      input wire [15:0] src13,
      input wire [15:0] src14,
      input wire [15:0] src15,
      input wire [15:0] src16,
      input wire [15:0] src17,
      input wire [15:0] src18,
      input wire [15:0] src19,
      input wire [15:0] src20,
      input wire [15:0] src21,
      input wire [15:0] src22,
      input wire [15:0] src23,
      input wire [15:0] src24,
      input wire [15:0] src25,
      input wire [15:0] src26,
      input wire [15:0] src27,
      input wire [15:0] src28,
      input wire [15:0] src29,
      input wire [15:0] src30,
      input wire [15:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [0:0] dst3,
      output wire [0:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [0:0] dst34,
      output wire [1:0] dst35);

   wire [15:0] stage0_0;
   wire [15:0] stage0_1;
   wire [15:0] stage0_2;
   wire [15:0] stage0_3;
   wire [15:0] stage0_4;
   wire [15:0] stage0_5;
   wire [15:0] stage0_6;
   wire [15:0] stage0_7;
   wire [15:0] stage0_8;
   wire [15:0] stage0_9;
   wire [15:0] stage0_10;
   wire [15:0] stage0_11;
   wire [15:0] stage0_12;
   wire [15:0] stage0_13;
   wire [15:0] stage0_14;
   wire [15:0] stage0_15;
   wire [15:0] stage0_16;
   wire [15:0] stage0_17;
   wire [15:0] stage0_18;
   wire [15:0] stage0_19;
   wire [15:0] stage0_20;
   wire [15:0] stage0_21;
   wire [15:0] stage0_22;
   wire [15:0] stage0_23;
   wire [15:0] stage0_24;
   wire [15:0] stage0_25;
   wire [15:0] stage0_26;
   wire [15:0] stage0_27;
   wire [15:0] stage0_28;
   wire [15:0] stage0_29;
   wire [15:0] stage0_30;
   wire [15:0] stage0_31;
   wire [6:0] stage1_0;
   wire [4:0] stage1_1;
   wire [8:0] stage1_2;
   wire [5:0] stage1_3;
   wire [5:0] stage1_4;
   wire [8:0] stage1_5;
   wire [10:0] stage1_6;
   wire [6:0] stage1_7;
   wire [5:0] stage1_8;
   wire [8:0] stage1_9;
   wire [5:0] stage1_10;
   wire [5:0] stage1_11;
   wire [10:0] stage1_12;
   wire [6:0] stage1_13;
   wire [6:0] stage1_14;
   wire [6:0] stage1_15;
   wire [9:0] stage1_16;
   wire [12:0] stage1_17;
   wire [5:0] stage1_18;
   wire [5:0] stage1_19;
   wire [5:0] stage1_20;
   wire [5:0] stage1_21;
   wire [8:0] stage1_22;
   wire [6:0] stage1_23;
   wire [6:0] stage1_24;
   wire [7:0] stage1_25;
   wire [10:0] stage1_26;
   wire [5:0] stage1_27;
   wire [7:0] stage1_28;
   wire [5:0] stage1_29;
   wire [11:0] stage1_30;
   wire [8:0] stage1_31;
   wire [2:0] stage1_32;
   wire [1:0] stage1_33;
   wire [0:0] stage1_34;
   wire [1:0] stage2_0;
   wire [1:0] stage2_1;
   wire [4:0] stage2_2;
   wire [1:0] stage2_3;
   wire [2:0] stage2_4;
   wire [5:0] stage2_5;
   wire [2:0] stage2_6;
   wire [2:0] stage2_7;
   wire [2:0] stage2_8;
   wire [5:0] stage2_9;
   wire [2:0] stage2_10;
   wire [1:0] stage2_11;
   wire [6:0] stage2_12;
   wire [3:0] stage2_13;
   wire [2:0] stage2_14;
   wire [1:0] stage2_15;
   wire [6:0] stage2_16;
   wire [4:0] stage2_17;
   wire [2:0] stage2_18;
   wire [5:0] stage2_19;
   wire [2:0] stage2_20;
   wire [2:0] stage2_21;
   wire [3:0] stage2_22;
   wire [1:0] stage2_23;
   wire [2:0] stage2_24;
   wire [6:0] stage2_25;
   wire [5:0] stage2_26;
   wire [1:0] stage2_27;
   wire [5:0] stage2_28;
   wire [4:0] stage2_29;
   wire [1:0] stage2_30;
   wire [5:0] stage2_31;
   wire [2:0] stage2_32;
   wire [1:0] stage2_33;
   wire [0:0] stage2_34;
   wire [0:0] stage2_35;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [0:0] stage3_2;
   wire [0:0] stage3_3;
   wire [0:0] stage3_4;
   wire [1:0] stage3_5;
   wire [1:0] stage3_6;
   wire [1:0] stage3_7;
   wire [1:0] stage3_8;
   wire [1:0] stage3_9;
   wire [1:0] stage3_10;
   wire [1:0] stage3_11;
   wire [1:0] stage3_12;
   wire [1:0] stage3_13;
   wire [1:0] stage3_14;
   wire [1:0] stage3_15;
   wire [1:0] stage3_16;
   wire [1:0] stage3_17;
   wire [1:0] stage3_18;
   wire [1:0] stage3_19;
   wire [1:0] stage3_20;
   wire [1:0] stage3_21;
   wire [1:0] stage3_22;
   wire [1:0] stage3_23;
   wire [1:0] stage3_24;
   wire [1:0] stage3_25;
   wire [1:0] stage3_26;
   wire [1:0] stage3_27;
   wire [1:0] stage3_28;
   wire [1:0] stage3_29;
   wire [1:0] stage3_30;
   wire [1:0] stage3_31;
   wire [1:0] stage3_32;
   wire [1:0] stage3_33;
   wire [0:0] stage3_34;
   wire [1:0] stage3_35;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage3_0;
   assign dst1 = stage3_1;
   assign dst2 = stage3_2;
   assign dst3 = stage3_3;
   assign dst4 = stage3_4;
   assign dst5 = stage3_5;
   assign dst6 = stage3_6;
   assign dst7 = stage3_7;
   assign dst8 = stage3_8;
   assign dst9 = stage3_9;
   assign dst10 = stage3_10;
   assign dst11 = stage3_11;
   assign dst12 = stage3_12;
   assign dst13 = stage3_13;
   assign dst14 = stage3_14;
   assign dst15 = stage3_15;
   assign dst16 = stage3_16;
   assign dst17 = stage3_17;
   assign dst18 = stage3_18;
   assign dst19 = stage3_19;
   assign dst20 = stage3_20;
   assign dst21 = stage3_21;
   assign dst22 = stage3_22;
   assign dst23 = stage3_23;
   assign dst24 = stage3_24;
   assign dst25 = stage3_25;
   assign dst26 = stage3_26;
   assign dst27 = stage3_27;
   assign dst28 = stage3_28;
   assign dst29 = stage3_29;
   assign dst30 = stage3_30;
   assign dst31 = stage3_31;
   assign dst32 = stage3_32;
   assign dst33 = stage3_33;
   assign dst34 = stage3_34;
   assign dst35 = stage3_35;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10]},
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage1_4[0],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[1],stage1_3[2],stage1_2[2],stage1_1[2]}
   );
   gpc606_5 gpc3 (
      {stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[2],stage1_3[3],stage1_2[3],stage1_1[3]}
   );
   gpc615_5 gpc4 (
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage0_3[12]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[2],stage1_4[3],stage1_3[4],stage1_2[4]}
   );
   gpc1343_5 gpc5 (
      {stage0_3[13], stage0_3[14], stage0_3[15]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9]},
      {stage0_5[0], stage0_5[1], stage0_5[2]},
      {stage0_6[0]},
      {stage1_7[0],stage1_6[1],stage1_5[3],stage1_4[4],stage1_3[5]}
   );
   gpc1406_5 gpc6 (
      {stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15]},
      {stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4]},
      {stage0_7[0]},
      {stage1_8[0],stage1_7[1],stage1_6[2],stage1_5[4],stage1_4[5]}
   );
   gpc606_5 gpc7 (
      {stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7], stage0_5[8]},
      {stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6]},
      {stage1_9[0],stage1_8[1],stage1_7[2],stage1_6[3],stage1_5[5]}
   );
   gpc615_5 gpc8 (
      {stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13]},
      {stage0_6[5]},
      {stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11], stage0_7[12]},
      {stage1_9[1],stage1_8[2],stage1_7[3],stage1_6[4],stage1_5[6]}
   );
   gpc615_5 gpc9 (
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10]},
      {stage0_7[13]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[2],stage1_8[3],stage1_7[4],stage1_6[5]}
   );
   gpc615_5 gpc10 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10]},
      {stage0_9[0]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[1],stage1_9[3],stage1_8[4]}
   );
   gpc615_5 gpc11 (
      {stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage0_9[1]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[2],stage1_9[4],stage1_8[5]}
   );
   gpc606_5 gpc12 (
      {stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[2],stage1_11[2],stage1_10[3],stage1_9[5]}
   );
   gpc606_5 gpc13 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[3],stage1_11[3],stage1_10[4],stage1_9[6]}
   );
   gpc615_5 gpc14 (
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], 1'b0},
      {stage0_11[12]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[2],stage1_12[4],stage1_11[4],stage1_10[5]}
   );
   gpc615_5 gpc15 (
      {stage0_11[13], stage0_11[14], stage0_11[15], 1'b0, 1'b0},
      {stage0_12[6]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[1],stage1_13[3],stage1_12[5],stage1_11[5]}
   );
   gpc1343_5 gpc16 (
      {stage0_12[7], stage0_12[8], stage0_12[9]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9]},
      {stage0_14[0], stage0_14[1], stage0_14[2]},
      {stage0_15[0]},
      {stage1_16[0],stage1_15[1],stage1_14[2],stage1_13[4],stage1_12[6]}
   );
   gpc623_5 gpc17 (
      {stage0_12[10], stage0_12[11], stage0_12[12]},
      {stage0_13[10], stage0_13[11]},
      {stage0_14[3], stage0_14[4], stage0_14[5], stage0_14[6], stage0_14[7], stage0_14[8]},
      {stage1_16[1],stage1_15[2],stage1_14[3],stage1_13[5],stage1_12[7]}
   );
   gpc615_5 gpc18 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], 1'b0},
      {stage0_14[9]},
      {stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5], stage0_15[6]},
      {stage1_17[0],stage1_16[2],stage1_15[3],stage1_14[4],stage1_13[6]}
   );
   gpc1343_5 gpc19 (
      {stage0_14[10], stage0_14[11], stage0_14[12]},
      {stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10]},
      {stage0_16[0], stage0_16[1], stage0_16[2]},
      {stage0_17[0]},
      {stage1_18[0],stage1_17[1],stage1_16[3],stage1_15[4],stage1_14[5]}
   );
   gpc1343_5 gpc20 (
      {stage0_14[13], stage0_14[14], stage0_14[15]},
      {stage0_15[11], stage0_15[12], stage0_15[13], stage0_15[14]},
      {stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage0_17[1]},
      {stage1_18[1],stage1_17[2],stage1_16[4],stage1_15[5],stage1_14[6]}
   );
   gpc606_5 gpc21 (
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[0],stage1_18[2],stage1_17[3],stage1_16[5]}
   );
   gpc606_5 gpc22 (
      {stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5], stage0_17[6], stage0_17[7]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[1],stage1_19[1],stage1_18[3],stage1_17[4]}
   );
   gpc615_5 gpc23 (
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10]},
      {stage0_19[6]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[1],stage1_20[2],stage1_19[2],stage1_18[4]}
   );
   gpc615_5 gpc24 (
      {stage0_18[11], stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15]},
      {stage0_19[7]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[2],stage1_20[3],stage1_19[3],stage1_18[5]}
   );
   gpc1343_5 gpc25 (
      {stage0_19[8], stage0_19[9], stage0_19[10]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15]},
      {stage0_21[0], stage0_21[1], stage0_21[2]},
      {stage0_22[0]},
      {stage1_23[0],stage1_22[2],stage1_21[3],stage1_20[4],stage1_19[4]}
   );
   gpc615_5 gpc26 (
      {stage0_19[11], stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15]},
      {1'b0},
      {stage0_21[3], stage0_21[4], stage0_21[5], stage0_21[6], stage0_21[7], stage0_21[8]},
      {stage1_23[1],stage1_22[3],stage1_21[4],stage1_20[5],stage1_19[5]}
   );
   gpc207_4 gpc27 (
      {stage0_21[9], stage0_21[10], stage0_21[11], stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15]},
      {stage0_23[0], stage0_23[1]},
      {stage1_24[0],stage1_23[2],stage1_22[4],stage1_21[5]}
   );
   gpc2135_5 gpc28 (
      {stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage0_23[2], stage0_23[3], stage0_23[4]},
      {stage0_24[0]},
      {stage0_25[0], stage0_25[1]},
      {stage1_26[0],stage1_25[0],stage1_24[1],stage1_23[3],stage1_22[5]}
   );
   gpc1163_5 gpc29 (
      {stage0_22[6], stage0_22[7], stage0_22[8]},
      {stage0_23[5], stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10]},
      {stage0_24[1]},
      {stage0_25[2]},
      {stage1_26[1],stage1_25[1],stage1_24[2],stage1_23[4],stage1_22[6]}
   );
   gpc606_5 gpc30 (
      {stage0_22[9], stage0_22[10], stage0_22[11], stage0_22[12], stage0_22[13], stage0_22[14]},
      {stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5], stage0_24[6], stage0_24[7]},
      {stage1_26[2],stage1_25[2],stage1_24[3],stage1_23[5],stage1_22[7]}
   );
   gpc615_5 gpc31 (
      {stage0_23[11], stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15]},
      {stage0_24[8]},
      {stage0_25[3], stage0_25[4], stage0_25[5], stage0_25[6], stage0_25[7], stage0_25[8]},
      {stage1_27[0],stage1_26[3],stage1_25[3],stage1_24[4],stage1_23[6]}
   );
   gpc606_5 gpc32 (
      {stage0_24[9], stage0_24[10], stage0_24[11], stage0_24[12], stage0_24[13], stage0_24[14]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[1],stage1_26[4],stage1_25[4],stage1_24[5]}
   );
   gpc1415_5 gpc33 (
      {stage0_25[9], stage0_25[10], stage0_25[11], stage0_25[12], stage0_25[13]},
      {stage0_26[6]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3]},
      {stage0_28[0]},
      {stage1_29[0],stage1_28[1],stage1_27[2],stage1_26[5],stage1_25[5]}
   );
   gpc615_5 gpc34 (
      {stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage0_27[4]},
      {stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5], stage0_28[6]},
      {stage1_30[0],stage1_29[1],stage1_28[2],stage1_27[3],stage1_26[6]}
   );
   gpc606_5 gpc35 (
      {stage0_27[5], stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[1],stage1_29[2],stage1_28[3],stage1_27[4]}
   );
   gpc615_5 gpc36 (
      {stage0_27[11], stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15]},
      {stage0_28[7]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[2],stage1_29[3],stage1_28[4],stage1_27[5]}
   );
   gpc606_5 gpc37 (
      {stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11], stage0_28[12], stage0_28[13]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[2],stage1_30[3],stage1_29[4],stage1_28[5]}
   );
   gpc615_5 gpc38 (
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], 1'b0},
      {stage0_30[6]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[1],stage1_31[3],stage1_30[4],stage1_29[5]}
   );
   gpc1163_5 gpc39 (
      {stage0_30[7], stage0_30[8], stage0_30[9]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {1'b0},
      {1'b0},
      {stage1_34[0],stage1_33[1],stage1_32[2],stage1_31[4],stage1_30[5]}
   );
   gpc1_1 gpc40 (
      {stage0_0[11]},
      {stage1_0[2]}
   );
   gpc1_1 gpc41 (
      {stage0_0[12]},
      {stage1_0[3]}
   );
   gpc1_1 gpc42 (
      {stage0_0[13]},
      {stage1_0[4]}
   );
   gpc1_1 gpc43 (
      {stage0_0[14]},
      {stage1_0[5]}
   );
   gpc1_1 gpc44 (
      {stage0_0[15]},
      {stage1_0[6]}
   );
   gpc1_1 gpc45 (
      {stage0_1[15]},
      {stage1_1[4]}
   );
   gpc1_1 gpc46 (
      {stage0_2[12]},
      {stage1_2[5]}
   );
   gpc1_1 gpc47 (
      {stage0_2[13]},
      {stage1_2[6]}
   );
   gpc1_1 gpc48 (
      {stage0_2[14]},
      {stage1_2[7]}
   );
   gpc1_1 gpc49 (
      {stage0_2[15]},
      {stage1_2[8]}
   );
   gpc1_1 gpc50 (
      {stage0_5[14]},
      {stage1_5[7]}
   );
   gpc1_1 gpc51 (
      {stage0_5[15]},
      {stage1_5[8]}
   );
   gpc1_1 gpc52 (
      {stage0_6[11]},
      {stage1_6[6]}
   );
   gpc1_1 gpc53 (
      {stage0_6[12]},
      {stage1_6[7]}
   );
   gpc1_1 gpc54 (
      {stage0_6[13]},
      {stage1_6[8]}
   );
   gpc1_1 gpc55 (
      {stage0_6[14]},
      {stage1_6[9]}
   );
   gpc1_1 gpc56 (
      {stage0_6[15]},
      {stage1_6[10]}
   );
   gpc1_1 gpc57 (
      {stage0_7[14]},
      {stage1_7[5]}
   );
   gpc1_1 gpc58 (
      {stage0_7[15]},
      {stage1_7[6]}
   );
   gpc1_1 gpc59 (
      {stage0_9[14]},
      {stage1_9[7]}
   );
   gpc1_1 gpc60 (
      {stage0_9[15]},
      {stage1_9[8]}
   );
   gpc1_1 gpc61 (
      {stage0_12[13]},
      {stage1_12[8]}
   );
   gpc1_1 gpc62 (
      {stage0_12[14]},
      {stage1_12[9]}
   );
   gpc1_1 gpc63 (
      {stage0_12[15]},
      {stage1_12[10]}
   );
   gpc1_1 gpc64 (
      {stage0_15[15]},
      {stage1_15[6]}
   );
   gpc1_1 gpc65 (
      {stage0_16[12]},
      {stage1_16[6]}
   );
   gpc1_1 gpc66 (
      {stage0_16[13]},
      {stage1_16[7]}
   );
   gpc1_1 gpc67 (
      {stage0_16[14]},
      {stage1_16[8]}
   );
   gpc1_1 gpc68 (
      {stage0_16[15]},
      {stage1_16[9]}
   );
   gpc1_1 gpc69 (
      {stage0_17[8]},
      {stage1_17[5]}
   );
   gpc1_1 gpc70 (
      {stage0_17[9]},
      {stage1_17[6]}
   );
   gpc1_1 gpc71 (
      {stage0_17[10]},
      {stage1_17[7]}
   );
   gpc1_1 gpc72 (
      {stage0_17[11]},
      {stage1_17[8]}
   );
   gpc1_1 gpc73 (
      {stage0_17[12]},
      {stage1_17[9]}
   );
   gpc1_1 gpc74 (
      {stage0_17[13]},
      {stage1_17[10]}
   );
   gpc1_1 gpc75 (
      {stage0_17[14]},
      {stage1_17[11]}
   );
   gpc1_1 gpc76 (
      {stage0_17[15]},
      {stage1_17[12]}
   );
   gpc1_1 gpc77 (
      {stage0_22[15]},
      {stage1_22[8]}
   );
   gpc1_1 gpc78 (
      {stage0_24[15]},
      {stage1_24[6]}
   );
   gpc1_1 gpc79 (
      {stage0_25[14]},
      {stage1_25[6]}
   );
   gpc1_1 gpc80 (
      {stage0_25[15]},
      {stage1_25[7]}
   );
   gpc1_1 gpc81 (
      {stage0_26[12]},
      {stage1_26[7]}
   );
   gpc1_1 gpc82 (
      {stage0_26[13]},
      {stage1_26[8]}
   );
   gpc1_1 gpc83 (
      {stage0_26[14]},
      {stage1_26[9]}
   );
   gpc1_1 gpc84 (
      {stage0_26[15]},
      {stage1_26[10]}
   );
   gpc1_1 gpc85 (
      {stage0_28[14]},
      {stage1_28[6]}
   );
   gpc1_1 gpc86 (
      {stage0_28[15]},
      {stage1_28[7]}
   );
   gpc1_1 gpc87 (
      {stage0_30[10]},
      {stage1_30[6]}
   );
   gpc1_1 gpc88 (
      {stage0_30[11]},
      {stage1_30[7]}
   );
   gpc1_1 gpc89 (
      {stage0_30[12]},
      {stage1_30[8]}
   );
   gpc1_1 gpc90 (
      {stage0_30[13]},
      {stage1_30[9]}
   );
   gpc1_1 gpc91 (
      {stage0_30[14]},
      {stage1_30[10]}
   );
   gpc1_1 gpc92 (
      {stage0_30[15]},
      {stage1_30[11]}
   );
   gpc1_1 gpc93 (
      {stage0_31[12]},
      {stage1_31[5]}
   );
   gpc1_1 gpc94 (
      {stage0_31[13]},
      {stage1_31[6]}
   );
   gpc1_1 gpc95 (
      {stage0_31[14]},
      {stage1_31[7]}
   );
   gpc1_1 gpc96 (
      {stage0_31[15]},
      {stage1_31[8]}
   );
   gpc606_5 gpc97 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc98 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], 1'b0},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1]}
   );
   gpc606_5 gpc99 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[1],stage2_4[2]}
   );
   gpc606_5 gpc100 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[2]}
   );
   gpc615_5 gpc101 (
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10]},
      {stage1_7[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[2],stage2_7[2],stage2_6[2]}
   );
   gpc606_5 gpc102 (
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[0],stage2_10[1],stage2_9[2]}
   );
   gpc606_5 gpc103 (
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[1],stage2_11[1],stage2_10[2]}
   );
   gpc606_5 gpc104 (
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[0],stage2_14[1],stage2_13[2]}
   );
   gpc117_4 gpc105 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage1_15[6]},
      {stage1_16[0]},
      {stage2_17[1],stage2_16[1],stage2_15[1],stage2_14[2]}
   );
   gpc1163_5 gpc106 (
      {stage1_16[1], stage1_16[2], stage1_16[3]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage1_18[0]},
      {stage1_19[0]},
      {stage2_20[0],stage2_19[0],stage2_18[0],stage2_17[2],stage2_16[2]}
   );
   gpc1163_5 gpc107 (
      {stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage1_18[1]},
      {stage1_19[1]},
      {stage2_20[1],stage2_19[1],stage2_18[1],stage2_17[3],stage2_16[3]}
   );
   gpc615_5 gpc108 (
      {stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5], 1'b0},
      {stage1_19[2]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[2]}
   );
   gpc1163_5 gpc109 (
      {stage1_21[0], stage1_21[1], stage1_21[2]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage1_23[0]},
      {stage1_24[0]},
      {stage2_25[0],stage2_24[0],stage2_23[0],stage2_22[1],stage2_21[1]}
   );
   gpc623_5 gpc110 (
      {stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage1_22[6], stage1_22[7]},
      {stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5], stage1_23[6]},
      {stage2_25[1],stage2_24[1],stage2_23[1],stage2_22[2],stage2_21[2]}
   );
   gpc606_5 gpc111 (
      {stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5], stage1_24[6]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[0],stage2_26[0],stage2_25[2],stage2_24[2]}
   );
   gpc615_5 gpc112 (
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4]},
      {stage1_26[6]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[1],stage2_27[1],stage2_26[1],stage2_25[3]}
   );
   gpc615_5 gpc113 (
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4]},
      {stage1_29[0]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[0],stage2_30[0],stage2_29[1],stage2_28[2]}
   );
   gpc1163_5 gpc114 (
      {stage1_29[1], stage1_29[2], stage1_29[3]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage1_31[0]},
      {stage1_32[0]},
      {stage2_33[0],stage2_32[1],stage2_31[1],stage2_30[1],stage2_29[2]}
   );
   gpc1325_5 gpc115 (
      {stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage1_32[1], stage1_32[2]},
      {stage1_33[0], stage1_33[1], 1'b0},
      {stage1_34[0]},
      {stage2_35[0],stage2_34[0],stage2_33[1],stage2_32[2],stage2_31[2]}
   );
   gpc1_1 gpc116 (
      {stage1_0[6]},
      {stage2_0[1]}
   );
   gpc1_1 gpc117 (
      {stage1_2[6]},
      {stage2_2[2]}
   );
   gpc1_1 gpc118 (
      {stage1_2[7]},
      {stage2_2[3]}
   );
   gpc1_1 gpc119 (
      {stage1_2[8]},
      {stage2_2[4]}
   );
   gpc1_1 gpc120 (
      {stage1_5[6]},
      {stage2_5[3]}
   );
   gpc1_1 gpc121 (
      {stage1_5[7]},
      {stage2_5[4]}
   );
   gpc1_1 gpc122 (
      {stage1_5[8]},
      {stage2_5[5]}
   );
   gpc1_1 gpc123 (
      {stage1_9[6]},
      {stage2_9[3]}
   );
   gpc1_1 gpc124 (
      {stage1_9[7]},
      {stage2_9[4]}
   );
   gpc1_1 gpc125 (
      {stage1_9[8]},
      {stage2_9[5]}
   );
   gpc1_1 gpc126 (
      {stage1_12[6]},
      {stage2_12[2]}
   );
   gpc1_1 gpc127 (
      {stage1_12[7]},
      {stage2_12[3]}
   );
   gpc1_1 gpc128 (
      {stage1_12[8]},
      {stage2_12[4]}
   );
   gpc1_1 gpc129 (
      {stage1_12[9]},
      {stage2_12[5]}
   );
   gpc1_1 gpc130 (
      {stage1_12[10]},
      {stage2_12[6]}
   );
   gpc1_1 gpc131 (
      {stage1_13[6]},
      {stage2_13[3]}
   );
   gpc1_1 gpc132 (
      {stage1_16[7]},
      {stage2_16[4]}
   );
   gpc1_1 gpc133 (
      {stage1_16[8]},
      {stage2_16[5]}
   );
   gpc1_1 gpc134 (
      {stage1_16[9]},
      {stage2_16[6]}
   );
   gpc1_1 gpc135 (
      {stage1_17[12]},
      {stage2_17[4]}
   );
   gpc1_1 gpc136 (
      {stage1_19[3]},
      {stage2_19[3]}
   );
   gpc1_1 gpc137 (
      {stage1_19[4]},
      {stage2_19[4]}
   );
   gpc1_1 gpc138 (
      {stage1_19[5]},
      {stage2_19[5]}
   );
   gpc1_1 gpc139 (
      {stage1_22[8]},
      {stage2_22[3]}
   );
   gpc1_1 gpc140 (
      {stage1_25[5]},
      {stage2_25[4]}
   );
   gpc1_1 gpc141 (
      {stage1_25[6]},
      {stage2_25[5]}
   );
   gpc1_1 gpc142 (
      {stage1_25[7]},
      {stage2_25[6]}
   );
   gpc1_1 gpc143 (
      {stage1_26[7]},
      {stage2_26[2]}
   );
   gpc1_1 gpc144 (
      {stage1_26[8]},
      {stage2_26[3]}
   );
   gpc1_1 gpc145 (
      {stage1_26[9]},
      {stage2_26[4]}
   );
   gpc1_1 gpc146 (
      {stage1_26[10]},
      {stage2_26[5]}
   );
   gpc1_1 gpc147 (
      {stage1_28[5]},
      {stage2_28[3]}
   );
   gpc1_1 gpc148 (
      {stage1_28[6]},
      {stage2_28[4]}
   );
   gpc1_1 gpc149 (
      {stage1_28[7]},
      {stage2_28[5]}
   );
   gpc1_1 gpc150 (
      {stage1_29[4]},
      {stage2_29[3]}
   );
   gpc1_1 gpc151 (
      {stage1_29[5]},
      {stage2_29[4]}
   );
   gpc1_1 gpc152 (
      {stage1_31[6]},
      {stage2_31[3]}
   );
   gpc1_1 gpc153 (
      {stage1_31[7]},
      {stage2_31[4]}
   );
   gpc1_1 gpc154 (
      {stage1_31[8]},
      {stage2_31[5]}
   );
   gpc1325_5 gpc155 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4]},
      {stage2_3[0], stage2_3[1]},
      {stage2_4[0], stage2_4[1], stage2_4[2]},
      {stage2_5[0]},
      {stage3_6[0],stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0]}
   );
   gpc2135_5 gpc156 (
      {stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage2_6[0], stage2_6[1], stage2_6[2]},
      {stage2_7[0]},
      {stage2_8[0], stage2_8[1]},
      {stage3_9[0],stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[1]}
   );
   gpc615_5 gpc157 (
      {stage2_7[1], stage2_7[2], 1'b0, 1'b0, 1'b0},
      {stage2_8[2]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[1],stage3_8[1],stage3_7[1]}
   );
   gpc623_5 gpc158 (
      {stage2_10[0], stage2_10[1], stage2_10[2]},
      {stage2_11[0], stage2_11[1]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[0],stage3_11[1],stage3_10[1]}
   );
   gpc135_4 gpc159 (
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], 1'b0},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[0],stage3_14[1],stage3_13[1]}
   );
   gpc207_4 gpc160 (
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6]},
      {stage2_18[0], stage2_18[1]},
      {stage3_19[0],stage3_18[0],stage3_17[0],stage3_16[1]}
   );
   gpc615_5 gpc161 (
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4]},
      {stage2_18[2]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[1],stage3_18[1],stage3_17[1]}
   );
   gpc1343_5 gpc162 (
      {stage2_20[0], stage2_20[1], stage2_20[2]},
      {stage2_21[0], stage2_21[1], stage2_21[2], 1'b0},
      {stage2_22[0], stage2_22[1], stage2_22[2]},
      {stage2_23[0]},
      {stage3_24[0],stage3_23[0],stage3_22[0],stage3_21[1],stage3_20[1]}
   );
   gpc1163_5 gpc163 (
      {stage2_24[0], stage2_24[1], stage2_24[2]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage2_26[0]},
      {stage2_27[0]},
      {stage3_28[0],stage3_27[0],stage3_26[0],stage3_25[0],stage3_24[1]}
   );
   gpc615_5 gpc164 (
      {stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage2_27[1]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[1]}
   );
   gpc2135_5 gpc165 (
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4]},
      {stage2_30[0], stage2_30[1], 1'b0},
      {stage2_31[0]},
      {stage2_32[0], stage2_32[1]},
      {stage3_33[0],stage3_32[0],stage3_31[0],stage3_30[1],stage3_29[1]}
   );
   gpc1325_5 gpc166 (
      {stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage2_32[2], 1'b0},
      {stage2_33[0], stage2_33[1], 1'b0},
      {stage2_34[0]},
      {stage3_35[0],stage3_34[0],stage3_33[1],stage3_32[1],stage3_31[1]}
   );
   gpc1_1 gpc167 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc168 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc169 (
      {stage2_1[0]},
      {stage3_1[0]}
   );
   gpc1_1 gpc170 (
      {stage2_1[1]},
      {stage3_1[1]}
   );
   gpc1_1 gpc171 (
      {stage2_12[6]},
      {stage3_12[1]}
   );
   gpc1_1 gpc172 (
      {stage2_15[1]},
      {stage3_15[1]}
   );
   gpc1_1 gpc173 (
      {stage2_22[3]},
      {stage3_22[1]}
   );
   gpc1_1 gpc174 (
      {stage2_23[1]},
      {stage3_23[1]}
   );
   gpc1_1 gpc175 (
      {stage2_25[6]},
      {stage3_25[1]}
   );
   gpc1_1 gpc176 (
      {stage2_35[0]},
      {stage3_35[1]}
   );
endmodule

module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [35:0] srcsum;
    wire [35:0] dstsum;
    wire test;
    compressor_CLA16_32 compressor_CLA16_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5de4d9850e2756c85d03fc681343d2214ffbbfd44162f7470add1e5b5cda0face5eb580f279d235363b8806529279102d3e230425dc24a26b61914ea301e984b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h4888ecc94d93d2b3848693a1dbcd24ca02123e444ce43230cf9752bb2e34f093e3a1a4a5ed483f138bea1659ff70ba3a2be72be77839896a1b807aa81ab4c4bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h72a9fbf2da01718fc322780291fe8f1486d533a6496762da99b82f04513dee70c7a83f46dc0d1d7635d222893f0151836fdad34301e5118d218889dc958a9808;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf9f86fd5e1b442863fd417b7da572586782857a8d56d030cd97380aef0fa2a3c4d03481a23a9d3ffda009c43a511889d6befc7b979216c862468ca6b4c47c81b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb51fc5917e7429108701e56020fc01ff6a3554e1563a5e84c71a4fc15b2c943a8ea9629921fb22f606c5e8c31c95387635eb962230e2a1b0cdc498fb56aa539a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc714c2a2ae78489c65f162fd994554bb2e4c1d928aba21d3c70fd8ba82a21eb81a5d7fca7c62f976ad58609a04558f3fe14f9724fcb46492641e7d909593937d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2469529477feca59f26084a7936890a075dc0265479b197c832395a360fbcb49fc11d998c675522586d50d9502128c38fdc753a05f2fba508127e049567d62c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd4059b3a69ac05c697fac4ffd326cd155e9f0a74c5b08c1b6f66cffb811d55cc566fc1df5368edbf5da67195d7a1862a4d112801ed6d60796ac08a9e8b91c6cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h53de82ccfc1dd00c4189009b07422d8d00220e73e485649fa69ccd63ba16061cb514c6361d7d04feafc258a470c738f7c90cc10a74a2fe662657b1a9a3735299;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h246d52d260d2560cdfabfbc576a390aebab1f2d29a4bfc9eb632c3ae9766628f8f37066b34f3cf6922478a9139c89416634be17140240f5fecbda167f66ccfb6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h40a8f70699e80276c19053a383351cab00212588f2a9cc398c23f9cd7487b67398fbde54d80cff01adf4bab373cb725daeced68cda690fd8fb2b4868514e4474;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hcb2b9f0478dfecea8a273871fd46fc3bfdb0989a623938faf96880c4c479fc6bf19e673de35d8b92a8925d6b90119549c1dc93ddcadd8fae549e7af65e33a194;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1580a35ded437b652c175dae2c96b596a1d1449864222494d4e7a33f10ba21d72f8f7e958ca8ec152296dd4381aa5f987e69e2124c86d7facaf60da2b602e85d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h96df8e146e5d10420b792063dd141d3373449cca020d91cba9846b7311b49dfb3d27bf5531bc0e939ee29d4e8e92191d6ccb0a23d51459b1b58efdac4096f12;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7eb2ac4fe569e696884ce9f18553aeb149d6e9d0aa5fe693d0b2e4f2f677f6b9fe55e994bf50fda3d824ea527e0f348eb1cc87640f5922bf8d405130520dfa9d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb7c50f734ac01c26ef72e11577dfdfeb58cac4a4a5fe6bea0ede5a19cf7f8f53976e3d68dcbe07c4695cfdcb0f0ac51fcbd7af32d2f5e854d317cafc7fa1520f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5f65e3bfb95509f3afd5a5901115928e9cb2705d4c01a779932edb44582b19cda4dc7260e2fff9b4334775473e05ae734a0ad28d3ba4bd3e66a92afee905c210;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc970a6e50002d224840ac03e5534a37ce3a040a6c923e4d8f4f3548c580a7cf178d6531771c69cdff76d2c79f309785ddd02e951ad4bf7a842e2779f6861ec1d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h88b01b8f64f8b89a4a48c572b11aa0506750fb6ea4dc76012d9824a1d8968fddc973f97b7502693fa733162897de16deccd607c6d783b321a440a0e2bfa4764e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf76232facfa8f5de9b791c8dc16fa2b71060414733dc5572883285d78c0d94d4615328762120a19a470125a582616b6abd3e16c0d22c456ed36f89da31a3f40f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1da2c4990916af1fd39b56eeabae28d5fc1c09f1eec28b5d06130c80e121b1d9329b7e7b9b1bf65ce58f2f3699891daff7c93d925db4e655fb88a9cbd720b2c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hfb4161437ac62a58bc4419fcd69986d460ff6875394f71630cf8d41aa9b06c328430c6807dab56be19dd13efdfb27b8ce4bd2d118e3336638bfb37776407e56e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hcc6676e45267b366bc79df5911ce5e382830b6031adb1596279f0e88c570bbf4852eb883bcfdb58957baa43f483328af2a06a660a3be080f78ebc7c73d39e56a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd55d1afa12c40af7ee3640218b25e3566307aab823590330d63af1a5a2db724fe85948c0d5869f4ca4c7da69d9c5b676b2861173634535fa91fd73189fa7ea34;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h862e6a857dbcfb87f41236d71f00040e1bd26bf1af142746bc75f4f1010a57ef381fc818d286fb75b84dc8d43e3c470e6f6c9b0dbb96df2e7b2aab0e3edd9357;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd0a4e3486a82f33482fe72c4d91f16356f6c0ae704ac223f84be53a8ade59b613d675b54c6f26aec17f72d8ac6c9f91d8dcfa59373becbd1f327361636c2eb32;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9cbafc23af057199b4c08233173dcc26da1643f149f50c1a26f5b3574b7800db2e8d8fe056f38f889aaba2f980c9d6d3c80df822eb35323d60916d2b274a4dc2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h19b677fdb9abbc3d9fc675fd75f172c21a9a2928896bb9e25a14b3502d2cba555273dbc4b904b603b90066d5d6b456feb3acee4cd4eedcbec9d019cb96b002e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hde32f4ba436e0830fb72df30cbd130532d4b4b72b1a624eb4c3ff4d93759737b8753483d31d937a464808df7b2754cc7c0bf0461029f3a22e2c5ef421a2f2d11;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h1498a334331e302c2a2521601ad2346be47fb5294a1f675913e3102b02f7210865dce88b0b45c4efc19111075f9377b1ab76f96a34b79fa8e2dfb35348247282;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf30ce659eaf5b8d9da4924d0a6a0671b9c29856b237b43cd7aee0d1da6a783ff0a2b29c1226c90cbe1fac7bbf5f8e8dcf757d5f4df2f6d868d7cefbe56fec7bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h3d8e786d1bdce61b15786135d97bfefc0f10e4396c919c4b1550829f8d95388972a11a432f509b558162fd28178d6b52f3c03f7e871a41382b76f12796691a05;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h72190e5c8796115682cc6df1aad8cf8e96d9dbedb69408bdba41c6465031ad268de7b8e1ced6bb02da3fa053cfad421dc425e2cf09a5e9dccd4f8d57ba43e965;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h42e31c17454ae860fdab85b46f1b3fd9876072f8364e41928dd1756638ae6007ea87762e456b255007a0def0228095b9ecadaec07bc20233a4c76f5db6cf0d8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb78c3a09907192fd157f3a4a8e514bf9d8dc5e81f30185cc8d42ff22d5daa084fe2db35562e195b7dd700875bec119b6d34a55d34786a0a287bc9947ada6d6ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h46315df19591a7c38818003e7a71b8fdd004e0dafc9bd1cc284c10d63bdee7666426874a039370351d53c19b475e9ca6457f6337ce8d28a942ea152a3d4ed52c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h25d8a9c4a8b6f125b3b80914488e83fc72a3dac30e06bca178387a231ffcd997fa651207d7bee6f10c618f38790e5909f60107f1ae2b132bc7154928cec73349;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd9fa2fe12adac677f2f48f007d4d694f35d4b890d124df7728ba256cd04fb3930d864bd1d326d39333c15dd4665ce7a82b96815ce7b369df0c00ac8e6e94b86b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb4a9958c00752b18a819217b46160206f4695d29effbe41fea78868505f9cdb9e3410f66ca8d9c3e1261fa279a1075ae9fb21cca1f123cffd1baad83b025a5b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'ha24c2bd721f2604a30f3f9963b5192f96ab6a575da2a19aefc3bd40994aefc9e6621ae2b4fc69c6c7066f2babfba86dc211691ffd26a086880bd63eb3f9fbce8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h8a88eb1052bdeac5781fde9a0bdc0bad9d7a44a114d0b0aa96fc1f4c200593aae8f5906ebb229951bd63d495606658384c81b9fd1dea5824c716b3ddb77219ac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5dc902bbff6a6a15991e4392271fb8a97c80624dc4a69adf810285026caf058a3ed1fc65b55e4670b94a9d697720c67e0cfd8e94e8b30dc7dc8a03661b04dd96;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'haaf6d43bf62794b4a96c036ece11673920c5047b90451777b07a8bbcc9e676ffc23896f6b38ad2f65478ba99a9f1ae0f91f3ac56762f8e677995630eb7a6d7a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h48009727f4f5a4ad47429dea13627b0ce485d83447674b6a325a7130e8d3351a641832476665b8fa7361fe64f00bcdcee63f66cc151e183b706b338a64d38d00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hada3c7505d082ad7ee93c410edeefc5d7a03d0bacc3ffd34512867608db14c15bd7f02504088e3cf1e0375b85d17753c98a7dc888d2cc4ab061582742811dd2a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2252353bd0ea9893e1f5e1880f2ec6535d02f1be9a41c49a982c84c266ae3f85f784f50c207b1feafbf3e5c076f61c00d270981a27f648cfc5f80ca70447b33b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2e1cb6b46c5a91702d916ca181e316f85bfbaa132494e0da0ce4c1c8c0747132251b408c7202355790e2672d3eb505687aca821323aa5ddb716643baedd57591;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9da383bb6bd246279d9a45c6c1843a0862a3ca9a639b96006c2bcb4445814e5ad0a3bd107dfb53a9169fbf9e106fc9523071ac8a6a448e3b8945f3eebb66ba30;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb074a393a4b9a5baccdade46933320947cb011497e17f450be0e276336cddb1882bf2944357dc32444aacdf00dbe250d86f3249b03ac7c41352454742d7c9239;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd73e875cdefeea8c137b6817a7d319638ef75143f446a9ca00a91aeb7af03d2fe931b529fa2b87acf34714cef21594bac5157648e20d66cd079225888bfe884e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h791c3098449ac933ae8222739232c49a756633a24c9e1d2d7d1ee63867b912eb3edc0fa4df6ffbd0c425665d4e723eba62280f90238affbaf389443dbaf3342c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf944d2ffdbf924bc979b3a0d0a8240775a439307433caf3f2ebed1f270c5f095283cf58711eb1092e7132b5558c70c10f13c3ef60bb775a8222159c34be8233c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2d6be60e2526261d1050a27c09951d1180f4a0dbf7cec2bc308f10981f928551346fece6c8f5cc58a0fd56b858d5e46f4cefa3b0c484d85c73c7a6885c775dcb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h7b15f81437b19831649ab690a9ba6cfcf9ada6c1d741ba0d5141bf0bd01a3d03d5efaffed169ad4bbc5d639a706df948e388eb5e23611e898c60ef83ed56459f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc8be011631c03e31657e5ac5cb35eefe7db87be9e289d4c7f4b12985ca634d11afe95539fce0cf053134c76f45217d9907d7c6cf0da1a75f9fb4d42d89754c41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he396526e5f11bd330c0e8e9dfa86fd89479d8139f0d076886ac0bcfe2ff13cbbdc996c15ec981616a57fb8308d75c4ca62f5007f2ba4f0194a1fd69f8726b2d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5fa5263614cfafa83d7b0f6257a3ed48171eb6a903d51f87f698af573aa4c06ad230de0689f70af2d7ab34f16d3f2207db087fb2c724a9d3e88b99a48a9352d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd330815a84ca1d0a0bf16de5414e76a66d73997f80f8f5d28e7ff4e6dbf63538256dd39eecbdd74c50f1052212ca691b43a9d2314596afc7e86793ae2babdb47;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h732d56e419f4bfab007f39ca80c035d70970639e5748835d890bbf63218db399246c025e0ae77db3fcca383278f8952e99f6da1ef8e9a402f43e7946f1b3b333;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6afd4935335bbd548a4a292de234d0609956ca9850c9d80371da644e74a5efb538cf6b4ac0e00c33f4002d6bcbf5dd7193a21c452655d036aac1b37ae9c3ec56;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hfe4279ae573176c565b7687cbc48b9ce127412cfc55e2321a02ec46843c41af421b9204926270e1905d7e0787a269741cdc4f20aecdb0283748f0832381b58c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h912ede1b0a4bdbb0c89e81704a96c5e5598396f1d63677694557d56bf93aaae23d904cfbac94dd1c58f693369e136f8d666649ab2decbe0fceb1a4ff7eecd099;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc195f84c4d2b59de0e292574cbd377f56c3520af099e04516e2ce9e8b5ce5254437cd0f2f1945fa3b92affde8bbbe4ebd57a961dfe05e6fa34151e129b062038;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc28585ce371107a2d94002ed2900c8743fa4ed1aae143bd01ac8f916adfa32138ca5e0cfbe4db60939eeff59065297353972ac5d675ff9f1c1015b2c38c7b2d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2d202c6326f5b42c9ebe6d7a45cc519e565879fc64adfe1ca3f14dd817530b6731c6339f8c50bdf030d99d366bdb38394b574d315db28f6e457bda6ddbdcf3a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h91131547102233c9c0efaa238520179fe899e25b725f3f765df05f3feac37a2ecb93e1112356f34754202ffdf5efbc3d3c33bff1da85d9dc6c0ed7278b94dda4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h886ce1ee199295524eafd0793f2d7feb9622d5eb955bbdffe91534a249932756df13ede5424d066dad7b8597e09e910487bca2258cf8259d5d6024cffd573160;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hc79bc6921bb869cdeaf00482432bef817a67950a9af6598b767d861cc535f3d1a77b6c90380899af5e6da258695c05aba169332049b8030ed58bbeec3ffec495;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h614d44ff3160be7143744712275eef50689f6b16ecfc554d677003af7f0f0bf094b0da58668f3163a44fcfe8dd4f02d4cf0fcf63584da1f05096bd951f6f7192;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'haf7a62864516b5f16349063462dcdda4ab822ab1985fc59dea3dd38730608e039186a8192c950f6e9121599a052e0bf8e23a431961f9c7e2706364748ba1b998;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hdf12f843b69fdf429321e210e75d3d87771c715afca46a1fde174363f391d2572b50d7f1ee28c13f5d19886e81341a4cf7f61d4451a5e8a81e8326ebe3b154c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hb67060c9d08674694aaf260751f37f7245420a92143e2145e9c1edd78fb556b786d513435038356f509c5ccce2a5868554dcdbc6288f1dbea158e2f057b3daeb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h887cb1d9140ca7923f6da1591b46d6f8b6e895b0116c70891ea8a3c82c715e0b397218e593f442515e6479dcdcd89288a5c19fe700f2e95640e19db7fe64ae40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h27bf44cb08a197cf6ff8608e316c6dbbf8f5ae56662da8a95f9cb17f7121cbde5b28fd45838c80feaf23b4fda2abceeb5247110534544b4bb535f5dfaf67878f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hf9992cc947b4ac01df769106166cfcb1fc552ae8089dd3e8b1aab5c487383c6bf2e9a97c5ed9f633b3129546eed4108dc82330f79a22b6f9bfb296917baa0a3b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hdc6e17b716626aa94ad7fce0b7109f47578e520e706158d4abc1c49a27cde22e78cdf50564c818500a44161e46e54e790d2b67a13fab4c95dae408588464456b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he2bf43c6fa092dd132bc11a5324955e6fa65101169c5e339223997cd231568f13be69eb6d8c14183973c4d9e64d2337f7b746940ffb73d5cd6f91f862a89ee1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h743b98d5c39f6120c8a9d78b5d13b4fbd1b67607106baa3696126f96d6293ec121d770ef41e3e0e5c6dffa477eeee38b5692a98c764e849da5fef74880437a36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h17df400543cdf723b133188ec524fed0b6186d60e6fa4b76be483a7bd7d2c9ea6d557db090d60dce6074d7bc1fd5982097cf888340facd8928264b302f6e191a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h5a95e45f97a649bc0fb0e777ced21669436adb691d9eb199e0d3c85251f148f404f6faadffc0ed5095284aa93ffd1deac48cceef3b42b2cf1b40d82c498768f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9cadd1935918b4a50bccb87e5b1c8f9314515d50aa15e7da9f5de315bc9d35501c25529f883f6fc7a77e4b6ebbcbc7e4cb3be1a3ac001ecdfd77cbb11412e167;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6917bfbac429c883ca6a7984229b6061e3b1fe7d64677984d4e51acea09bf3f74c6363692d5f112d204f2093296f9e202016986d67a9e1b70fa11d137c3ccd91;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h469d5722f7455d13b6dcf691ec95f1e78c290b6915098c79b2595117c640e4cafe96e8a14117069728d9f071becad493cad2e4d573459e2c47376b5106b743;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h24da592abd02f2cae7a4d8451bf981f13e2bc8ca46503e9054e1aa3684e815d7fd5b03ad9ee8dd14dd61a98a999adca646ac5e147be6b5fd1d56849a4cea4f4c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hba41d5ffae2d5a4df9ec63f506f7a83bbd896b659bd218c6cab54794ad1ca1d7808faad1d5e4836b5d016e8b2d8f8ecef0d438014d23c79fd1d7938c00ab4854;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he96b80116fca28d8fc92b3ecbcf420619cc560365da9ecec5cbc6a661ed4e610a1c10509e66b8cc704611eb37db0349b257467e72d0af7d416142e94207a4cc4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h79e46190310f39fa4d8db761c116aa8513ad9e4ab26e69d5b79d59f2f66eef4044c978069746b9c350783ded623773f36768ca191ba60065bfaf67234eedf7bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h2ce35c3e4adab9998a940425b0de6e0454b3055a17bc8ff2ea57a606e7147daa12be29b7f0d7040bf90b08e42f3db95bd1c9ceaa03381cd3e14375bf38575710;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h79cddc207c58cfbcb2f8bd7439f1405cbaec8dc6afb1f1c05c9c45b9e8acdb06aaa8937bf74655e88fd66b1909fe5e64aafa3dcaf7528abbd4811566a1176050;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h9e9c0d540c58d513218b5b39ef71846bbddbcb3d17fef8409004b58caaf2628d65df7b2026b68b82fe0d0f878e4b4a91e854cdbe09c55adbaf6974c6e444ef4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h87277c7b3cfae36587a393ca4d9d173c298c908c78dc77e3dc2f01c49c9e2e7bc1f2c20d01899b2357d32d27d850c2d83aec8bca60cd10bb2dadcd95e96e8d16;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hfb7c6cf52ef2552206ec51979e9e0adc47e8c4eec465abdc1946c045eba33595a439e0e56178c3d2b7724cfd668e67a4006a596c4d8ae700d06d8256cae7d030;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h6cec14c31ed18df958530f7feba4614dc87ce38cffa78ca1efbfba4099e3eb1817cae7523a9fd944117c87e615ea546e7b70f980e794215fd68dddb4315f5650;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd197401e13fdb5c98451b3388908815528d57f0f7cf27f09dcb8c02a5c46ecc3f6ce4579b89b990512d09a3f8a2c675b83055a3af9512dbc5bab27b71b6364ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hac8ec8b6cc079793cb89c0955d74bc1269a8cd3e9d5d675e9a65f7bad654bed81ef95dd536e13a8ae4b99b6c8df707fec0f5aa417da97c09357839f75976ff98;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hde5515b30b0092c9b0b92d23624688967a6a1c920c78a369942eb7a9d6080b20a9636037023b862280dd3b0dd7a064d42cbe096460e13909ec196f24d15941cf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'h750b33c73328b38b2e0c4147078eeb7caa83e0a14955ab70dec3f3f5540511467b1cc739466d3414d88cc16d3b2d748f4034c1e1f05d0d2fe08ee74611ddee00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hd6dca67c594d08c4079e0efe97401adcbd27326b3a33597e2bc46eb4d6b4970b8e91f0ffcd800ce1542bc50c434b0bd973061a365a7ee860ea75628dde3a6fe1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'hec76f9732cc9c1c0be65051c9c23190f50f37e1ec39ee928f938ea01a8253eab9eaf7b5bf851e9535985bca4e18c2940cbc3d04fb247795f5ebc1fd8cb87d21f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 512'he1d9f1b6e3d6ff13425211d9cbe5d3763d1933e260b255ecce82ca047a8f5f13fe2f3e081178898de0a5676f4f43f4f59fe9b7faf8e107d9a8e5c6ec501c32d1;
        #1
        $finish();
    end
endmodule
