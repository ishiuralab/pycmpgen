module testbench();
    reg [10:0] src0;
    reg [10:0] src1;
    reg [10:0] src2;
    reg [10:0] src3;
    reg [10:0] src4;
    reg [10:0] src5;
    reg [10:0] src6;
    reg [10:0] src7;
    reg [10:0] src8;
    reg [10:0] src9;
    reg [10:0] src10;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [14:0] srcsum;
    wire [14:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ffffffffffffffffffffffffffffff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd0706acf0a12b8f4958995bcab1233;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18d12ae57aaed73e6f7072b553285bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h367811b3d412ae1009b2d6ce1b668c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hef46473d7c57f2631bf4207e69b1e4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c4abbef4432263e34f3ad2f79f07;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a990be570e25690820a72472b7d50;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1255afdb6661760f054c50703aa1a0f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2a4135256cbf32140b2bff3287931;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf5854ebb358d954601df02ce12c662;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h69e2750e608f3c173bf8e4ae2cd4dd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e7fa36034aeea67c079ba72c156376;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h156ecc9dbd57d0942d9938257f39905;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h162c95d5d8cb3fa548a869cd2eaa960;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b804cd6c9293df0f759f27f22e5f93;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h671ff5a013b4b559bc3383c7974b8d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h668f06e178ed257b511a5c0a68f42;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb43688f57ad7cd58aa34334fb1302;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10fe8af17cfcb2b2959194d1431c933;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h505657c6534defbc180305807c9086;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb6836c64f56f28cf06b5c68e626e60;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e0cf1f1f16d15c34201108f12cbb93;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b164ae374d7e9efce62c6b95ec1b16;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10f4074b03b3a78d527dba0d20dde83;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5f3a8ca871993d2a008e810a43a648;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce5f2ced9517364207f9d26c34aadc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4656f55c1fd7702893442e77bfe2a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb05555ef3dc465ff0ab6b9408865a3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h170921e1c7b121b0382224e900c02fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b9fe23f810c486ac5a5fbfc6eaa76c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1192c2cd409a9f03605573f1f02d1ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h164dd41beb51e347c60c8926ad78a20;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1893680a09b337127f6b4d95fb4f34;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha0d6b59527ff939055f4835e644ef1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d20a92d131b8df90364ca22ef5c930;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h85a0bd75154a8b91e02c3dbed68f65;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h140a251c0749387719598d6690210f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcd444b3cfa3d7f6914ad94ea9ac52d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha992b27aaaf369b53da27685fb239e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7799703d441bedff29eda3f6f17546;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heef621d1ab9c6f48585bc96ae75af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ea6c1bc31f4d37185e683d1485afe5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12cd113cdf7b1ec3424aaf9e39a1de7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc1e3c231f0b25fd46f14db9a13d85d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e97054f6d052d6ff6919f6b32cf2a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1927d6a7cce4d4fb9cd46612643ba03;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a1dcce6686fc9ac6e922c6c44f59be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h181ed4d89910dea904417a581dab34d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10906ce953e1e45930a167a0a64d91d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h131495074336a54cfc39f47026f776b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h42a83c17fdc10f634e5bc770c7072e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1902701d164badeb078b249911aedbe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h128f82a75fd46491af2a5db536e8790;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h280332bb6d9a4c39535d2a2d7e1d67;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h108e063abbb5202e2eac6ff908e8662;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19c51b851fad927a6f4c3041fb7c29f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d5e66521a8e89d2c3923dd31edd04d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h853995b2b174391f1f1f1908ee311a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6c58bb53ff054d5542f6ab0eb048cb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h166f81fb2400a87820e518e96a2ba13;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cb9890bd4836d8ab2581737118cd93;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3391285a75b861c17cd4ae2a90ab20;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hab5ee67342512a687c22b42eeba638;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc87012c07ec8f9871780bb1e2d60d8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2e089274db6950da829aa3ad58c559;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15c38bc88e6abafe76a11ab54ff397b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10b1b408f709daaf49612b026fbcb6f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec4a55b1fe07370c90845cc5d117b9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha6fc7df9a83f02427feb3574d0dff6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h117d64762b16eed0fb5097b1e6a73ef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90bd9e23c8972ef8e9e692dc8a8a80;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8cf5c74647c2bcfc652f4c94c17880;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d5c82b075fd6ad001265b50126053;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h921543130a5c9812162d10d2a28b71;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a985a8666d81d416dcfd5493fc7b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17a7e4fd735b612bd4dc8915b24291c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43fccf8797f7b0f927baab27f349ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1efe2cf1f43df121ab53aeafe812b8b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14c935337ddf74cadd8cc2b3893ce4c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d851439b271faafdca8eee929505cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16dc08278f03790e0d131e118843dda;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf0a6528885ff153a7832b8a8b04bf2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb884f7bd3d97dd78db8d71ae3343bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8961b9bde9f7317162d1aa9921d87b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a3a3f14455d9d7bfbd5db24ac04bd2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf5098f1d11dc8a1c447e8feee182d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbf538131e25f177d5c6e01521d38c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16a504ebe7defe5bd3548ce3c723f25;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7eaf9db99b728be15d682e33f3d49c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfd11964505981c4c338498655f9e6c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd4557e09d6630189526ca2acf2673a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a7d97b0637a954df6e49c238c5314;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a6a7b43545d2e72e24fed86ec9e31f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc6bc2ff075183af2a45fc1a7a3a881;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145f13612510590faf8ae3cc2ec27f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h42328b03c34917159f440d2b421f8c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d79405647dd013291ee84c3bf18a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a0bcbbd1a456359728b4c5dd152618;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18260796ad917bf7d30522b2088affd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h156642fc4221a903bfb2f5daa1d10f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h153dafb45c3ee8c639457709ace4916;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heb99f856bd818fdba04a5ce71ec76c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6e574c15514b2a4ba504fa772ee8fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2213017bc40a885c05e3e50f893aee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd80b33dac466a2eb9f5d621280374b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc2f5750984429aee4e349d3a60bf03;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h64c029db8f7c1cd66816deb8c1e2d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h41da981135a8ce642ca7f2f5aa0cc2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha4143497947c0f94005d90b72babe5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17d663f66816f6af68090f466379ff9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e89d6ce78833012edc51453111b30d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b420d095bc225cfdb533a967374de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18d80fd355a1b5f3cb63f9034862754;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c2631b5ce5b0ab731789c648bf872f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc80c935bfe8ae487b5718cf471331d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fe404f56168b913ace8bb33c3a92bc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1407ed1cfc5fa3a81badb9a3a79e7a0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ebbd170e5b593b23f5e94892866565;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8afff79f93a94fbec7aeb77688efc9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he814630291d50b6dc6896d30f2e916;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12e93aa2dff1999a8f45bee53d5e729;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15334710e5cd0b56252b86273fee5e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111c682ffbc889f6231585d422481b7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h72f7d0e9ab31b8d6a200631e4536c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d34ed523a3e550d770f620bf0580d6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ef9cfab8c0a7cad4f7d5a4baeca14d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5573c1ac5d8f9b0fb8bd4f9d6fe8d0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h147d8338ad1ae4bf0e2e720f9e61d80;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13058c6308c0de550210e4f3f88d84b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ee8acf23ebe86df62283f981441e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h193902e2b8c5ab2b7e836eaec8d399;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a963cdb6fb883281ab29f8ca554fa6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8bf7fc2c5d659c86f2d1dba23f103a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h139ca64d7ab862ad2c570b29754a8a0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4156759292e08d7849b47b38af7d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18395eaa8832d0827f31787ee283c18;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfc15cd98ddbb66f7034124908ab172;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d89a2ecf701cddb6856a46320060be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h449763269d88a12a37140cf511096f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h148a6648a66a5f1c233d72792e95656;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19220c3790897f520b884416ad6fefd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h52829a234af66d9538cbb6a4c2beaa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e82eb54a82249ca4fe48c5ea5d6b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h161b78a8edb95daee4f073fc40b54cc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cef6430a1081e8e8b0bd1e87440903;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1efa1122e6ac993089173fb0b058803;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h707bb36faa9fce44c36b1c1f0287ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b9822f07cb52bce6733c5de4b70ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1973313a7d56113b024c4ae00f337fd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a6cde403425c1ac84a068a04ee7a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6b15300fe24bc210b98cd01eac460;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1614802b890a97e54e78047c9f1d386;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h115b603e292e7f49100109fbf62fa74;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha83e4e8ac194c182e08feef0c10b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16fb6240b52479e4acc6c5b67dadb0e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hadcd9a5f1083c4c4c8e7022fa1a8c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h803fd2873505bfe767b08877c6bb1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h855131839776003bfa86c5af151888;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe8436744a5320eb795c8a35214ff1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd72798db4395cb4052e5f012674551;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b62afa993e2f00805447327d122013;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h108d2786b98b570e0e2d8fba226064f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h411835317a342c8bd3d225128f992e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd89f8b6a22bf9de4958c87f3f921a2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heaf1e8562077e590a10274ce6eca31;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e9714438c5ca5a8fc81cf6cec0491e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ca60b64ff2f51034dfce1a5539a96;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c560bec7fcec444148f6f3c8005be4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f9d5a49a0e712a8c10e28c93e96a2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e606e5e5f1ee950e097db64f1b2c1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df9d11439887d3d5c5983e65904476;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc8108ba990824c7af31e85aab0551;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1323fc423b26aa534fc32aee4f1bb1c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h162d347004d93d6c312444096a751f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h280bf37a8f7d0e92c0236db536b00b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha0900e61a6c83c1d9708f742be462;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b5978c47f0d0cf247f3ae7b601c511;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he2f4b75e67ae31b705d829cf4944a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1600cc9ab58a8704e035efef57f07a3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16bfb49ad343c47e310ac81980a7d52;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd766b64575d316565d20277bbcf8ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h129c9cb4269c69210be8fbc4e99745a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h799f3b24ae0083e41226de1cca4fc0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11eb163e889141df57979f8f7d8836c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h805c787d8a0ad0d63973fdbc7593;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15dc00be033304964ad9df9a41cdcda;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb3e300f330bb4c2a3a14dfa7828bad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he3c0c04b45ae4dfa4fbcd82217f44d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13746ddf07803253b5aa2f4091922a3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h612984c108dcc4c7679fa569a54b88;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1200073e11b2a4f50ae51a2775880ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h183739a52d2c9cce4e52c1bfedab14b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5410d4b4c9346a73b2cb075f165de3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107b5a8664d3e99dae5ce2c66493afd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6713de489f6c4fb47958e63c7cc20d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e309144d8bdb048e00dc1f404a62fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h351974719b133e83fb4a77c41d42c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fe3151356c3a816ac424bd7c52c95e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33a24cb4b81c6f3e04cdd64ca9a21f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h83204081a3ee74a9421e8536337f05;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15434a76f8ca54c3f7201198c9e229c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cbdb8abda0f56a4cb577054ac6a39f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h171b7838a9edb068733817c2655cc42;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1319d5d4c42b4952468a9956088cd94;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75dcda95313c082b4c0d6e11974523;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ee2804421d40862b69a4d8e235b848;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f79da551a72653be81a0ae6646ff6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a871ad329412dd2791ebbb811329c2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6e44c30ff078ab95c37736dd96c57c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b62e5d9377112d329b8591c9be0e92;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha34df635278b858f7cd4aaf88d7a8b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h170f4272fdb71696b8e36ea31c87881;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ed4274dc3248a06eed360ec972e72e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e304e31e38f87da1cc5325644e230;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha54d070335e178746da9760e32b4b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa879e6c4eef0138139ad319ca968d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9c51d85855224be85414859dcc9f81;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f62c8585f27e42bf8221143f15fedc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hea23f284e4f6e77e665a068495a15f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f47621e938cca6289694e522b043d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ea579b00dc285ca3d214a255540811;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha7b941dba3851e4fda05a0cfa6d60a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75be682cdb974ec648116500c57c4b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h175c3388821773af3a05281511f5d03;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17542e39b305a3f9b20aab3562b18ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h214bcc14258a1c82df201d263bb4d8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h128ccecfd9addb65a0cf450a925ddd5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc7b8d66d9e941687e24839b26c84b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5dada654d89d7f748b26b81cd2f761;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f7e5dee5c2df00f16103d2fd3d1a81;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197190894f3f3b7511123f0fcb8e469;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a80a7e9b55e40a3269a4b1aeccfa1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h123f24d3eed067de11bfc24b271e17;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha7bd44a44d32e3e49efdaadd768b80;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6cd29c77e0014ad96ecc59d2fe469;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h324c326be395ebe89e1c014ab0602d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159bec8aea5c87ca2838851be879b91;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h190bae0afed6f266d5a1c7e08b127b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e79d350e12f6b674b9149d5343c5b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5492279473f66a0a8fe8d3a2e525c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b6e58277ae31164227e041e533dd00;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f17c8a4b16e2db3e7ac87cb5718df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7a52967f3163b52550fb630f51949f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc97f900532e9d6fd3340cec95f4a83;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h69b5397a0e2dd9c4a8d0f88105c3fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ff96f83d9b61bdc75ce3aa0fe891f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1142271b30f9cbbbe5df93b3b283c1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h171429a8bcb22a923f40cc696930f7a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f8cde14edc5d6ef1795e4d49c8f2fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb5073b8dfb220b2488ea7c44ec5a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e4ff7b8667250e147324d95a0942fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159fb567ed904867cd50f12d1dfc361;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he61884e24475cd6e3e2e45a80aa17b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1025cf74271d3e024460d882b88ba99;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb5fb525499472e834c4d8ec622329;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h86d43858c54fb94dda0ccbfcde5688;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hae8f44587eac8d88699176c5e5f96b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e40c78c63eebb36d4325864ad6c6b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heed188babdb5ad774d5f12e395535a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h314ef71cd40908f249fcf157050e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1744c02ea3c400775f3d6a60d85e488;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3c031dbbeb794069968304bacd4070;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b8d85ca16284b233aa95ac883d095c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a69b0e25fa6881c20628b11fba567;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15c0974c935e8067078b437206c1cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1beed8d62160172e8b95c26db8a3b7c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha37b66b67fe8e9352d8ee21970604a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f54d83dc140538be261e525410afee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb0c52d78ce00777c2772ceae2e432d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4b9eeafec4673b8e8bde96ba48804a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19db116641d2e84cfbbee262179eeab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a819d3f1439eefe136d01f1f3a9324;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19ecb4478ed995c6a38a527ea7e6d21;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe2e80a72afbbb773b542ba55093fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha3a4d5c76273cf839d12583cc803d7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17148d3f0253fd2d57d83efa058ef8e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fbfba10f33f944565a592f873d3ffb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ead0589ead71c884052569d747d40;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf7f0eef38b99b2619d422a3c6f7858;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1606a7b120e820675bcc2e858fa2bb9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb7016f727b8e2544d1e4b2a125918e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12189496d9c4583ccceba49705dcd1d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hecf4c680dfc7a3e3dbac0afb540737;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6bc94ec775db496e18556f1f029e3b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f38f6113e04839aea22ea1de7c22a0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b53b70578c61ad0ff373514992702;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15ecfd4720ef391ac1b03fe5527e188;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c26bc9cf0181acae209462080975db;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1309e60ecf7ce79eb6ea1de89dc1503;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9dfebef56cbfefa00c522c5604fb59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159a2767b9284b262e4ae3c41fd6983;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17fceda42878c12704802de2985a79a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he273c4380d32c37a1e8d758e8099af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e13ea6acaa647bd7959eb9a3853ab5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h196980a298088498ad0013134278bfc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17bb6230c79b665a46da68ee7f5ffd1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16132e3eaa03c65f4ca47195190ec93;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h186cbc1b520a193d46352e6431b69aa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4667b0209ba9eb736ccaaa140520d5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h29bc67fac81129fb828b64f8eb8c56;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8f38705c8d1e797c341d61ce0828b7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a2e0bc7110939d98d034e5510e475;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h36f807b1d6b4e608d89608e6996194;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b363284f3bd3aad85f3d7e6f6f3ddb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d147ba28efab4775d08e4fc9c08c23;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18db1f773d0e1b81eb3dd85105ce38d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haed8d050c5515fbaeeff5c4aab7ce8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c446cfa35f474b97f32ce7d885caf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124b6d3ba981ccf2f86fe856d77d1c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14c44422b2232e963c67b2bc4406a49;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15d76681194850219385d817a40ad1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h152455e4146e446bab10666688cc5a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15388eb500a5ec3f373a3eb50d8bf8b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h32c042399c4677742e186431d63e00;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd35fe6fed7da64c374374c15df515;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h95b88da41952b8c22505e43018835c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c5210937946d98b207915bf2ec72b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12577d7c18a0690d3675ca91a746092;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8ad01be18d5fe936c922b225f4680e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6cdfa3b8994779d467b65d16e0842e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf6314563bb09f37d35abceac316418;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he0c96dfcd9e925d075802d797d208a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11eee17845bdca053b654f4d7aad332;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd70e13c01b53ff9cbd18c6d009967;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc009daa7ab41cac9f7b0d0a34eaabb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2bda15e5c5cdf0be893461a271435e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11d2e837de9293b57cb77b2e8907869;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1503bfdb97cf66621c193fb25730c3e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha2066bfb886bab190e58f87a44f9be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a361779ebda1f80b4e6ae3ccfed953;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec395b620bba08f714234a36e3309a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f3b3d79c499f24980dc006e435470;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h143cad7e09c2bf9007c982429700226;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcd93b646f5bde25d652ecd34808129;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc0c80d153e52995061501dd419c6ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90903f99f8d518def939a4d84a9fd5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3000f06adfef8b1fc2bbd7e1a7ac67;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10258eaae8bf55519305edbf33341f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9d628f7798cc5b13a11661ad72d002;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1861dda5ba8153a7a6f9fec6acfd6db;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1361069d06995f1d3d94fef369719f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19290dec704dbcfef0e28ee6ec6f7e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f33874de78141fb26c5410e08d6aa0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9e5b7e33bf1f58d48adcff6c8c573;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1412ee3791a021468a3c57d114a3c39;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf99a628f470709518f7c5dbd3248a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he1288d64b84db164f1a5781b32a25;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he55a0fd40e9ae44910211558e1cde4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b36b7de572a2874ba8e68a0b4cf72a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e05665bb61f143e63f0fa3173a71d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h171f5145be5f637f5f3b04eed8ccec3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h151008ef9ce4c0c7f8dd40bdcd62075;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a56b59096aadc77b74dbb5af52f20f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a877f7bbc60ce03a6ea87e7f5e6b20;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f4ee3c3a841cec4b00bc484df9069;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1890a91b5d12a2fb0b28373ffb7dd6b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ece118b11b233c965d08db269ed704;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb7d3aee973e986288309ad8a8b4e16;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19fb849eb865069335217e2c55f63c9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8af6e4cb8b28495ab675f9e9dec6da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4d9ca4cde3ed6faeee2e7629e57154;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2dea58be31a1dd5b3e9bf111713646;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18128484b6df40ba29e3d815e4ab1f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10a5dac365a68e7a54d44c7532f71e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf11f8761ab64800c7e36153c889470;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13484dd7ebc61dcc1d6906966abb8b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1239b7399b0ddf9d11e81058e13af3b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hff195d3711ec0c30cc03df345f395b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5e11518ecc46892b75f2f5a13efbfe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1141c33d1c4f9ead9727883569c5545;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h158f887bb12011246ea6a9e92525a14;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hea696f61b580a337515cc566047341;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43c06cdd0b9535e88b9f5c651d2601;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6bcaf67d396833c341d294ab88dbad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8b2a6c9d8360926991b0e7bd030427;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h162a6255f5d23e87609bef6e84c41aa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19f4fd395edf50404574badb36ff20c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb6bc26307e3d4a8cb5f7a3a936bfb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1369f49a6dea460a749e762e9c25338;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a93990c0b99be55727dd99aa76a5e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13b60fbab63201bfd0cf1b477afc5a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hab195f5c92709d1bc88104d8d32881;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d558807091a8c7b1da6139d5a572bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb918af70283e77582abde68232e1f6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12794413896b7e63f301c51f13fb8f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haacf9dfae75c05d63ca7971c5a1c4a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118460b34b8e0fb18975eb5399805dc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33a1dc69f66109bb162f8d483abc8b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha9b3d5de1448ab4531ea7985a5289;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7cfc2d14e9559c41e6f1cecd394ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec6578c13f80f72488e5e7a2b81516;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c42963949c5f51de21ca0534528a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11879c04a2ed2004ec59d6f478df5e4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3cdb531c31f68385bae0c4852c0c6c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12e1a5a5f8d365645926b822818e88c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11dd0810fca601adcc456b5b77612b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae3b001f75913aca80435b6be17d9e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8b9d5975e8e8fafa859edf0d064291;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7dfef16ecca9c34be1335f0fd90dc8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h220712744b58dfdee16d26f0ed7e36;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18246f954a155da61b02c30d89f8034;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13288f0a6ca94a45abb834b5bc0b1ee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hba33caf9f3a0070aaa85c51146b410;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h131450fe80fa755c4068f45937a1f27;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d1c3590a20926b34bd2d23f304bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16559c2f19fbc90dfee2098c4bf96ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cbc2ea23115c464f8e86b5d986fc3d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10645236b2d30ac01a8465b061bee82;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9eda03fc78ebc4e6e308eacc64c0c0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha6f7574522b0d576495a5630681542;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7c8bd93ff81071ca72a4fc148f8467;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd9c1d477b6fd86b7531e739ee15e4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce30d30b65e02f0a3528ac27393f02;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfafbf5886a32536bf40b682e264bdc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h527dc05f6cb83ab01d2eeaf8f043f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h683b3171033846e1f9041bc11ed233;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d1d08c3c5ce706288c469a000a9012;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe3b5ec7e9a3781da207037ab12e2e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1403916496c6a4d0e23709da76195a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hceedec0d5caba313dae7017b938f18;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1170389da800927c65d3eb47a354781;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e20eeb40752af38bee02efb4b926b7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bf9e1f5411123bc6169d8d1132ff22;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5bbf1eb77cdcd8dbd8700a0ca9fe9b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7695eb36acc9a714109bb360eafa05;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f97cd255b12c853e3270ca6c67366a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haf65b54d2f8f23d5bf3b7e3f6c62e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e8a4ce4cab19b8e74aad9b60363b11;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c43bb20151964e84fe03900cb987ed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc91d30426dabfb49781a0aefa69ed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h28b2fbe7e8e50a79ce0701e24622d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18630c060422e75de303d15b8bb6b13;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159ad9142faeeb283da55ae2e6f4d14;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8c41d730c96fec9fb3182246888162;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d58c0d29b94562ffb1c2bbc78ff21a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h130ce5ca10e8a5ba6c7a0dad1d33d21;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h390548823618f4c3b9dc6cf618d001;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2bbd4a64c9d0cced74e9f952e2fadb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a4cf17e5637082520982ca5db84f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19ccea4357a04adb308fbbbdee34502;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bf8416657d91f8559c722acf7d17c9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e6ec71a104328f15ba17a41482069a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8c7c182e69e4f016e4538be937a8ef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h113245adbc02d7b0d9ea7d4d9313885;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h742681cc837ab8b0b2ad5ebbe34ffe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf05ad56feb40db8f45be459a32d904;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14ddc7cf75631752847d6bde6b79758;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h934302462153d44781562bb869b1c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ba2d2c0ef18bc90ba602c57afa46c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d34544f232840558fd1adf647c932b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1336314b8add76aec44f2e42806156c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h176e0646c9f088e3bb3e7d4ef57142a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14567982ba876117e3d63eed5a65d15;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1687d05adf5d50ee804bc1cc08e997;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heb857b9b5d97301273efb2d3784cd8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111cf532778b04e8d0a603e7ffd8c97;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haea281e7d75e071426e282de84de87;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fce8235e99217535a6f8ff8bff7198;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b9db21e4490a0045350c869e8c221;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfeb42d79faa837d45a6dd5b6b2918a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h78de0598fc997c30551092a32efa3f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eef2b63c2835141a17ce221cd54b1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdc64f741159e1e21680fce33b0249a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16062bf2831ae23c45729bccccd3bfd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h168abd1caf97d2f3588c044f13d76;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c0c6078d2aff46d3c4a28bbfd964bb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf04412b8e004c64688ad2ffe15b755;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1213c8861b68b131f1a119692fc343b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11a5bae4e58eba44747ddec6dd3fdca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcea0bad2f915a1d19881bd3a8379a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b7053085c6dc0da86dcdf2f784b3da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h226a19376aa2b8fa744768d9dbe889;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10653c460b48ab7c71dba3dbc9887cf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1091ea2e7df89e5f78852953132d0b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5b5766d34243d9e9770ec3bf6e29;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3809a7f43389f89a5f993c5bbe8d36;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he49310b1ed8434eb0514ebec08e89f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha9be931830f63586530cbaa93d7eed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf9988459cc23b13532f5693412e5f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a5d959e8dd92ca51dab2bfa066fec7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbef1b540d86a291d52b80e53f427d4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3cdcc7b5d23b9c8e642db7533cc393;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb264b8f038e6165e4fe7997e5ee74f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h195b502c076774c4f4222ffa3cd171a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h177a7703a6c3ca69ff8b4f4e0ce0866;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13a0f984a97ab54eb3dab796bebea34;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc936af965df56847e9f1e295d47f9e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fa9aa4fd5c8eb3ea71fb0bffe86ccf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc1f938e11b92ef6d32f842dbca5e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12cd33ce5de0bc4c7349df13d6c1dae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h152a81f048bc053d8dbb28af7f10312;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17e304009ba2e08b9dcb786f8e3a610;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h130b1d5f78a6277cd2b916004a26421;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12dcd68b08f938b99589764defe127b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h123b5d2c93ce1503f333da460cfe6d5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ccfbc74bda2959f976781882d699a0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c139658631668004c6aecb8b72c1e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18cc044adc95f029d8c16cde0ffe6b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1708721c59b988a8f851c5dba0cbe63;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha61c259d47a77b457a289e8cde816c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9dba9491227c7a6441aad88c47064d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13aaa4e1dec096eb62e96dfe699cf5f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h161378d67fe7e936ab0c9b85058ecb3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a68b78ec6ab4c67d9ba341d89ec60;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h90c8f7c43c3b40c65a143019556ea0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h24843aecdcf5eb9b5aba43f8e1f4c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd78be980ef3bed50560f8b24c33112;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc2ec955b2d0a386c73e55039ef0672;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6cde9f6b7625f8fe9b005b8d347e34;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h58de6e73e79431811bf6bd09341f61;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4ccbada06ce9608e997588b6dfacc2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf1c7a99913687e08d87c3d3c43dc48;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a7eb5ee7aa6dbb66abca1f3c7c0d75;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be25ed46f759bf22d9c947bd50defe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12b4ddb14514ff8c4f6d2d67f2c07eb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1160331752fe08a5e1a22425ee7b9a5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec6f52e4397927ede9f03f06dfe2a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hba473b2a11852d8b35d9ae09c3580c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1313f2ff09c98bd99242b424f81f605;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h121eb19e54156700ec1662065f6dda1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d63c4df3100405394fdf043c4886fd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10034afff6c46c539b315e14d71002f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a0484fa381448273779dc00c78ab4b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h69ac612fb591dc2cc7ca4fe93f9fbc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc77d7f573c9e057f1309b8a9caa574;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10162dd9da4b93495d3cdc58df8908f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6566cac650dfd8ae65970836aad09d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dc18fc7f34425a9922f5c24eb8dee7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h54d1bbf5bae13af1b1fe32cf1512e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha2e14b1d2be6a7bbb8580825fa3d41;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ab5018cc6c90f61406daad18eff91f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h35771730734718127e231a669e6c3f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h63a55c13f2f71af253958dc3ca4b02;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'had9157ed864032ac5fdaee5526262b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8c6cb39f849ed777d19a5a302b6f77;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7b19573a352f72c5a23b27752c46c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1399d69eea20d5ddb8082f21699f42e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5129f452a49d1a5997854519f2277;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h911e323297944260c080d209c29414;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h26e1c3c0ba392b68d826483af8f2c5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160a7fb13e37bb139ebc9023851c59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h23cc67c962fc0d87448dc2b32373ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce8a5b6689c40a956c43cfb69e771e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfc7180bfbbc336f83d0054a0abb65f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14a2b9c30bd48c3079081a818a0fffa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e1ae5b683e9ec574017408a0519fa8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f6e0b521ba1063056d62ccb350996c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd89f747462a97d00017c9f57f20cf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d8ed8dacdfcfd2bc85a94843b6a1f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9af5caa8d4ed6a4f963d16bffccb91;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4df5c2ff74cdb43c025ba1a5520cac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8b38560b9cf0d7c0cca4e44ddaaea7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4d7188e603e76dad4d8e2200c20887;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'habf4543fa4f466c162d4fa6c1cf95f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c81b30eb7f3919fc616cc363becd95;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8a2b707a4790be86442cfa8fdf4b92;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h194d12e3d8cc7bdc45ebfd5a74ced7f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd734f92a8e715e82e52c600f795284;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h965212836e38a491f1d6ae52835d93;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d613a664a05fc82dcc37609c7024c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a08249fe5774364b30dcb79d7f040c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h626e8256dd191e3545da17dfd33901;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf82dfd6c0cb95d3c9fb6a4b49e6a09;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h189b6a6f06684b2ded27a750fba2f48;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd306507c8626783ad490333f25ae61;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c4fc322a8e52ecf0a00f370cd023ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1472af291ae19e49df2d7fbd8215ef8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f678185a8d112445aaed721adcf11;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2d7f00d3fb140520a1227fc3ae81a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75654a0628121c04af03485cbc9f7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a25a1ac13ebca03d76aa6911c6243;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h167a24adafc59dcfd99f39695faaffe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heb1c7cb9e8f3fc3d0a3e0bdda299d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h180a51376fb0b13d3d4ab5cb21db6c2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18ce82758b30bd4ddaa472f94969805;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h133192b439ec1154dfe31ed99348a9c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15fca53551e27e5229ec6318138aa63;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc37620c1f73ce5452e4a51fde0959b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2ef9b3e37222e6e2d1fe638f18cc42;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c1147515afca93f276a154fd90969;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h143d430c6daadc810f22dcc939d750d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha20202d4fe56bafd5bd4681e3cf1a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h137c27b81fceff68bc45cb71c4dea95;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15912c7a2910aa4762017932fc7f503;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4618347542d82d64185d304cebaec7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c92c980f728f126c4c75e79208fdb0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c1c6758b129fd8ce0f057287dd0543;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11060eb17a5428322ad855943945d1f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf49fa95386510115531fea5c4a471f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdde8027523e0c644bb1eed2631e7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha9d5a7afb55875d8b3e62354ad4747;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5275e0d953521245e98b58be6bc6f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h136105d054e449c5e74ac5aeea807c9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h647364f0ad3012455a4a5a56fcde0a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7b450aa185cc3fc6cb82e2efea5c1d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h122fff0062adef4c0a2c3b15742b323;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h29a48b7dc1655231a595f4066d07af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h364c375db0de5f736947c8c182a49c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15141126aeca3342bf73d406d53ba6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'had4e6591733f1c90c467a041b7be89;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f5e6cdc7f8446d00ea6042967f385d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5bad255344be487d25c786461760f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16ad1419f558651e4ff290c20f25a47;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13389c03dd103a83190e091166fd0b7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12df7a5b815f87c38c6914428be0e7e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb97bf063e49751c95fcef75da30f5b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2983445541db724095fca2c60f1c68;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb6bf4ed77cce400520467803fd9080;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15184e4280c8aedfa902fd5ad61136d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a8563de1cf49e289a1fe10a0d8bcda;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1885babadb13eac71049cdacb6d9cfb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1701a0895d19f25b3afe4170e835b89;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14656fdfb005e5e0ce8573cd0f13aac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18013b6c122cd2614387e3135de954d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h194462d515f21422bb9e34de8d2c03a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h193837d8178a6bfb7ba4d0d65872946;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h169a22a6e3d0a3e2a07a969beac2592;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19df3f1009ee6c627c2541513657c16;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h101c022033e12d07d6a4ed9734eb609;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4269e9439fd128485b0cdabd583782;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b157dca231897706ae304905eff70e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf650dfa36cf94b885250a1e3231c58;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15bda5181917c68082dc2a7bb6625e2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a2c0551f0f213b3634523617140ef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1737a82816f1dad3c4675a0a016b210;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eefa9859d8598338beb6906f5dc487;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ad86528f72cea115674576c984fdf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e7824a51d469dc99b19dd3734645c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcc2e53cd3416c8b6f64989fa3a7c38;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d3a4fd234176c98535174b959847b5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc7e78afd8094556902c1419c227ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14795182a1df15a8c06887de480a1e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18c1f5d4040eca4b072dd396d8c00e0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15f9ca5c37955592d4bb7a470971a1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4fa7619af7512b23988d6b5e7b25b7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6d4542ecebae6ffcd41096d402770d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h95b824bb615f1e32474d0a8aab08af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14b1f3884e60cbb787639df4d9b4493;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d98fb7ef5a2e3fb2fd295cd18c175;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5c5532694f75fef9a241a37484c9e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ab19a78c1b0840b83d2b7e6cd18089;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb9c748eec22784fb85efe06cfaa8e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h954d2a6e0d6604ca0275ab60c5055a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e86d853c2dfe3982f04b38f968e30;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9905b45473f105269038c55bac2f42;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb20d33304bcd813c1e651c26a8498c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hae6b84dc2a9e628bb4ed90fac62c4b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4e601b107927fdb2d9a139711e13bc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h185ffa072853691ab6659a39b7c328a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dadbca2e06e4fd5a2f66e2230d71e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h352d119009bec68819f026cec79e59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b14f7128335efeb5679f2df5111601;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e9dc2b86731945b6a9522f45aa77b0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11743bc1350b6f2ede1c96eb6991a67;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13fca74cf5cdd2c289262b6f942205d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd031ab7b0a9110c9d5126a3ff85165;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h112474eae5af86b489923c4cf9bacab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h182db73cc8b307201e1eb6d28f58906;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h26115a58afb68e7cdd024d41d9dcc7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h81cbe5e637716667152a2ca39fc1f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h147089cda53457f62bd568ce444bba3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2d9c92ebc27fc8512e3a864335187f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h426ec8501109087ba0fa5d1dfd5682;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h140f908ce2e84032d020a30f50232c0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfaac35699a6746bb792a46c2c84d6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h189efa01b5bc3c2c911a89e7c96ddd8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h104d3c9853d39cfc169591040636f1e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h815b86d4050f125faaf26b4a9690ec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd0af10fd4e8a30db40d1d1d4855e59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e3885b0cf460e50b1a7e451a86b645;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc000f3b271689efd1095ebd7eec65d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6b835f1e12aa37cad00c063eb2f02;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h31ef3a6cfd59394ab0cb797a49d238;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbceebe63b851ee6913ff13f4d08faa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5c2d682c60b8b324660f4a916626ec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h65580aab5e72803796b3002e2004ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1317401b1f7b5b2117c79ed41d4ffd9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d982b370b68712956b26c1e080a533;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d18983bb004a5646102ffa859e51c1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9aa9f01a64034c80ec9fe31fd79037;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15bb090d59e88a5d8151297f0abe540;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16a929faccc2440c8bf86b4c454f7a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3756271d116d211000a238f0dfe3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h30c281fdae45a77de48fab47e8476;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h70336107de69762b70e77c1264a046;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a521e60166ce2fa32d1b83ea7e094e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h483e73e7d7bf3b4a561a903711df94;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h293df233deca757f4dd48fc381bcac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a4e20a8586b5644dc73d73c3a12e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2852e95732589f44a80c1461a125ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18b3801b5723e0e315b1190e972877b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h175fdc2741a955a1a94eb2fef24a6c8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c9f3950cb9890f9ac85356b532aba2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h146e152a8fd29518a78004cf435f658;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1666186e018e09804e69d424579dd9a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4e83fee5caaac0c644848b02381fb5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h234deb4f9ff35064743dbc1331b4f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15be815f58adbd4e2a5b9da05669700;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12b00d4548f1cb724cee60a42de4b83;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13315445b4ba189e62e8de14487dc11;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1008ca810f75497545f8d05e65aada1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h542109eebb5aa3bdf3aa1aaebcf20a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h383d519c1d179eb164715f59589ad5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1239f27335bf1bb4a9781f16d541bc4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd58674dc7e90bf56999435f2b9c10b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dec4708e4e6235703fc62c4866095e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h198a85cf615bdfa1faa38d8b526b1ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he5d85e8c96e57d67f574c4b15ff385;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h379ab29f4112dc1a3acbcfd3eeb233;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h391f055478725880c732915ad9406e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h449196ed7a8ec200c366329c9fe85a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14d74115458efafa800ec6b029616b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac6d04deb76d0314c7ef7d691c00b1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h458e8a8497cf93e95e9c5befdfdcb8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd4a5d5de04864248620a4139f799e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1559e9c97d64d50e4b30e38aa69feb7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h355f449f0d58bb68158b2086b5650;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e1bd03d600d0c2c94ccf2dc8884e7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dba1dbceed05852d74823df8279b40;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13175ce3f45bb7dab2928f64dd76d9f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd585c49cae111d5783d301c7d53a95;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha806e7183bc0f3d3c0ff7972bb926f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hda6ab5cacda130e816a0c5aca7f5a0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13154454ce117bbd841bc53c119bf62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h149a2ccb7841390d59d70fa89c3ce24;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbe9dcf96990f44f34aaa19852781c9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h481869461c915483a2e341cc93759b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h183fd4f7b0911c53d0d88179c25e36e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1359a84c38dc30de046db47e0e24da6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h114f49f8f66d647c9f022b240e3e650;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h92ba331693f5c0f3acde19058da5b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160c1d35dadc14c12a378eb94085b2a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf3917c2b41851fcc67c0f57c2c8d09;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111d1ea712c11c6cac0293380814607;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ebb8fe99d021ac31b54c86b1f3316;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd4bcc05d8c1ea585e88db24663689a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd0766bcbc0e7914ad130094a728689;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h38caa184f26eedc473a5be522f08b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17a855f64b1c3da740295089b128a08;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f6068d320d28423bb68da158b26e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h65276b6e35f6528d1a00da873ec3cf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h34f52f71177411b2fc52403dc4b69c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h178ed601c68e9c9788b6088da2752fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1968ab6cfdc8c80704241d7d05396ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h918f720aebbb1df4a5332c6e9813cb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c11a13648ca8f7bb4a030aba11505;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d14a1204d0bfd8967f912b3ad905f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h490c0020372a936da4f4bccef87a3f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a54180bb989e59f0cdaf187607b9ca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3accd2463e76bc0f43a172c62ae1e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bfdc863d1e4f864e11c10c9edef235;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c28e39fbed20954411e36ebce84080;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2c0410f2d7a916c4deb1637b28e2e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h152edfd939f527605e88ad87fe342bc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13be16c1cc68dc8eaa6713a8188e467;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h59b501c2f8fd768862d6c776c4eac4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18f922d3cf29a0673790397760a3676;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h150fb4bdaf77224ea72df60edb64b1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h84c2533dd530768a7c405c5c05c7c9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f019adc3c92bdfd8a20b8788fff80d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcef39e8e592932d0923bc5aa075b4b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d61ccd69c98883e563a2f1dd350b79;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h56525b784843938d749e08f49586af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f8c5720f74021c364d99c06e69d77f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c565fca7d11fa53c1e3c717268d42e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdba95e4caf479a9859d31f927c4cc5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h20b0a4a9bba80915302bad539be65e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c88f80bb5575372c4a574626d9bcd0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd260e2339f2b7902cb063cd1d8449;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfbc8fabc45636bc2c8921061458f67;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e1d685c18545845b93f0e28adbf90c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h131987447b9aba03e13be854425e92;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18b4a860dc6871557ade37f1351cbd5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha204df22d078b490296be5b0f45591;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb09abbbd4cfb6d2bbe216e1a1d43c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdf5c0eba6c6426da6fda545df9f1bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ea00ed72bc1bbe65c106a24532c0d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9fa38b4a4cb79edcd9ced17c1a0cd0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h168d7268a65260a7cad4d1d91dcc93d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdfc6ccaaf85ceead00910be959d78b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4fe2685f1808719fa212c1f3642b2d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11735e4d24b8e4461592794ab1564b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h65fa31236b07036aa873ae82bfd664;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11211e4caef9a2fb2ec8ac08016c47e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d96acdb04549bb340a77a04db146e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h824fd8cbed570248c0aecf7bc26793;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a3ad500627a5551a0d694a700c66;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h93fc50ca9682c4d4dd2a58c3b99ee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f3cda4de095908834cdb090c1da74;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c83b2eae3484385b871df45411723;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb97c898bcced20b89181c77fb75ace;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfbf5265f2862497e25241330b27d5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5f05e0dab9c7ba540c36e37794aa89;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he39271bbe95449c36deec117cdfd01;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c051d18dcf9f7d3e9985115d6b8fd2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ea46a625b4e75dd6256d32ea7b56fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15837277b8c9ede3cd5aae9f5b844be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h381272a6aeb3f97ac00544381d4c83;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12634ab92f75ceb0f62703b0d754f89;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1034269c3803ea1d86516f20b9f5400;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h60738dde61e36caff139d40c9a5c38;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h95d128597ea7e9858947472c2dff95;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h816517cbb37a66fdb3632127a0dc9f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf580a6e0d69b4cf0c70e2d60e41d73;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe0bf2009ada19fc002ce3968b0d7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfcd76194d69cc14f41eb232f82bcd5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6349fdb4278b88a976a7c596c2179f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a1edb05662de8445a558aeb031787;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f65b5dbe248ae7c76597b65f95bbb0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14c87c3060b253687e1093c36d4cd6e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11f9832beba8383138b71a0da8a0a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1940ed570f49f620e9b992cbb406a37;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3fe09657a1c3007b1287ef9ed6b4d9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13dc0df878a69d26b69f5684e6bb13f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h39ffb8d18d834f33c49ddcd11431ca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haaeb3549ea01eb5a6150482acb5cbf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he9770498b87951736d8be25c69f9f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc259d9303bedebdb7f527a5c20571;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14dcb5ec9ec9b69a9a301ea153316cb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cb5df086e9c57ca0f5a14075e19b8c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b1a43475cfc73f280826013ba7730a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10e9e3ac8acfe6c93e36513cf789150;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17617e71e46b41d5c99ac81df35891c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h98d2b1c067786bde9ec606b7b897ca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf79ea8ecd9ad60aa7b6d0fe54c267b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13d966062d05ca803f6a8aee401fdc3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11a8d488f419235dad3e2514c4878a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h137f9eff4cfe91c33f96339723fcb87;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb6b1e2cac8d8afd9be35508803542c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h193e08c3fe63b835e8c6f09e72c798b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e98657d3debb7ffbdf94517908261a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h119d70989d1d526066b345487b7f244;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha631541e6b3834b2834529cc7c2728;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d35b903ee0db68af621d35cfb9eed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h82bfc8dd5b49fc2127eb824261bd3d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dad7985c2b4c62b8f40f150c935eb2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd8d1517ead4f7df9598a5aa45463b1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h35354c8f793db8874d859a7e7398a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b6454d45677cca91d6f2eca92936f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d9d2950fb2989969b0ee3b2ed2dfd5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h156a6214739ddde9787e8382f331a97;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7d88a450754a429adc2dd54026992d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e97378b5297b12a70016a1fd04447b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124d99954a22bac4284157a0d29890b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h102a24d5b80325db5e14ff6142710e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h61988f778cbddda572972c194aed95;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcd4505fe3b4f7b5f403adcdbcbec79;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5d3970440d318180bd8c735431bcfb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7524452dba8eb9c694c76f92140c1f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16091f50d1937f017ffe152556c6faa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc9b34ecd0ce560cc3b4961fbe191b3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb73b6c119abce70f881b542fb66f71;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h22c1917401574acf392e8335a2dfe4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf6ee523ac0bb78c32f5771b187f050;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12fe64d23df40147e216a61eb2dfd88;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf1d656d0e11829ba85bd9423630f3e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb9e5565da8357874792302c5bb6172;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9fd624ea37952bc0822b0768a82651;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e130273bdf6ee05cb6b5f4729c39d9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4da942015f5109540d2023ca2a4198;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1177b0870ceaf0822f62b59e57b5bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h26026f1cb2a63c9d5147b83f2bb9f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf10d03893d4f2ea6bccbfae53d1ad5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h644ea74a43e32b93450f732ac3516b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac7381720376470d7da2523c0fe0f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cf510af629bf49827d8c7ee04ebaf2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h68e76fdf0d5ba9b257931e2aa33889;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cdb8120d90e9cceb6eef06be79d14f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f3d245e2a57e9caf814715439d771;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1992b73d369a3cf10b77fc96984abaa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h786683ca0330d1c21c60f2e9ba6d29;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5bda0dd7212149246b67354c1108d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1500b7fe09949b436ee98de0120f123;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c52bd9d97ebb752e6294784613f6cf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aa3c93af7d3261ca7956ba15755437;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fed62557a5092c25ab1637a28b11a1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12b8643c713c9099952d48d215627ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb1483c4bab0e14a43e21e08acde403;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1029021e367ff87d9df9eb343a6b22b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4871224198f1abb18c0857d197b8ed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hefa2c885b3e890290c21bcc6069bfc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18dcd40360d49ece5e18d1965c68e2b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2ba6aa6e89511003f90ff3458d6a56;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157bb1f9ae638644e8dd050715dffa8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb1324200c8e0e2c3090c5d71dc325;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h147db0284e7a253f0b09eace16adc62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8efc831848647ac524fe29f1203ecb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7fdf1a9f4c5ed51a877dffbc79fe23;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7703bbacd26d3a3201beb9e6f9b265;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1434752cd05e11829cb8b587ca82b5d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13bc14f366e2f30fac44e16dd02fdf9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h509a533d6f95ae7d94fbc1433fad6a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43d67ef0953da0fe6710bf741ec2c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b0c5893bd9dc5fa9d7c12ef1f5cb9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h869880c410808d540a35f8d8ce6ad5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h188ae127a2365c17adae41eef81835f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160bbf925a47a0e0a1692a130dc3763;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7735c4e48ac93827d5a39729d96a44;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd4886d103da94b9b8b43b0fd25f10d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b21f80e3a6aac3889ed9a1b1a5d3d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a2e97f9f374d0c16029e1d9d5c38b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h184fa45123372aecd5d9ea1264ea304;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d60a0f13a199a19119f0fd2468ee50;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac076f0180a76df949575e35ec34e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc8fbf181cd7ba26c1b115a709aff86;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc8317c4e36452cf1765f83e8b5b56e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a120a9d594cb9e9ef94bd043378ca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd3162054d0210734e2568ddb9289e2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc2775bd6a30d06e8b3fc1d4ae9b53;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1681ce11134d08197d6b6701cde1073;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c00399c3af1ddaf485944cbf0bb9e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hef857ea93ac27e712d36dea77229dd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5bc58a86175a756b85fd8c2aeb66e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f2ce411c94f651a9058c8954beac5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc22cc820c3c6f227a62697ae39dc65;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hea8ee3b2a966329cc9f634cea0d849;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a0077f23ea4bd471f7ea2fac197f6f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h207f3568c06f8f0f981096cbd1c857;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f8094d127bfc7ff3d9d4e1569842e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ee8d8a32ae9f9467cc2f1bb1d8e8f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10fe0abc3e300a80cafc8baa0a4a3ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h166c8e76e583a238df38cd37283fd7a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h48cb0bce2a299a3bbeef31527f5bdb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75ea44c4a4c29211714d08fd58d169;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf98e1dbab4c815e7bf55806cf6ba98;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1306cd030ccafd892ef7c9bb09766f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4c474fbe9f969a55cc08cf58eefa54;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d6b0d60b7f9b811a47b8fbbf1e9f0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ec439f9d555c7df22595b0774fbad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h31d99ba0125e7a125d513ebb59313e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h130b6aabffb1a56c439b6486716dbcd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ad6791839415375c452dbc885c7d89;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ab64f09d7380571d42e7eab9830761;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h65d901d1f571c1d04b7bd800fd2ca1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ee2794994467c58f64de7c5e963cf8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1674b2b91b34fdb43cf2153319e1e2a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5ef6617bfbd2ee36044414068c6bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae621ca329ffc6ffc94194c9dc06bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9eeacedff59e6e95d38959ef5928d7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha8a64539277752852f6b774f88246e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he73316fc639a2412ee5c1ed9142424;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1004037d1fa8b45ee30ef8d533a1d88;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e92221ad4010a4e5da8cfc3b650b36;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197bbe5eae4dc4f9199807fa88aee44;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c577b1c13c3ec85a454bcd3010a812;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13f75b82cd74ebe9b4f3b051fb9e9cb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha9f28c5ca980c249e62c7a09f39cc6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a995e78f642832bb70f31fbc6c7cb2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138af39f0ed002f26b114385a1b5498;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbc2a9eb06f3b5b90952bce2f461ef5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd83e46496d8942e4805c87df1ebbed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heb0bf9dce03ad7dfeb75b1d379d35d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heea437a86b2a683308f3f2ed43e07e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b03aaaa01ce2e25ee9294a619c595;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f0d6cc410f2eb624d4e278ca629af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1303a2b0c4cf511dacb6c3e34a5384e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h47235746a0656451bf5064e4de71be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d3a22bdecb58727144b4e704d8af32;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h96bc9116ca4adde49c360d29ac15be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha058d4e838ddbceb7d364233dee108;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2ce0c029a63fb5d5f51b3b525b16de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb5cf6b1b16b86586315e12b0d845d8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc871f7e0eedc74b2fa161a2c636b42;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcec16659171c648eb5655aa3d9a01a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde1e482e962f1f83cb31cafd3abb42;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b0acf0178c699aafc06d6ec006861b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd6e066963d31d9844e541bdb973798;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ed7a1a90d900d41a0c20b8010577b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h195acc58f4632047440305aafe3732a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1530e62d049b25b3bf80fb0963f1132;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e2d02cbc78c1758aafe1c88735fc8c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h894dd44de3dbca71d3ccc51be55a3d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha5c075dd54ba32f5cf9a6e52257999;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c809c84b17da414bb03bd48fe18fa5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h30ea9771b3bcbec2fbf3221c2c39b0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5dc638335109280fc0bb1af4a81a33;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8e03fc33de852f88c713e7dc2c9950;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10861f641b8ffbe4f3cb17c72a789ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f3159deda633fa812531c787643b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h25888394ed26e10cf8d5341909943f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h65b933669a165e6e873e5c6958996c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16a90c7ae3b53250d4102e491080e91;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h350fdd9aece858fa0541b76be62e6d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1008ed9dfbc79fcb8ee3d8557bcc0b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d3f6ae98b313cbdda0111164253cb2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18d958315ba200c5b6cb6cee79fa8bc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8356600780ea07d7dc42c9dc195914;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a3463a0905e59aeceeaf3f261ee79;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5eba8313118269419dec011bde9a53;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h191ce8785f7d1d3e531e22beb97c8cb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h242c5d4d021eaa07ebe02df5c294fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8993f57662778651a5179701a14516;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h126c24b787084afbe492fed3cee311d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10f2f244640743301211ace539a38a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5314f02d8e46d6843980d7cb67d3c2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12968acf1fb2c32a35388d8b6bc0f0b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e3eb4e7e6e434c5f8a4e864867a52d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h81d4998c1891601260fc0651e19653;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16f7184c4931d4e2dc1fcde648ec2eb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a8c0a3536aab9fd81cabec7890123;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1612b339656cfdd19aa86e7a7bd3bf3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3e252c6848606bd597966f15e897ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f5da9d6cb8305623d7b82f347410fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h54288dc53f6a17a3388b237527069a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14c595a84e0e6de991d6c75952e3724;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec7d69f2f3f973f0287d4f5c7ce3cb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2ab277021eab761be7bbc91fcb3e6d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c758738f3be70355249c658662e777;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df599cfb90bc32cec535213016e440;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cf601216eaeba43ee999e457717b35;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf269e97abf5e127fe569fa47db6628;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h519bf8c6d8759528b1659980a0a52f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h158412d3ad2a647b8323a8efd624538;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b612218b350a58eaeddd043e25a63;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3818322388b1556bb19950a65fb8c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h57634b0bd1d51c90aec6794be371e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6329cf9fb1ce8902c0d5d84f3f06f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f786859cdf3c49da9bb0496c4278f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6c877bf67e03bd3a20e2c752426a2b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12dcf7e2fcdccb3ed869cdb1d206e9f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18fcff80425043ce533a5464fd12251;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h36f0dee377ec5cc119d10f2746a501;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17de658e379a8adcb39d03922c4ca4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h39d8a13949227d15b53f079b3c9523;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h56d95d8f16c9f271a2362f7afb682;
        #1
        $finish();
    end
endmodule
