module compressor2_1_54_16_shiftregister(input clk, input in_data0, input in_data1, input in_data2, input in_data3, input in_data4, input in_data5, input in_data6, input in_data7, input in_data8, input in_data9, input in_data10, input in_data11, input in_data12, input in_data13, input in_data14, input in_data15, input in_data16, input in_data17, input in_data18, input in_data19, input in_data20, input in_data21, input in_data22, input in_data23, input in_data24, input in_data25, input in_data26, input in_data27, input in_data28, input in_data29, input in_data30, input in_data31, input in_data32, input in_data33, input in_data34, input in_data35, input in_data36, input in_data37, input in_data38, input in_data39, input in_data40, input in_data41, input in_data42, input in_data43, input in_data44, input in_data45, input in_data46, input in_data47, input in_data48, input in_data49, input in_data50, input in_data51, input in_data52, input in_data53, output [21:0]dst);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    compressor2_1_54_16 compressor2_1_54_16(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .src32(src32), .src33(src33), .src34(src34), .src35(src35), .src36(src36), .src37(src37), .src38(src38), .src39(src39), .src40(src40), .src41(src41), .src42(src42), .src43(src43), .src44(src44), .src45(src45), .src46(src46), .src47(src47), .src48(src48), .src49(src49), .src50(src50), .src51(src51), .src52(src52), .src53(src53), .dst(dst));
    initial begin
        src0 <= 0;
        src1 <= 0;
        src2 <= 0;
        src3 <= 0;
        src4 <= 0;
        src5 <= 0;
        src6 <= 0;
        src7 <= 0;
        src8 <= 0;
        src9 <= 0;
        src10 <= 0;
        src11 <= 0;
        src12 <= 0;
        src13 <= 0;
        src14 <= 0;
        src15 <= 0;
        src16 <= 0;
        src17 <= 0;
        src18 <= 0;
        src19 <= 0;
        src20 <= 0;
        src21 <= 0;
        src22 <= 0;
        src23 <= 0;
        src24 <= 0;
        src25 <= 0;
        src26 <= 0;
        src27 <= 0;
        src28 <= 0;
        src29 <= 0;
        src30 <= 0;
        src31 <= 0;
        src32 <= 0;
        src33 <= 0;
        src34 <= 0;
        src35 <= 0;
        src36 <= 0;
        src37 <= 0;
        src38 <= 0;
        src39 <= 0;
        src40 <= 0;
        src41 <= 0;
        src42 <= 0;
        src43 <= 0;
        src44 <= 0;
        src45 <= 0;
        src46 <= 0;
        src47 <= 0;
        src48 <= 0;
        src49 <= 0;
        src50 <= 0;
        src51 <= 0;
        src52 <= 0;
        src53 <= 0;
    end
    always @(posedge clk) begin
        src0 <= {src0[14:0], in_data0};
        src1 <= {src1[14:0], in_data1};
        src2 <= {src2[14:0], in_data2};
        src3 <= {src3[14:0], in_data3};
        src4 <= {src4[14:0], in_data4};
        src5 <= {src5[14:0], in_data5};
        src6 <= {src6[14:0], in_data6};
        src7 <= {src7[14:0], in_data7};
        src8 <= {src8[14:0], in_data8};
        src9 <= {src9[14:0], in_data9};
        src10 <= {src10[14:0], in_data10};
        src11 <= {src11[14:0], in_data11};
        src12 <= {src12[14:0], in_data12};
        src13 <= {src13[14:0], in_data13};
        src14 <= {src14[14:0], in_data14};
        src15 <= {src15[14:0], in_data15};
        src16 <= {src16[14:0], in_data16};
        src17 <= {src17[14:0], in_data17};
        src18 <= {src18[14:0], in_data18};
        src19 <= {src19[14:0], in_data19};
        src20 <= {src20[14:0], in_data20};
        src21 <= {src21[14:0], in_data21};
        src22 <= {src22[14:0], in_data22};
        src23 <= {src23[14:0], in_data23};
        src24 <= {src24[14:0], in_data24};
        src25 <= {src25[14:0], in_data25};
        src26 <= {src26[14:0], in_data26};
        src27 <= {src27[14:0], in_data27};
        src28 <= {src28[14:0], in_data28};
        src29 <= {src29[14:0], in_data29};
        src30 <= {src30[14:0], in_data30};
        src31 <= {src31[14:0], in_data31};
        src32 <= {src32[14:0], in_data32};
        src33 <= {src33[14:0], in_data33};
        src34 <= {src34[14:0], in_data34};
        src35 <= {src35[14:0], in_data35};
        src36 <= {src36[14:0], in_data36};
        src37 <= {src37[14:0], in_data37};
        src38 <= {src38[14:0], in_data38};
        src39 <= {src39[14:0], in_data39};
        src40 <= {src40[14:0], in_data40};
        src41 <= {src41[14:0], in_data41};
        src42 <= {src42[14:0], in_data42};
        src43 <= {src43[14:0], in_data43};
        src44 <= {src44[14:0], in_data44};
        src45 <= {src45[14:0], in_data45};
        src46 <= {src46[14:0], in_data46};
        src47 <= {src47[14:0], in_data47};
        src48 <= {src48[14:0], in_data48};
        src49 <= {src49[14:0], in_data49};
        src50 <= {src50[14:0], in_data50};
        src51 <= {src51[14:0], in_data51};
        src52 <= {src52[14:0], in_data52};
        src53 <= {src53[14:0], in_data53};
    end
endmodule

module compressor2_1_54_16(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    input [15:0]src16,
    input [15:0]src17,
    input [15:0]src18,
    input [15:0]src19,
    input [15:0]src20,
    input [15:0]src21,
    input [15:0]src22,
    input [15:0]src23,
    input [15:0]src24,
    input [15:0]src25,
    input [15:0]src26,
    input [15:0]src27,
    input [15:0]src28,
    input [15:0]src29,
    input [15:0]src30,
    input [15:0]src31,
    input [15:0]src32,
    input [15:0]src33,
    input [15:0]src34,
    input [15:0]src35,
    input [15:0]src36,
    input [15:0]src37,
    input [15:0]src38,
    input [15:0]src39,
    input [15:0]src40,
    input [15:0]src41,
    input [15:0]src42,
    input [15:0]src43,
    input [15:0]src44,
    input [15:0]src45,
    input [15:0]src46,
    input [15:0]src47,
    input [15:0]src48,
    input [15:0]src49,
    input [15:0]src50,
    input [15:0]src51,
    input [15:0]src52,
    input [15:0]src53,
    output [21:0]dst);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [0:0] comp_out20;
    wire [1:0] comp_out21;
    wire [22:0] out;
    compressor compressor_inst(
        .src0({src53[0], src52[0], src51[0], src50[0], src49[0], src48[0], src47[0], src46[0], src45[0], src44[0], src43[0], src42[0], src41[0], src40[0], src39[0], src38[0], src37[0], src36[0], src35[0], src34[0], src33[0], src32[0], src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}),
        .src1({src53[1], src52[1], src51[1], src50[1], src49[1], src48[1], src47[1], src46[1], src45[1], src44[1], src43[1], src42[1], src41[1], src40[1], src39[1], src38[1], src37[1], src36[1], src35[1], src34[1], src33[1], src32[1], src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}),
        .src2({src53[2], src52[2], src51[2], src50[2], src49[2], src48[2], src47[2], src46[2], src45[2], src44[2], src43[2], src42[2], src41[2], src40[2], src39[2], src38[2], src37[2], src36[2], src35[2], src34[2], src33[2], src32[2], src31[2], src30[2], src29[2], src28[2], src27[2], src26[2], src25[2], src24[2], src23[2], src22[2], src21[2], src20[2], src19[2], src18[2], src17[2], src16[2], src15[2], src14[2], src13[2], src12[2], src11[2], src10[2], src9[2], src8[2], src7[2], src6[2], src5[2], src4[2], src3[2], src2[2], src1[2], src0[2]}),
        .src3({src53[3], src52[3], src51[3], src50[3], src49[3], src48[3], src47[3], src46[3], src45[3], src44[3], src43[3], src42[3], src41[3], src40[3], src39[3], src38[3], src37[3], src36[3], src35[3], src34[3], src33[3], src32[3], src31[3], src30[3], src29[3], src28[3], src27[3], src26[3], src25[3], src24[3], src23[3], src22[3], src21[3], src20[3], src19[3], src18[3], src17[3], src16[3], src15[3], src14[3], src13[3], src12[3], src11[3], src10[3], src9[3], src8[3], src7[3], src6[3], src5[3], src4[3], src3[3], src2[3], src1[3], src0[3]}),
        .src4({src53[4], src52[4], src51[4], src50[4], src49[4], src48[4], src47[4], src46[4], src45[4], src44[4], src43[4], src42[4], src41[4], src40[4], src39[4], src38[4], src37[4], src36[4], src35[4], src34[4], src33[4], src32[4], src31[4], src30[4], src29[4], src28[4], src27[4], src26[4], src25[4], src24[4], src23[4], src22[4], src21[4], src20[4], src19[4], src18[4], src17[4], src16[4], src15[4], src14[4], src13[4], src12[4], src11[4], src10[4], src9[4], src8[4], src7[4], src6[4], src5[4], src4[4], src3[4], src2[4], src1[4], src0[4]}),
        .src5({src53[5], src52[5], src51[5], src50[5], src49[5], src48[5], src47[5], src46[5], src45[5], src44[5], src43[5], src42[5], src41[5], src40[5], src39[5], src38[5], src37[5], src36[5], src35[5], src34[5], src33[5], src32[5], src31[5], src30[5], src29[5], src28[5], src27[5], src26[5], src25[5], src24[5], src23[5], src22[5], src21[5], src20[5], src19[5], src18[5], src17[5], src16[5], src15[5], src14[5], src13[5], src12[5], src11[5], src10[5], src9[5], src8[5], src7[5], src6[5], src5[5], src4[5], src3[5], src2[5], src1[5], src0[5]}),
        .src6({src53[6], src52[6], src51[6], src50[6], src49[6], src48[6], src47[6], src46[6], src45[6], src44[6], src43[6], src42[6], src41[6], src40[6], src39[6], src38[6], src37[6], src36[6], src35[6], src34[6], src33[6], src32[6], src31[6], src30[6], src29[6], src28[6], src27[6], src26[6], src25[6], src24[6], src23[6], src22[6], src21[6], src20[6], src19[6], src18[6], src17[6], src16[6], src15[6], src14[6], src13[6], src12[6], src11[6], src10[6], src9[6], src8[6], src7[6], src6[6], src5[6], src4[6], src3[6], src2[6], src1[6], src0[6]}),
        .src7({src53[7], src52[7], src51[7], src50[7], src49[7], src48[7], src47[7], src46[7], src45[7], src44[7], src43[7], src42[7], src41[7], src40[7], src39[7], src38[7], src37[7], src36[7], src35[7], src34[7], src33[7], src32[7], src31[7], src30[7], src29[7], src28[7], src27[7], src26[7], src25[7], src24[7], src23[7], src22[7], src21[7], src20[7], src19[7], src18[7], src17[7], src16[7], src15[7], src14[7], src13[7], src12[7], src11[7], src10[7], src9[7], src8[7], src7[7], src6[7], src5[7], src4[7], src3[7], src2[7], src1[7], src0[7]}),
        .src8({src53[8], src52[8], src51[8], src50[8], src49[8], src48[8], src47[8], src46[8], src45[8], src44[8], src43[8], src42[8], src41[8], src40[8], src39[8], src38[8], src37[8], src36[8], src35[8], src34[8], src33[8], src32[8], src31[8], src30[8], src29[8], src28[8], src27[8], src26[8], src25[8], src24[8], src23[8], src22[8], src21[8], src20[8], src19[8], src18[8], src17[8], src16[8], src15[8], src14[8], src13[8], src12[8], src11[8], src10[8], src9[8], src8[8], src7[8], src6[8], src5[8], src4[8], src3[8], src2[8], src1[8], src0[8]}),
        .src9({src53[9], src52[9], src51[9], src50[9], src49[9], src48[9], src47[9], src46[9], src45[9], src44[9], src43[9], src42[9], src41[9], src40[9], src39[9], src38[9], src37[9], src36[9], src35[9], src34[9], src33[9], src32[9], src31[9], src30[9], src29[9], src28[9], src27[9], src26[9], src25[9], src24[9], src23[9], src22[9], src21[9], src20[9], src19[9], src18[9], src17[9], src16[9], src15[9], src14[9], src13[9], src12[9], src11[9], src10[9], src9[9], src8[9], src7[9], src6[9], src5[9], src4[9], src3[9], src2[9], src1[9], src0[9]}),
        .src10({src53[10], src52[10], src51[10], src50[10], src49[10], src48[10], src47[10], src46[10], src45[10], src44[10], src43[10], src42[10], src41[10], src40[10], src39[10], src38[10], src37[10], src36[10], src35[10], src34[10], src33[10], src32[10], src31[10], src30[10], src29[10], src28[10], src27[10], src26[10], src25[10], src24[10], src23[10], src22[10], src21[10], src20[10], src19[10], src18[10], src17[10], src16[10], src15[10], src14[10], src13[10], src12[10], src11[10], src10[10], src9[10], src8[10], src7[10], src6[10], src5[10], src4[10], src3[10], src2[10], src1[10], src0[10]}),
        .src11({src53[11], src52[11], src51[11], src50[11], src49[11], src48[11], src47[11], src46[11], src45[11], src44[11], src43[11], src42[11], src41[11], src40[11], src39[11], src38[11], src37[11], src36[11], src35[11], src34[11], src33[11], src32[11], src31[11], src30[11], src29[11], src28[11], src27[11], src26[11], src25[11], src24[11], src23[11], src22[11], src21[11], src20[11], src19[11], src18[11], src17[11], src16[11], src15[11], src14[11], src13[11], src12[11], src11[11], src10[11], src9[11], src8[11], src7[11], src6[11], src5[11], src4[11], src3[11], src2[11], src1[11], src0[11]}),
        .src12({src53[12], src52[12], src51[12], src50[12], src49[12], src48[12], src47[12], src46[12], src45[12], src44[12], src43[12], src42[12], src41[12], src40[12], src39[12], src38[12], src37[12], src36[12], src35[12], src34[12], src33[12], src32[12], src31[12], src30[12], src29[12], src28[12], src27[12], src26[12], src25[12], src24[12], src23[12], src22[12], src21[12], src20[12], src19[12], src18[12], src17[12], src16[12], src15[12], src14[12], src13[12], src12[12], src11[12], src10[12], src9[12], src8[12], src7[12], src6[12], src5[12], src4[12], src3[12], src2[12], src1[12], src0[12]}),
        .src13({src53[13], src52[13], src51[13], src50[13], src49[13], src48[13], src47[13], src46[13], src45[13], src44[13], src43[13], src42[13], src41[13], src40[13], src39[13], src38[13], src37[13], src36[13], src35[13], src34[13], src33[13], src32[13], src31[13], src30[13], src29[13], src28[13], src27[13], src26[13], src25[13], src24[13], src23[13], src22[13], src21[13], src20[13], src19[13], src18[13], src17[13], src16[13], src15[13], src14[13], src13[13], src12[13], src11[13], src10[13], src9[13], src8[13], src7[13], src6[13], src5[13], src4[13], src3[13], src2[13], src1[13], src0[13]}),
        .src14({src53[14], src52[14], src51[14], src50[14], src49[14], src48[14], src47[14], src46[14], src45[14], src44[14], src43[14], src42[14], src41[14], src40[14], src39[14], src38[14], src37[14], src36[14], src35[14], src34[14], src33[14], src32[14], src31[14], src30[14], src29[14], src28[14], src27[14], src26[14], src25[14], src24[14], src23[14], src22[14], src21[14], src20[14], src19[14], src18[14], src17[14], src16[14], src15[14], src14[14], src13[14], src12[14], src11[14], src10[14], src9[14], src8[14], src7[14], src6[14], src5[14], src4[14], src3[14], src2[14], src1[14], src0[14]}),
        .src15({src53[15], src52[15], src51[15], src50[15], src49[15], src48[15], src47[15], src46[15], src45[15], src44[15], src43[15], src42[15], src41[15], src40[15], src39[15], src38[15], src37[15], src36[15], src35[15], src34[15], src33[15], src32[15], src31[15], src30[15], src29[15], src28[15], src27[15], src26[15], src25[15], src24[15], src23[15], src22[15], src21[15], src20[15], src19[15], src18[15], src17[15], src16[15], src15[15], src14[15], src13[15], src12[15], src11[15], src10[15], src9[15], src8[15], src7[15], src6[15], src5[15], src4[15], src3[15], src2[15], src1[15], src0[15]}),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21)
    );
    rowadder2_1_22 rowadder2_1inst(
        .src0({comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({comp_out21[1], 1'h0, comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0(out)
    );
    assign dst = out[21:0];
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      input wire [53:0] src12,
      input wire [53:0] src13,
      input wire [53:0] src14,
      input wire [53:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [0:0] dst20,
      output wire [1:0] dst21);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [53:0] stage0_12;
   wire [53:0] stage0_13;
   wire [53:0] stage0_14;
   wire [53:0] stage0_15;
   wire [13:0] stage1_0;
   wire [16:0] stage1_1;
   wire [22:0] stage1_2;
   wire [17:0] stage1_3;
   wire [34:0] stage1_4;
   wire [24:0] stage1_5;
   wire [18:0] stage1_6;
   wire [18:0] stage1_7;
   wire [25:0] stage1_8;
   wire [26:0] stage1_9;
   wire [18:0] stage1_10;
   wire [17:0] stage1_11;
   wire [25:0] stage1_12;
   wire [25:0] stage1_13;
   wire [17:0] stage1_14;
   wire [23:0] stage1_15;
   wire [16:0] stage1_16;
   wire [7:0] stage1_17;
   wire [7:0] stage2_0;
   wire [2:0] stage2_1;
   wire [7:0] stage2_2;
   wire [8:0] stage2_3;
   wire [11:0] stage2_4;
   wire [9:0] stage2_5;
   wire [11:0] stage2_6;
   wire [10:0] stage2_7;
   wire [7:0] stage2_8;
   wire [11:0] stage2_9;
   wire [12:0] stage2_10;
   wire [6:0] stage2_11;
   wire [8:0] stage2_12;
   wire [10:0] stage2_13;
   wire [8:0] stage2_14;
   wire [7:0] stage2_15;
   wire [9:0] stage2_16;
   wire [6:0] stage2_17;
   wire [2:0] stage2_18;
   wire [2:0] stage2_19;
   wire [0:0] stage2_20;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [1:0] stage3_2;
   wire [5:0] stage3_3;
   wire [3:0] stage3_4;
   wire [5:0] stage3_5;
   wire [2:0] stage3_6;
   wire [5:0] stage3_7;
   wire [4:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [2:0] stage3_14;
   wire [3:0] stage3_15;
   wire [5:0] stage3_16;
   wire [3:0] stage3_17;
   wire [3:0] stage3_18;
   wire [0:0] stage3_19;
   wire [0:0] stage3_20;
   wire [0:0] stage3_21;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [0:0] stage4_20;
   wire [1:0] stage4_21;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;
   assign dst21 = stage4_21;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1406_5 gpc8 (
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3]},
      {stage0_4[0]},
      {stage1_5[0],stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8]}
   );
   gpc1406_5 gpc9 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7]},
      {stage0_4[1]},
      {stage1_5[1],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[2],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[3],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[4],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[5],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[6],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[7],stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15]}
   );
   gpc606_5 gpc16 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[8],stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16]}
   );
   gpc615_5 gpc17 (
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], 1'b0},
      {stage0_4[2]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[0],stage1_5[9],stage1_4[17],stage1_3[17]}
   );
   gpc606_5 gpc18 (
      {stage0_4[3], stage0_4[4], stage0_4[5], stage0_4[6], stage0_4[7], stage0_4[8]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[1],stage1_5[10],stage1_4[18]}
   );
   gpc606_5 gpc19 (
      {stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[2],stage1_6[2],stage1_5[11],stage1_4[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19], stage0_4[20]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[3],stage1_6[3],stage1_5[12],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[4],stage1_6[4],stage1_5[13],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[5],stage1_6[5],stage1_5[14],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[6],stage1_6[6],stage1_5[15],stage1_4[23]}
   );
   gpc615_5 gpc24 (
      {stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_5[6]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[7],stage1_6[7],stage1_5[16],stage1_4[24]}
   );
   gpc606_5 gpc25 (
      {stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[7],stage1_7[8],stage1_6[8],stage1_5[17]}
   );
   gpc606_5 gpc26 (
      {stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[8],stage1_7[9],stage1_6[9],stage1_5[18]}
   );
   gpc606_5 gpc27 (
      {stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[9],stage1_7[10],stage1_6[10],stage1_5[19]}
   );
   gpc606_5 gpc28 (
      {stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[10],stage1_7[11],stage1_6[11],stage1_5[20]}
   );
   gpc606_5 gpc29 (
      {stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[11],stage1_7[12],stage1_6[12],stage1_5[21]}
   );
   gpc606_5 gpc30 (
      {stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[12],stage1_7[13],stage1_6[13],stage1_5[22]}
   );
   gpc606_5 gpc31 (
      {stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[13],stage1_7[14],stage1_6[14],stage1_5[23]}
   );
   gpc615_5 gpc32 (
      {stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_6[42]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[14],stage1_7[15],stage1_6[15],stage1_5[24]}
   );
   gpc615_5 gpc33 (
      {stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage0_7[48]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[8],stage1_8[15],stage1_7[16],stage1_6[16]}
   );
   gpc615_5 gpc34 (
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52]},
      {stage0_7[49]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[9],stage1_8[16],stage1_7[17],stage1_6[17]}
   );
   gpc615_5 gpc35 (
      {stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53], 1'b0},
      {stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[2],stage1_9[10],stage1_8[17],stage1_7[18]}
   );
   gpc606_5 gpc36 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[1],stage1_10[3],stage1_9[11],stage1_8[18]}
   );
   gpc615_5 gpc37 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_9[6]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[2],stage1_10[4],stage1_9[12],stage1_8[19]}
   );
   gpc615_5 gpc38 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28]},
      {stage0_9[7]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[3],stage1_10[5],stage1_9[13],stage1_8[20]}
   );
   gpc615_5 gpc39 (
      {stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_9[8]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[4],stage1_10[6],stage1_9[14],stage1_8[21]}
   );
   gpc615_5 gpc40 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38]},
      {stage0_9[9]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[5],stage1_10[7],stage1_9[15],stage1_8[22]}
   );
   gpc615_5 gpc41 (
      {stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_9[10]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[6],stage1_10[8],stage1_9[16],stage1_8[23]}
   );
   gpc615_5 gpc42 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_9[11]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[7],stage1_10[9],stage1_9[17],stage1_8[24]}
   );
   gpc615_5 gpc43 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_9[12]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[8],stage1_10[10],stage1_9[18],stage1_8[25]}
   );
   gpc606_5 gpc44 (
      {stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[8],stage1_11[9],stage1_10[11],stage1_9[19]}
   );
   gpc606_5 gpc45 (
      {stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[9],stage1_11[10],stage1_10[12],stage1_9[20]}
   );
   gpc615_5 gpc46 (
      {stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage0_10[48]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[10],stage1_11[11],stage1_10[13],stage1_9[21]}
   );
   gpc615_5 gpc47 (
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34]},
      {stage0_10[49]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[11],stage1_11[12],stage1_10[14],stage1_9[22]}
   );
   gpc615_5 gpc48 (
      {stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39]},
      {stage0_10[50]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[12],stage1_11[13],stage1_10[15],stage1_9[23]}
   );
   gpc615_5 gpc49 (
      {stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44]},
      {stage0_10[51]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[13],stage1_11[14],stage1_10[16],stage1_9[24]}
   );
   gpc615_5 gpc50 (
      {stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49]},
      {stage0_10[52]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[14],stage1_11[15],stage1_10[17],stage1_9[25]}
   );
   gpc615_5 gpc51 (
      {stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53], 1'b0},
      {stage0_10[53]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[15],stage1_11[16],stage1_10[18],stage1_9[26]}
   );
   gpc606_5 gpc52 (
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[0],stage1_13[8],stage1_12[16],stage1_11[17]}
   );
   gpc606_5 gpc53 (
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[1],stage1_13[9],stage1_12[17]}
   );
   gpc606_5 gpc54 (
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[2],stage1_13[10],stage1_12[18]}
   );
   gpc606_5 gpc55 (
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[3],stage1_13[11],stage1_12[19]}
   );
   gpc606_5 gpc56 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[4],stage1_13[12],stage1_12[20]}
   );
   gpc606_5 gpc57 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[5],stage1_14[5],stage1_13[13],stage1_12[21]}
   );
   gpc606_5 gpc58 (
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[6],stage1_14[6],stage1_13[14],stage1_12[22]}
   );
   gpc606_5 gpc59 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[7],stage1_14[7],stage1_13[15],stage1_12[23]}
   );
   gpc606_5 gpc60 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[8],stage1_14[8],stage1_13[16],stage1_12[24]}
   );
   gpc606_5 gpc61 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[9],stage1_14[9],stage1_13[17],stage1_12[25]}
   );
   gpc606_5 gpc62 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[9],stage1_15[10],stage1_14[10],stage1_13[18]}
   );
   gpc606_5 gpc63 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[10],stage1_15[11],stage1_14[11],stage1_13[19]}
   );
   gpc606_5 gpc64 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[11],stage1_15[12],stage1_14[12],stage1_13[20]}
   );
   gpc606_5 gpc65 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[12],stage1_15[13],stage1_14[13],stage1_13[21]}
   );
   gpc606_5 gpc66 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[13],stage1_15[14],stage1_14[14],stage1_13[22]}
   );
   gpc606_5 gpc67 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[14],stage1_15[15],stage1_14[15],stage1_13[23]}
   );
   gpc606_5 gpc68 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[15],stage1_15[16],stage1_14[16],stage1_13[24]}
   );
   gpc606_5 gpc69 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[16],stage1_15[17],stage1_14[17],stage1_13[25]}
   );
   gpc1_1 gpc70 (
      {stage0_0[48]},
      {stage1_0[8]}
   );
   gpc1_1 gpc71 (
      {stage0_0[49]},
      {stage1_0[9]}
   );
   gpc1_1 gpc72 (
      {stage0_0[50]},
      {stage1_0[10]}
   );
   gpc1_1 gpc73 (
      {stage0_0[51]},
      {stage1_0[11]}
   );
   gpc1_1 gpc74 (
      {stage0_0[52]},
      {stage1_0[12]}
   );
   gpc1_1 gpc75 (
      {stage0_0[53]},
      {stage1_0[13]}
   );
   gpc1_1 gpc76 (
      {stage0_2[48]},
      {stage1_2[17]}
   );
   gpc1_1 gpc77 (
      {stage0_2[49]},
      {stage1_2[18]}
   );
   gpc1_1 gpc78 (
      {stage0_2[50]},
      {stage1_2[19]}
   );
   gpc1_1 gpc79 (
      {stage0_2[51]},
      {stage1_2[20]}
   );
   gpc1_1 gpc80 (
      {stage0_2[52]},
      {stage1_2[21]}
   );
   gpc1_1 gpc81 (
      {stage0_2[53]},
      {stage1_2[22]}
   );
   gpc1_1 gpc82 (
      {stage0_4[44]},
      {stage1_4[25]}
   );
   gpc1_1 gpc83 (
      {stage0_4[45]},
      {stage1_4[26]}
   );
   gpc1_1 gpc84 (
      {stage0_4[46]},
      {stage1_4[27]}
   );
   gpc1_1 gpc85 (
      {stage0_4[47]},
      {stage1_4[28]}
   );
   gpc1_1 gpc86 (
      {stage0_4[48]},
      {stage1_4[29]}
   );
   gpc1_1 gpc87 (
      {stage0_4[49]},
      {stage1_4[30]}
   );
   gpc1_1 gpc88 (
      {stage0_4[50]},
      {stage1_4[31]}
   );
   gpc1_1 gpc89 (
      {stage0_4[51]},
      {stage1_4[32]}
   );
   gpc1_1 gpc90 (
      {stage0_4[52]},
      {stage1_4[33]}
   );
   gpc1_1 gpc91 (
      {stage0_4[53]},
      {stage1_4[34]}
   );
   gpc1_1 gpc92 (
      {stage0_6[53]},
      {stage1_6[18]}
   );
   gpc1_1 gpc93 (
      {stage0_15[48]},
      {stage1_15[18]}
   );
   gpc1_1 gpc94 (
      {stage0_15[49]},
      {stage1_15[19]}
   );
   gpc1_1 gpc95 (
      {stage0_15[50]},
      {stage1_15[20]}
   );
   gpc1_1 gpc96 (
      {stage0_15[51]},
      {stage1_15[21]}
   );
   gpc1_1 gpc97 (
      {stage0_15[52]},
      {stage1_15[22]}
   );
   gpc1_1 gpc98 (
      {stage0_15[53]},
      {stage1_15[23]}
   );
   gpc1163_5 gpc99 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc100 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc101 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], 1'b0},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc102 (
      {stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3]}
   );
   gpc606_5 gpc103 (
      {stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc606_5 gpc104 (
      {stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc615_5 gpc105 (
      {stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7]},
      {stage1_4[18]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[3],stage2_5[3],stage2_4[6],stage2_3[6]}
   );
   gpc615_5 gpc106 (
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage1_4[19]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[4],stage2_5[4],stage2_4[7],stage2_3[7]}
   );
   gpc615_5 gpc107 (
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage1_4[20]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[5],stage2_5[5],stage2_4[8],stage2_3[8]}
   );
   gpc207_4 gpc108 (
      {stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27]},
      {stage1_6[0], stage1_6[1]},
      {stage2_7[3],stage2_6[6],stage2_5[6],stage2_4[9]}
   );
   gpc606_5 gpc109 (
      {stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[0],stage2_7[4],stage2_6[7],stage2_5[7],stage2_4[10]}
   );
   gpc606_5 gpc110 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[5],stage2_6[8],stage2_5[8]}
   );
   gpc615_5 gpc111 (
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage1_7[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[2],stage2_7[6],stage2_6[9]}
   );
   gpc615_5 gpc112 (
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_7[7]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[2],stage2_8[3],stage2_7[7],stage2_6[10]}
   );
   gpc615_5 gpc113 (
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_8[12]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[2],stage2_9[3],stage2_8[4],stage2_7[8]}
   );
   gpc615_5 gpc114 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage1_8[13]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[3],stage2_9[4],stage2_8[5],stage2_7[9]}
   );
   gpc606_5 gpc115 (
      {stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[2],stage2_10[4],stage2_9[5],stage2_8[6]}
   );
   gpc606_5 gpc116 (
      {stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[3],stage2_10[5],stage2_9[6],stage2_8[7]}
   );
   gpc606_5 gpc117 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[2],stage2_11[4],stage2_10[6],stage2_9[7]}
   );
   gpc606_5 gpc118 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[3],stage2_11[5],stage2_10[7],stage2_9[8]}
   );
   gpc1163_5 gpc119 (
      {stage1_10[12], stage1_10[13], stage1_10[14]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage1_12[0]},
      {stage1_13[0]},
      {stage2_14[0],stage2_13[2],stage2_12[4],stage2_11[6],stage2_10[8]}
   );
   gpc117_4 gpc120 (
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6], stage1_12[7]},
      {stage1_13[1]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[1],stage2_13[3],stage2_12[5]}
   );
   gpc606_5 gpc121 (
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[0],stage2_15[1],stage2_14[2],stage2_13[4],stage2_12[6]}
   );
   gpc606_5 gpc122 (
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage2_16[1],stage2_15[2],stage2_14[3],stage2_13[5],stage2_12[7]}
   );
   gpc606_5 gpc123 (
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], 1'b0},
      {stage2_16[2],stage2_15[3],stage2_14[4],stage2_13[6],stage2_12[8]}
   );
   gpc606_5 gpc124 (
      {stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[3],stage2_15[4],stage2_14[5],stage2_13[7]}
   );
   gpc606_5 gpc125 (
      {stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[4],stage2_15[5],stage2_14[6],stage2_13[8]}
   );
   gpc606_5 gpc126 (
      {stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[5],stage2_15[6],stage2_14[7],stage2_13[9]}
   );
   gpc606_5 gpc127 (
      {stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[6],stage2_15[7],stage2_14[8],stage2_13[10]}
   );
   gpc117_4 gpc128 (
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage1_17[0]},
      {1'b0},
      {stage2_19[0],stage2_18[0],stage2_17[4],stage2_16[7]}
   );
   gpc117_4 gpc129 (
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12], stage1_16[13]},
      {stage1_17[1]},
      {1'b0},
      {stage2_19[1],stage2_18[1],stage2_17[5],stage2_16[8]}
   );
   gpc1163_5 gpc130 (
      {stage1_16[14], stage1_16[15], stage1_16[16]},
      {stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5], stage1_17[6], stage1_17[7]},
      {1'b0},
      {1'b0},
      {stage2_20[0],stage2_19[2],stage2_18[2],stage2_17[6],stage2_16[9]}
   );
   gpc1_1 gpc131 (
      {stage1_0[9]},
      {stage2_0[3]}
   );
   gpc1_1 gpc132 (
      {stage1_0[10]},
      {stage2_0[4]}
   );
   gpc1_1 gpc133 (
      {stage1_0[11]},
      {stage2_0[5]}
   );
   gpc1_1 gpc134 (
      {stage1_0[12]},
      {stage2_0[6]}
   );
   gpc1_1 gpc135 (
      {stage1_0[13]},
      {stage2_0[7]}
   );
   gpc1_1 gpc136 (
      {stage1_2[21]},
      {stage2_2[6]}
   );
   gpc1_1 gpc137 (
      {stage1_2[22]},
      {stage2_2[7]}
   );
   gpc1_1 gpc138 (
      {stage1_4[34]},
      {stage2_4[11]}
   );
   gpc1_1 gpc139 (
      {stage1_5[24]},
      {stage2_5[9]}
   );
   gpc1_1 gpc140 (
      {stage1_6[18]},
      {stage2_6[11]}
   );
   gpc1_1 gpc141 (
      {stage1_7[18]},
      {stage2_7[10]}
   );
   gpc1_1 gpc142 (
      {stage1_9[24]},
      {stage2_9[9]}
   );
   gpc1_1 gpc143 (
      {stage1_9[25]},
      {stage2_9[10]}
   );
   gpc1_1 gpc144 (
      {stage1_9[26]},
      {stage2_9[11]}
   );
   gpc1_1 gpc145 (
      {stage1_10[15]},
      {stage2_10[9]}
   );
   gpc1_1 gpc146 (
      {stage1_10[16]},
      {stage2_10[10]}
   );
   gpc1_1 gpc147 (
      {stage1_10[17]},
      {stage2_10[11]}
   );
   gpc1_1 gpc148 (
      {stage1_10[18]},
      {stage2_10[12]}
   );
   gpc207_4 gpc149 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5], stage2_0[6]},
      {stage2_2[0], stage2_2[1]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc150 (
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7]},
      {stage2_3[0]},
      {stage2_4[0]},
      {stage3_5[0],stage3_4[0],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc615_5 gpc151 (
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage2_4[1]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[2]}
   );
   gpc615_5 gpc152 (
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6]},
      {stage2_5[6]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[1],stage3_6[1],stage3_5[2],stage3_4[2]}
   );
   gpc615_5 gpc153 (
      {stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_5[7]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[2],stage3_6[2],stage3_5[3],stage3_4[3]}
   );
   gpc615_5 gpc154 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[3]}
   );
   gpc615_5 gpc155 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[1]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[4]}
   );
   gpc606_5 gpc156 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6], stage2_8[7]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[2],stage3_10[2],stage3_9[2],stage3_8[4]}
   );
   gpc7_3 gpc157 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11], stage2_10[12]},
      {stage3_12[1],stage3_11[3],stage3_10[3]}
   );
   gpc606_5 gpc158 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[4]}
   );
   gpc1343_5 gpc159 (
      {stage2_12[0], stage2_12[1], stage2_12[2]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9]},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[3]}
   );
   gpc615_5 gpc160 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7]},
      {stage2_13[10]},
      {stage2_14[3], stage2_14[4], stage2_14[5], stage2_14[6], stage2_14[7], stage2_14[8]},
      {stage3_16[1],stage3_15[2],stage3_14[2],stage3_13[2],stage3_12[4]}
   );
   gpc117_4 gpc161 (
      {stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6], stage2_15[7]},
      {stage2_16[0]},
      {stage2_17[0]},
      {stage3_18[0],stage3_17[0],stage3_16[2],stage3_15[3]}
   );
   gpc7_3 gpc162 (
      {stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6], stage2_16[7]},
      {stage3_18[1],stage3_17[1],stage3_16[3]}
   );
   gpc1325_5 gpc163 (
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage2_18[0], stage2_18[1]},
      {stage2_19[0], stage2_19[1], stage2_19[2]},
      {stage2_20[0]},
      {stage3_21[0],stage3_20[0],stage3_19[0],stage3_18[2],stage3_17[2]}
   );
   gpc1_1 gpc164 (
      {stage2_0[7]},
      {stage3_0[1]}
   );
   gpc1_1 gpc165 (
      {stage2_3[6]},
      {stage3_3[3]}
   );
   gpc1_1 gpc166 (
      {stage2_3[7]},
      {stage3_3[4]}
   );
   gpc1_1 gpc167 (
      {stage2_3[8]},
      {stage3_3[5]}
   );
   gpc1_1 gpc168 (
      {stage2_5[8]},
      {stage3_5[4]}
   );
   gpc1_1 gpc169 (
      {stage2_5[9]},
      {stage3_5[5]}
   );
   gpc1_1 gpc170 (
      {stage2_7[10]},
      {stage3_7[5]}
   );
   gpc1_1 gpc171 (
      {stage2_11[6]},
      {stage3_11[5]}
   );
   gpc1_1 gpc172 (
      {stage2_12[8]},
      {stage3_12[5]}
   );
   gpc1_1 gpc173 (
      {stage2_16[8]},
      {stage3_16[4]}
   );
   gpc1_1 gpc174 (
      {stage2_16[9]},
      {stage3_16[5]}
   );
   gpc1_1 gpc175 (
      {stage2_17[6]},
      {stage3_17[3]}
   );
   gpc1_1 gpc176 (
      {stage2_18[2]},
      {stage3_18[3]}
   );
   gpc2135_5 gpc177 (
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4]},
      {stage3_4[0], stage3_4[1], stage3_4[2]},
      {stage3_5[0]},
      {stage3_6[0], stage3_6[1]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0]}
   );
   gpc615_5 gpc178 (
      {stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_6[2]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[1]}
   );
   gpc135_4 gpc179 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1]}
   );
   gpc1163_5 gpc180 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc181 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], stage3_14[2]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc1163_5 gpc182 (
      {stage3_15[1], stage3_15[2], stage3_15[3]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage3_17[0]},
      {stage3_18[0]},
      {stage4_19[0],stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1]}
   );
   gpc1163_5 gpc183 (
      {stage3_17[1], stage3_17[2], stage3_17[3]},
      {stage3_18[1], stage3_18[2], stage3_18[3], 1'b0, 1'b0, 1'b0},
      {stage3_19[0]},
      {stage3_20[0]},
      {stage4_21[0],stage4_20[0],stage4_19[1],stage4_18[1],stage4_17[1]}
   );
   gpc1_1 gpc184 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc185 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc186 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc187 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc188 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc189 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc190 (
      {stage3_3[5]},
      {stage4_3[1]}
   );
   gpc1_1 gpc191 (
      {stage3_4[3]},
      {stage4_4[1]}
   );
   gpc1_1 gpc192 (
      {stage3_21[0]},
      {stage4_21[1]}
   );
endmodule
module rowadder2_1_22(input [21:0] src0, input [21:0] src1, output [22:0] dst0);
    wire [21:0] gene;
    wire [21:0] prop;
    wire [23:0] out;
    wire [23:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_20_gene (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(gene[20])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_20_prop (
        .I0(src0[20]),
        .I1(src1[20]),
        .O(prop[20])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_21_gene (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(gene[21])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_21_prop (
        .I0(src0[21]),
        .I1(src1[21]),
        .O(prop[21])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_23_20 (
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CI(carryout[19]),
        .CYINIT(1'h0),
        .DI({2'h0, gene[21:20]}),
        .S({2'h0, prop[21:20]})
    );
    assign dst0 = {carryout[21], out[21:0]};
endmodule


module comp2_1test_54_16();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    reg [15:0] src16;
    reg [15:0] src17;
    reg [15:0] src18;
    reg [15:0] src19;
    reg [15:0] src20;
    reg [15:0] src21;
    reg [15:0] src22;
    reg [15:0] src23;
    reg [15:0] src24;
    reg [15:0] src25;
    reg [15:0] src26;
    reg [15:0] src27;
    reg [15:0] src28;
    reg [15:0] src29;
    reg [15:0] src30;
    reg [15:0] src31;
    reg [15:0] src32;
    reg [15:0] src33;
    reg [15:0] src34;
    reg [15:0] src35;
    reg [15:0] src36;
    reg [15:0] src37;
    reg [15:0] src38;
    reg [15:0] src39;
    reg [15:0] src40;
    reg [15:0] src41;
    reg [15:0] src42;
    reg [15:0] src43;
    reg [15:0] src44;
    reg [15:0] src45;
    reg [15:0] src46;
    reg [15:0] src47;
    reg [15:0] src48;
    reg [15:0] src49;
    reg [15:0] src50;
    reg [15:0] src51;
    reg [15:0] src52;
    reg [15:0] src53;
    reg [21:0] exp;
    wire [21:0] dst;
    assign test = dst == exp;
    compressor2_1_54_16 compressor2_1_54_16_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .dst(dst)
    );
    initial begin
        $monitor("0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x %x", src0, src1, src2, src3, src4, src5, src6, src7, src8, src9, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, src32, src33, src34, src35, src36, src37, src38, src39, src40, src41, src42, src43, src44, src45, src46, src47, src48, src49, src50, src51, src52, src53, dst, exp, test);
        src0 <= 16'h47bb;
        src1 <= 16'h7638;
        src2 <= 16'h4936;
        src3 <= 16'h289;
        src4 <= 16'hc6e0;
        src5 <= 16'hccfa;
        src6 <= 16'h218c;
        src7 <= 16'h5bb9;
        src8 <= 16'hf2fd;
        src9 <= 16'h2f06;
        src10 <= 16'h23a3;
        src11 <= 16'h3f7a;
        src12 <= 16'h409c;
        src13 <= 16'h200b;
        src14 <= 16'haf67;
        src15 <= 16'h65c;
        src16 <= 16'hf564;
        src17 <= 16'h75ef;
        src18 <= 16'h4c50;
        src19 <= 16'h9b10;
        src20 <= 16'hd87;
        src21 <= 16'h8d23;
        src22 <= 16'h784;
        src23 <= 16'h6614;
        src24 <= 16'hd41e;
        src25 <= 16'hb167;
        src26 <= 16'h1aed;
        src27 <= 16'hd2dc;
        src28 <= 16'h2439;
        src29 <= 16'hf9a9;
        src30 <= 16'hfd24;
        src31 <= 16'hed45;
        src32 <= 16'h6f5f;
        src33 <= 16'h2146;
        src34 <= 16'h8663;
        src35 <= 16'hf31b;
        src36 <= 16'h7464;
        src37 <= 16'h8457;
        src38 <= 16'ha874;
        src39 <= 16'h516f;
        src40 <= 16'hd59c;
        src41 <= 16'hc21;
        src42 <= 16'hfcb3;
        src43 <= 16'h5813;
        src44 <= 16'h748e;
        src45 <= 16'h52df;
        src46 <= 16'hf442;
        src47 <= 16'h7b6d;
        src48 <= 16'h19e3;
        src49 <= 16'h29f2;
        src50 <= 16'h4fec;
        src51 <= 16'habe6;
        src52 <= 16'hf738;
        src53 <= 16'h8107;
        exp <= 22'h19af2f;
        #1
        src0 <= 16'h71fc;
        src1 <= 16'hcde7;
        src2 <= 16'hc3c3;
        src3 <= 16'h9216;
        src4 <= 16'h2a16;
        src5 <= 16'h60dc;
        src6 <= 16'h6405;
        src7 <= 16'hde6f;
        src8 <= 16'h87dc;
        src9 <= 16'h4305;
        src10 <= 16'h29fc;
        src11 <= 16'hd7b7;
        src12 <= 16'hfaea;
        src13 <= 16'hc01a;
        src14 <= 16'h1579;
        src15 <= 16'h3cbc;
        src16 <= 16'h34ab;
        src17 <= 16'h4535;
        src18 <= 16'hfb80;
        src19 <= 16'h2995;
        src20 <= 16'h1e66;
        src21 <= 16'he071;
        src22 <= 16'h53b5;
        src23 <= 16'h8545;
        src24 <= 16'hc9c9;
        src25 <= 16'hf7f4;
        src26 <= 16'h6071;
        src27 <= 16'h921;
        src28 <= 16'h7228;
        src29 <= 16'h2e7c;
        src30 <= 16'h3d78;
        src31 <= 16'he67b;
        src32 <= 16'hcd72;
        src33 <= 16'h29f4;
        src34 <= 16'h917b;
        src35 <= 16'hbb88;
        src36 <= 16'h6b78;
        src37 <= 16'h6bf4;
        src38 <= 16'hd563;
        src39 <= 16'h792b;
        src40 <= 16'ha08;
        src41 <= 16'h2fd;
        src42 <= 16'hdef4;
        src43 <= 16'h606f;
        src44 <= 16'hab7e;
        src45 <= 16'h20cb;
        src46 <= 16'he34c;
        src47 <= 16'h4d4e;
        src48 <= 16'h89af;
        src49 <= 16'h9b41;
        src50 <= 16'h5c;
        src51 <= 16'h2d1d;
        src52 <= 16'ha2d;
        src53 <= 16'h794e;
        exp <= 22'h192d2d;
        #1
        src0 <= 16'h78f8;
        src1 <= 16'hc569;
        src2 <= 16'hfb0d;
        src3 <= 16'h47a2;
        src4 <= 16'hb020;
        src5 <= 16'h7185;
        src6 <= 16'h99ac;
        src7 <= 16'hac54;
        src8 <= 16'hd899;
        src9 <= 16'h9118;
        src10 <= 16'hed7c;
        src11 <= 16'h1ea7;
        src12 <= 16'h2b31;
        src13 <= 16'hd92a;
        src14 <= 16'h9fed;
        src15 <= 16'h4280;
        src16 <= 16'h3de0;
        src17 <= 16'hec4;
        src18 <= 16'hd123;
        src19 <= 16'hffac;
        src20 <= 16'hc7ce;
        src21 <= 16'h222d;
        src22 <= 16'h59af;
        src23 <= 16'h2339;
        src24 <= 16'h36ba;
        src25 <= 16'hf503;
        src26 <= 16'hd64b;
        src27 <= 16'h6704;
        src28 <= 16'h48d5;
        src29 <= 16'hdf02;
        src30 <= 16'h1da1;
        src31 <= 16'hfbf8;
        src32 <= 16'h5c9a;
        src33 <= 16'h8127;
        src34 <= 16'h65af;
        src35 <= 16'h4856;
        src36 <= 16'hf632;
        src37 <= 16'h2e99;
        src38 <= 16'hdfc7;
        src39 <= 16'hea3d;
        src40 <= 16'h9b6b;
        src41 <= 16'h5594;
        src42 <= 16'h492f;
        src43 <= 16'h98b2;
        src44 <= 16'h6c5f;
        src45 <= 16'h606f;
        src46 <= 16'hff67;
        src47 <= 16'h4ff1;
        src48 <= 16'h3318;
        src49 <= 16'hca5f;
        src50 <= 16'hbc0b;
        src51 <= 16'h6762;
        src52 <= 16'he5e6;
        src53 <= 16'h989c;
        exp <= 22'h1d7d24;
        #1
        src0 <= 16'h98f1;
        src1 <= 16'hf727;
        src2 <= 16'h59f2;
        src3 <= 16'hdd0a;
        src4 <= 16'h21ce;
        src5 <= 16'h1068;
        src6 <= 16'h4241;
        src7 <= 16'h4ce7;
        src8 <= 16'he4f3;
        src9 <= 16'h1122;
        src10 <= 16'h32bb;
        src11 <= 16'hc834;
        src12 <= 16'h8ddb;
        src13 <= 16'he789;
        src14 <= 16'h42d4;
        src15 <= 16'h2729;
        src16 <= 16'h44ba;
        src17 <= 16'haf46;
        src18 <= 16'hab74;
        src19 <= 16'hcb71;
        src20 <= 16'h2de8;
        src21 <= 16'h6586;
        src22 <= 16'hd5bf;
        src23 <= 16'hb546;
        src24 <= 16'hdf1;
        src25 <= 16'h7521;
        src26 <= 16'hd842;
        src27 <= 16'h1a07;
        src28 <= 16'h767;
        src29 <= 16'heb70;
        src30 <= 16'h8dca;
        src31 <= 16'h8423;
        src32 <= 16'hfac9;
        src33 <= 16'hfa52;
        src34 <= 16'hbd9e;
        src35 <= 16'h3c86;
        src36 <= 16'hd557;
        src37 <= 16'h7ac5;
        src38 <= 16'h8b85;
        src39 <= 16'h4b9f;
        src40 <= 16'h2187;
        src41 <= 16'h6ff4;
        src42 <= 16'hd88;
        src43 <= 16'hf621;
        src44 <= 16'h2ed9;
        src45 <= 16'h3e82;
        src46 <= 16'hf04e;
        src47 <= 16'h1f92;
        src48 <= 16'h392a;
        src49 <= 16'h1d6e;
        src50 <= 16'h3e66;
        src51 <= 16'h3738;
        src52 <= 16'hedd2;
        src53 <= 16'h9f38;
        exp <= 22'h19de6c;
        #1
        src0 <= 16'h82f9;
        src1 <= 16'hda0b;
        src2 <= 16'he9bb;
        src3 <= 16'h1cd2;
        src4 <= 16'h122d;
        src5 <= 16'h607d;
        src6 <= 16'h6ade;
        src7 <= 16'hc002;
        src8 <= 16'h6b9f;
        src9 <= 16'hf57f;
        src10 <= 16'h17b2;
        src11 <= 16'h7427;
        src12 <= 16'h973e;
        src13 <= 16'he57d;
        src14 <= 16'h5b96;
        src15 <= 16'hcdf5;
        src16 <= 16'h1b4;
        src17 <= 16'h161a;
        src18 <= 16'h984;
        src19 <= 16'haff;
        src20 <= 16'ha753;
        src21 <= 16'hf033;
        src22 <= 16'ha233;
        src23 <= 16'h16fe;
        src24 <= 16'hb75f;
        src25 <= 16'hbbb0;
        src26 <= 16'hc384;
        src27 <= 16'h22d2;
        src28 <= 16'h9560;
        src29 <= 16'hb50c;
        src30 <= 16'h96f0;
        src31 <= 16'h3c36;
        src32 <= 16'h4ea9;
        src33 <= 16'h72e7;
        src34 <= 16'hbcb8;
        src35 <= 16'h2996;
        src36 <= 16'hb305;
        src37 <= 16'h9cd4;
        src38 <= 16'h3b5f;
        src39 <= 16'hcce7;
        src40 <= 16'h1386;
        src41 <= 16'hcd24;
        src42 <= 16'h32ba;
        src43 <= 16'ha9c8;
        src44 <= 16'h8308;
        src45 <= 16'h75ce;
        src46 <= 16'h44fc;
        src47 <= 16'h283;
        src48 <= 16'h8822;
        src49 <= 16'h11c0;
        src50 <= 16'h23f9;
        src51 <= 16'h2133;
        src52 <= 16'hee72;
        src53 <= 16'h3174;
        exp <= 22'h1884c9;
        #1
        src0 <= 16'hef4a;
        src1 <= 16'h2a70;
        src2 <= 16'hdf1d;
        src3 <= 16'hf5f6;
        src4 <= 16'h5c88;
        src5 <= 16'h910a;
        src6 <= 16'h535a;
        src7 <= 16'hc311;
        src8 <= 16'hf8a7;
        src9 <= 16'he7f1;
        src10 <= 16'h3f8e;
        src11 <= 16'h2d2a;
        src12 <= 16'h70fd;
        src13 <= 16'h5138;
        src14 <= 16'h982b;
        src15 <= 16'h6294;
        src16 <= 16'h805f;
        src17 <= 16'h2dab;
        src18 <= 16'he196;
        src19 <= 16'h3784;
        src20 <= 16'h6b54;
        src21 <= 16'h474d;
        src22 <= 16'h9478;
        src23 <= 16'h7aea;
        src24 <= 16'h4369;
        src25 <= 16'h58d7;
        src26 <= 16'h6275;
        src27 <= 16'he3d0;
        src28 <= 16'h6d5f;
        src29 <= 16'hc9e5;
        src30 <= 16'h52af;
        src31 <= 16'hd960;
        src32 <= 16'hd1ab;
        src33 <= 16'h738a;
        src34 <= 16'hebcb;
        src35 <= 16'he198;
        src36 <= 16'he201;
        src37 <= 16'hd76f;
        src38 <= 16'h9811;
        src39 <= 16'h1fca;
        src40 <= 16'h245c;
        src41 <= 16'h62cb;
        src42 <= 16'h4b54;
        src43 <= 16'h99e0;
        src44 <= 16'ha6e6;
        src45 <= 16'hcc7c;
        src46 <= 16'h7822;
        src47 <= 16'h8d55;
        src48 <= 16'h2c49;
        src49 <= 16'h75a5;
        src50 <= 16'hd077;
        src51 <= 16'h6e50;
        src52 <= 16'h8fe7;
        src53 <= 16'h16c4;
        exp <= 22'h1cbc84;
        #1
        src0 <= 16'h93c1;
        src1 <= 16'h93bb;
        src2 <= 16'hc684;
        src3 <= 16'hec90;
        src4 <= 16'h27e1;
        src5 <= 16'h7808;
        src6 <= 16'h4641;
        src7 <= 16'h8724;
        src8 <= 16'h547d;
        src9 <= 16'hf450;
        src10 <= 16'hb21f;
        src11 <= 16'hc010;
        src12 <= 16'ha595;
        src13 <= 16'h91e0;
        src14 <= 16'h6d49;
        src15 <= 16'h9680;
        src16 <= 16'h9952;
        src17 <= 16'h21ab;
        src18 <= 16'h8536;
        src19 <= 16'h28ca;
        src20 <= 16'h23c4;
        src21 <= 16'hfff7;
        src22 <= 16'hc7b1;
        src23 <= 16'h1311;
        src24 <= 16'h8b38;
        src25 <= 16'hc040;
        src26 <= 16'h7ccb;
        src27 <= 16'h4c96;
        src28 <= 16'h707;
        src29 <= 16'he72;
        src30 <= 16'h488b;
        src31 <= 16'h4271;
        src32 <= 16'h62c7;
        src33 <= 16'h7428;
        src34 <= 16'hf3d;
        src35 <= 16'hac1d;
        src36 <= 16'hd0ca;
        src37 <= 16'h2433;
        src38 <= 16'h5980;
        src39 <= 16'h9ae8;
        src40 <= 16'hc38d;
        src41 <= 16'h52cb;
        src42 <= 16'h4c5a;
        src43 <= 16'hb7cc;
        src44 <= 16'h1e18;
        src45 <= 16'h5203;
        src46 <= 16'h747;
        src47 <= 16'h6251;
        src48 <= 16'h6576;
        src49 <= 16'hb2be;
        src50 <= 16'h604f;
        src51 <= 16'h87c7;
        src52 <= 16'hfd55;
        src53 <= 16'h9b2b;
        exp <= 22'h196389;
        #1
        src0 <= 16'h9da2;
        src1 <= 16'hf99a;
        src2 <= 16'h6bb7;
        src3 <= 16'h923;
        src4 <= 16'ha70;
        src5 <= 16'hc34e;
        src6 <= 16'he7ed;
        src7 <= 16'hee82;
        src8 <= 16'hb033;
        src9 <= 16'hb5b;
        src10 <= 16'h67c;
        src11 <= 16'h2f57;
        src12 <= 16'h38c0;
        src13 <= 16'had6f;
        src14 <= 16'hd910;
        src15 <= 16'h50ad;
        src16 <= 16'h69df;
        src17 <= 16'h1738;
        src18 <= 16'h270f;
        src19 <= 16'h2331;
        src20 <= 16'hcd10;
        src21 <= 16'h43af;
        src22 <= 16'hd741;
        src23 <= 16'ha21c;
        src24 <= 16'hff6e;
        src25 <= 16'h344b;
        src26 <= 16'h2e09;
        src27 <= 16'h9aa3;
        src28 <= 16'hfcc2;
        src29 <= 16'h210f;
        src30 <= 16'hf4e5;
        src31 <= 16'hcc97;
        src32 <= 16'h4835;
        src33 <= 16'h8e54;
        src34 <= 16'hf79f;
        src35 <= 16'hf547;
        src36 <= 16'hfc52;
        src37 <= 16'h1a1f;
        src38 <= 16'hedb2;
        src39 <= 16'hb53a;
        src40 <= 16'ha06a;
        src41 <= 16'hdab5;
        src42 <= 16'h4ccd;
        src43 <= 16'hb9b7;
        src44 <= 16'hc857;
        src45 <= 16'hd3b;
        src46 <= 16'h1b3e;
        src47 <= 16'h8ca5;
        src48 <= 16'h4dd2;
        src49 <= 16'h3657;
        src50 <= 16'h6a3;
        src51 <= 16'h9012;
        src52 <= 16'h92e3;
        src53 <= 16'h7813;
        exp <= 22'h1b846d;
        #1
        src0 <= 16'h9edc;
        src1 <= 16'hd66;
        src2 <= 16'h52d;
        src3 <= 16'hbfa6;
        src4 <= 16'h895a;
        src5 <= 16'h287e;
        src6 <= 16'hd50a;
        src7 <= 16'h666;
        src8 <= 16'ha8fd;
        src9 <= 16'h1312;
        src10 <= 16'h7693;
        src11 <= 16'h6d78;
        src12 <= 16'ha9d0;
        src13 <= 16'h27cd;
        src14 <= 16'ha2ac;
        src15 <= 16'h112e;
        src16 <= 16'hfe05;
        src17 <= 16'hba38;
        src18 <= 16'h3050;
        src19 <= 16'h7728;
        src20 <= 16'hb416;
        src21 <= 16'he4d;
        src22 <= 16'h96c0;
        src23 <= 16'h67fd;
        src24 <= 16'hae42;
        src25 <= 16'hb9b1;
        src26 <= 16'h957f;
        src27 <= 16'hff60;
        src28 <= 16'he6f5;
        src29 <= 16'h1776;
        src30 <= 16'hde96;
        src31 <= 16'h294;
        src32 <= 16'h872e;
        src33 <= 16'h17d9;
        src34 <= 16'h93c3;
        src35 <= 16'hd6e7;
        src36 <= 16'h93a0;
        src37 <= 16'he9d4;
        src38 <= 16'h2d6d;
        src39 <= 16'h6281;
        src40 <= 16'h804a;
        src41 <= 16'h6c59;
        src42 <= 16'h7077;
        src43 <= 16'h81b9;
        src44 <= 16'h6850;
        src45 <= 16'he257;
        src46 <= 16'h9f3a;
        src47 <= 16'hbb5;
        src48 <= 16'h5412;
        src49 <= 16'h3e23;
        src50 <= 16'h576c;
        src51 <= 16'hebf6;
        src52 <= 16'h28a7;
        src53 <= 16'h17ee;
        exp <= 22'h1922d2;
        #1
        src0 <= 16'hbaca;
        src1 <= 16'hfbae;
        src2 <= 16'h5b41;
        src3 <= 16'h4b03;
        src4 <= 16'h7ec0;
        src5 <= 16'hdae4;
        src6 <= 16'hbc3b;
        src7 <= 16'h18db;
        src8 <= 16'hfc29;
        src9 <= 16'h5416;
        src10 <= 16'ha9d2;
        src11 <= 16'h46b4;
        src12 <= 16'h74e3;
        src13 <= 16'h2871;
        src14 <= 16'hafc3;
        src15 <= 16'h7a2b;
        src16 <= 16'ha518;
        src17 <= 16'hfc9a;
        src18 <= 16'h5629;
        src19 <= 16'h1c03;
        src20 <= 16'hf2c3;
        src21 <= 16'h8df3;
        src22 <= 16'h9dcf;
        src23 <= 16'hcd06;
        src24 <= 16'h3197;
        src25 <= 16'h3c6;
        src26 <= 16'heaf7;
        src27 <= 16'h4e6b;
        src28 <= 16'h2eff;
        src29 <= 16'hdc26;
        src30 <= 16'h5cb4;
        src31 <= 16'h6aa5;
        src32 <= 16'hf0e8;
        src33 <= 16'h5958;
        src34 <= 16'h9369;
        src35 <= 16'hd46b;
        src36 <= 16'hd888;
        src37 <= 16'h79be;
        src38 <= 16'hea37;
        src39 <= 16'h4d5b;
        src40 <= 16'h68f3;
        src41 <= 16'h4dbc;
        src42 <= 16'hef90;
        src43 <= 16'h2067;
        src44 <= 16'hefe0;
        src45 <= 16'h3e6d;
        src46 <= 16'hf104;
        src47 <= 16'h48ef;
        src48 <= 16'h1ce0;
        src49 <= 16'h5105;
        src50 <= 16'hb810;
        src51 <= 16'h7e10;
        src52 <= 16'hfd72;
        src53 <= 16'he7c1;
        exp <= 22'h1dc82d;
        #1
        src0 <= 16'h9869;
        src1 <= 16'hdae4;
        src2 <= 16'h4749;
        src3 <= 16'hd7a3;
        src4 <= 16'h4295;
        src5 <= 16'ha5f3;
        src6 <= 16'h9424;
        src7 <= 16'hd535;
        src8 <= 16'hb200;
        src9 <= 16'h2b21;
        src10 <= 16'hc12d;
        src11 <= 16'hd227;
        src12 <= 16'h87ec;
        src13 <= 16'h7395;
        src14 <= 16'ha276;
        src15 <= 16'h2285;
        src16 <= 16'h62f1;
        src17 <= 16'h2d7e;
        src18 <= 16'h7f99;
        src19 <= 16'h7b87;
        src20 <= 16'hc2a9;
        src21 <= 16'hfd0;
        src22 <= 16'h5641;
        src23 <= 16'h5a6d;
        src24 <= 16'he8e3;
        src25 <= 16'hc2b;
        src26 <= 16'hb10a;
        src27 <= 16'he5b0;
        src28 <= 16'h1930;
        src29 <= 16'h4de4;
        src30 <= 16'h7a20;
        src31 <= 16'h4346;
        src32 <= 16'h8334;
        src33 <= 16'hae20;
        src34 <= 16'ha3b3;
        src35 <= 16'h68c9;
        src36 <= 16'hcc7;
        src37 <= 16'ha07d;
        src38 <= 16'h6c90;
        src39 <= 16'h1b1c;
        src40 <= 16'hd5;
        src41 <= 16'h825a;
        src42 <= 16'hb04c;
        src43 <= 16'h5cf0;
        src44 <= 16'h55e4;
        src45 <= 16'h3172;
        src46 <= 16'h87c0;
        src47 <= 16'h9980;
        src48 <= 16'hb464;
        src49 <= 16'he8fb;
        src50 <= 16'h4b6a;
        src51 <= 16'he826;
        src52 <= 16'h3b85;
        src53 <= 16'h6415;
        exp <= 22'h19f04d;
        #1
        src0 <= 16'h3d67;
        src1 <= 16'h53b6;
        src2 <= 16'h1396;
        src3 <= 16'ha297;
        src4 <= 16'h221e;
        src5 <= 16'h7f41;
        src6 <= 16'hf95c;
        src7 <= 16'h4e5e;
        src8 <= 16'ha8be;
        src9 <= 16'hccfc;
        src10 <= 16'h6cff;
        src11 <= 16'hc851;
        src12 <= 16'h65f8;
        src13 <= 16'hbe61;
        src14 <= 16'h2f24;
        src15 <= 16'h8354;
        src16 <= 16'h37e6;
        src17 <= 16'h4674;
        src18 <= 16'hd67c;
        src19 <= 16'hb7a9;
        src20 <= 16'h5e07;
        src21 <= 16'h55b1;
        src22 <= 16'he8ec;
        src23 <= 16'h4f3c;
        src24 <= 16'hbef6;
        src25 <= 16'h7c7f;
        src26 <= 16'h7cf4;
        src27 <= 16'hd50d;
        src28 <= 16'hc50c;
        src29 <= 16'ha689;
        src30 <= 16'h828b;
        src31 <= 16'hf2e2;
        src32 <= 16'h80c1;
        src33 <= 16'h87fc;
        src34 <= 16'h256;
        src35 <= 16'h42da;
        src36 <= 16'hb3b2;
        src37 <= 16'h5d32;
        src38 <= 16'h6365;
        src39 <= 16'h5547;
        src40 <= 16'hdb77;
        src41 <= 16'h6ffa;
        src42 <= 16'h1728;
        src43 <= 16'he7a7;
        src44 <= 16'hf11a;
        src45 <= 16'hc2e5;
        src46 <= 16'hc60;
        src47 <= 16'h5356;
        src48 <= 16'h92c2;
        src49 <= 16'hbbe1;
        src50 <= 16'hf959;
        src51 <= 16'h782c;
        src52 <= 16'h74fe;
        src53 <= 16'h2fd7;
        exp <= 22'h1bf384;
        #1
        src0 <= 16'h5c8e;
        src1 <= 16'h8e46;
        src2 <= 16'h5171;
        src3 <= 16'h9212;
        src4 <= 16'hdbe9;
        src5 <= 16'h5352;
        src6 <= 16'h3d29;
        src7 <= 16'h8d67;
        src8 <= 16'h4e69;
        src9 <= 16'hfd9c;
        src10 <= 16'hd026;
        src11 <= 16'hf0a4;
        src12 <= 16'h1dde;
        src13 <= 16'h9de9;
        src14 <= 16'hfd3e;
        src15 <= 16'hfa9e;
        src16 <= 16'h2d6f;
        src17 <= 16'h3047;
        src18 <= 16'h30b6;
        src19 <= 16'hc053;
        src20 <= 16'hff9a;
        src21 <= 16'h33e0;
        src22 <= 16'h525f;
        src23 <= 16'hb8ba;
        src24 <= 16'hb974;
        src25 <= 16'h93c9;
        src26 <= 16'he83f;
        src27 <= 16'h47d3;
        src28 <= 16'h98e4;
        src29 <= 16'h5f74;
        src30 <= 16'h9397;
        src31 <= 16'h1e6;
        src32 <= 16'h46be;
        src33 <= 16'h62f7;
        src34 <= 16'h7fab;
        src35 <= 16'hc59;
        src36 <= 16'h1813;
        src37 <= 16'he947;
        src38 <= 16'h2301;
        src39 <= 16'h1c4;
        src40 <= 16'h65af;
        src41 <= 16'h2ec6;
        src42 <= 16'h5fe2;
        src43 <= 16'h267c;
        src44 <= 16'hff69;
        src45 <= 16'he1da;
        src46 <= 16'h8bad;
        src47 <= 16'ha7d8;
        src48 <= 16'ha4bd;
        src49 <= 16'he9ba;
        src50 <= 16'hcc4;
        src51 <= 16'h5a3;
        src52 <= 16'hc128;
        src53 <= 16'h7125;
        exp <= 22'h1a7fa8;
        #1
        src0 <= 16'h4b90;
        src1 <= 16'h2161;
        src2 <= 16'h6b56;
        src3 <= 16'h6404;
        src4 <= 16'h407;
        src5 <= 16'h7c04;
        src6 <= 16'h65c2;
        src7 <= 16'hd4b3;
        src8 <= 16'hbfe4;
        src9 <= 16'hea4d;
        src10 <= 16'h3d0;
        src11 <= 16'h23f;
        src12 <= 16'hca2e;
        src13 <= 16'h8589;
        src14 <= 16'hf211;
        src15 <= 16'h422c;
        src16 <= 16'h81ea;
        src17 <= 16'h587d;
        src18 <= 16'hb802;
        src19 <= 16'h306e;
        src20 <= 16'h97a2;
        src21 <= 16'h5142;
        src22 <= 16'h5b65;
        src23 <= 16'h6cb6;
        src24 <= 16'h7cd7;
        src25 <= 16'h8e34;
        src26 <= 16'h54d5;
        src27 <= 16'hdada;
        src28 <= 16'h97b3;
        src29 <= 16'h800a;
        src30 <= 16'hd114;
        src31 <= 16'hab57;
        src32 <= 16'h47b2;
        src33 <= 16'h87d9;
        src34 <= 16'hf178;
        src35 <= 16'h99af;
        src36 <= 16'hd897;
        src37 <= 16'h203a;
        src38 <= 16'he64e;
        src39 <= 16'h7993;
        src40 <= 16'h11c7;
        src41 <= 16'h5cec;
        src42 <= 16'h1176;
        src43 <= 16'h3583;
        src44 <= 16'hdd4c;
        src45 <= 16'h222;
        src46 <= 16'h5be1;
        src47 <= 16'hc134;
        src48 <= 16'h465f;
        src49 <= 16'h5812;
        src50 <= 16'h5f4c;
        src51 <= 16'h5edf;
        src52 <= 16'h6545;
        src53 <= 16'h3967;
        exp <= 22'h18ce92;
        #1
        src0 <= 16'h86d0;
        src1 <= 16'h69a4;
        src2 <= 16'h22d2;
        src3 <= 16'h2d31;
        src4 <= 16'h5080;
        src5 <= 16'hd779;
        src6 <= 16'hba80;
        src7 <= 16'h39a5;
        src8 <= 16'h1a14;
        src9 <= 16'h9d10;
        src10 <= 16'h8915;
        src11 <= 16'hf5e1;
        src12 <= 16'hb127;
        src13 <= 16'h88ef;
        src14 <= 16'h8fd7;
        src15 <= 16'h40f3;
        src16 <= 16'h8e3d;
        src17 <= 16'h51b4;
        src18 <= 16'h5c73;
        src19 <= 16'hd6f6;
        src20 <= 16'h918d;
        src21 <= 16'h5fa7;
        src22 <= 16'h6546;
        src23 <= 16'h8ac9;
        src24 <= 16'hd1ec;
        src25 <= 16'hf939;
        src26 <= 16'hf75;
        src27 <= 16'h1939;
        src28 <= 16'hd20e;
        src29 <= 16'ha48f;
        src30 <= 16'h392f;
        src31 <= 16'h3218;
        src32 <= 16'h70d4;
        src33 <= 16'hc6b0;
        src34 <= 16'h35c3;
        src35 <= 16'he6;
        src36 <= 16'h82f6;
        src37 <= 16'hd10b;
        src38 <= 16'hea36;
        src39 <= 16'ha9a9;
        src40 <= 16'h3a63;
        src41 <= 16'h6f68;
        src42 <= 16'h4ab8;
        src43 <= 16'h2ca4;
        src44 <= 16'h73da;
        src45 <= 16'h13ec;
        src46 <= 16'h1c94;
        src47 <= 16'he0bf;
        src48 <= 16'h4a69;
        src49 <= 16'h7de2;
        src50 <= 16'h8427;
        src51 <= 16'h46dd;
        src52 <= 16'h747c;
        src53 <= 16'hdd9c;
        exp <= 22'h194997;
        #1
        src0 <= 16'hca1c;
        src1 <= 16'h32d5;
        src2 <= 16'hca85;
        src3 <= 16'h7328;
        src4 <= 16'hb109;
        src5 <= 16'h7a81;
        src6 <= 16'hcdb6;
        src7 <= 16'h8739;
        src8 <= 16'hc29;
        src9 <= 16'hc07a;
        src10 <= 16'h6b37;
        src11 <= 16'h2dc3;
        src12 <= 16'h6db5;
        src13 <= 16'hd66b;
        src14 <= 16'h413d;
        src15 <= 16'h9812;
        src16 <= 16'h974f;
        src17 <= 16'he7ec;
        src18 <= 16'h4887;
        src19 <= 16'h6505;
        src20 <= 16'h9bcb;
        src21 <= 16'h6d4e;
        src22 <= 16'he118;
        src23 <= 16'h4666;
        src24 <= 16'h67d1;
        src25 <= 16'hb7e1;
        src26 <= 16'ha9c4;
        src27 <= 16'hfdba;
        src28 <= 16'h43cb;
        src29 <= 16'h8af2;
        src30 <= 16'hc944;
        src31 <= 16'hd28f;
        src32 <= 16'hfb66;
        src33 <= 16'h4211;
        src34 <= 16'hcb85;
        src35 <= 16'h5101;
        src36 <= 16'h6027;
        src37 <= 16'he8c2;
        src38 <= 16'hd027;
        src39 <= 16'h59e0;
        src40 <= 16'h18ec;
        src41 <= 16'h28ac;
        src42 <= 16'hf58a;
        src43 <= 16'h4a8f;
        src44 <= 16'hdffb;
        src45 <= 16'h6771;
        src46 <= 16'hcd13;
        src47 <= 16'hc1ef;
        src48 <= 16'h7f6a;
        src49 <= 16'h7f98;
        src50 <= 16'h2988;
        src51 <= 16'h111c;
        src52 <= 16'h7b8;
        src53 <= 16'h71d7;
        exp <= 22'h1ca582;
        #1
        src0 <= 16'h152b;
        src1 <= 16'h9e9e;
        src2 <= 16'hd6d6;
        src3 <= 16'hde1c;
        src4 <= 16'h9d2e;
        src5 <= 16'h1c9;
        src6 <= 16'hdae9;
        src7 <= 16'he69c;
        src8 <= 16'hf46;
        src9 <= 16'h62d3;
        src10 <= 16'hb9f6;
        src11 <= 16'h95a1;
        src12 <= 16'hd5c2;
        src13 <= 16'h6a99;
        src14 <= 16'h3a30;
        src15 <= 16'he531;
        src16 <= 16'ha15e;
        src17 <= 16'h4970;
        src18 <= 16'he9cf;
        src19 <= 16'h6fcd;
        src20 <= 16'h6e00;
        src21 <= 16'hfed9;
        src22 <= 16'h6713;
        src23 <= 16'hbdac;
        src24 <= 16'heb6e;
        src25 <= 16'hd83d;
        src26 <= 16'ha5af;
        src27 <= 16'hcd27;
        src28 <= 16'h2e3d;
        src29 <= 16'h46bf;
        src30 <= 16'h1782;
        src31 <= 16'h9b55;
        src32 <= 16'h5255;
        src33 <= 16'h4b8f;
        src34 <= 16'h169e;
        src35 <= 16'h5172;
        src36 <= 16'ha0e2;
        src37 <= 16'h9afd;
        src38 <= 16'h8b9a;
        src39 <= 16'h975b;
        src40 <= 16'h3bc6;
        src41 <= 16'h4394;
        src42 <= 16'h9910;
        src43 <= 16'hd81;
        src44 <= 16'h6cd6;
        src45 <= 16'h27e4;
        src46 <= 16'h9403;
        src47 <= 16'hcdc7;
        src48 <= 16'hbc31;
        src49 <= 16'hafdb;
        src50 <= 16'hedc6;
        src51 <= 16'h8df;
        src52 <= 16'he0d1;
        src53 <= 16'h96fc;
        exp <= 22'h1c7aae;
        #1
        src0 <= 16'h74da;
        src1 <= 16'hc88d;
        src2 <= 16'h7c38;
        src3 <= 16'h5f6e;
        src4 <= 16'h8e7b;
        src5 <= 16'hcb24;
        src6 <= 16'h2ad7;
        src7 <= 16'h3cb2;
        src8 <= 16'h27af;
        src9 <= 16'h677;
        src10 <= 16'hf8df;
        src11 <= 16'h2d3c;
        src12 <= 16'h265e;
        src13 <= 16'h4141;
        src14 <= 16'h5f42;
        src15 <= 16'h4a7c;
        src16 <= 16'hfcc1;
        src17 <= 16'h6f6d;
        src18 <= 16'h71cd;
        src19 <= 16'hfdd0;
        src20 <= 16'hbc20;
        src21 <= 16'h1b69;
        src22 <= 16'he5d4;
        src23 <= 16'h1c89;
        src24 <= 16'h870f;
        src25 <= 16'h7d8a;
        src26 <= 16'ha832;
        src27 <= 16'h2817;
        src28 <= 16'h707b;
        src29 <= 16'h773e;
        src30 <= 16'hae1e;
        src31 <= 16'h1d59;
        src32 <= 16'h43be;
        src33 <= 16'h902c;
        src34 <= 16'h82b6;
        src35 <= 16'ha5af;
        src36 <= 16'h77e0;
        src37 <= 16'h8c95;
        src38 <= 16'h24b2;
        src39 <= 16'haebd;
        src40 <= 16'h9132;
        src41 <= 16'hd246;
        src42 <= 16'h4fda;
        src43 <= 16'hf7cf;
        src44 <= 16'h5693;
        src45 <= 16'h7b87;
        src46 <= 16'h6ccf;
        src47 <= 16'hb7a8;
        src48 <= 16'h2388;
        src49 <= 16'hc9fc;
        src50 <= 16'he3dd;
        src51 <= 16'he7db;
        src52 <= 16'hdcb5;
        src53 <= 16'hd220;
        exp <= 22'h1b5b8c;
        #1
        src0 <= 16'h9977;
        src1 <= 16'hb6e3;
        src2 <= 16'h6358;
        src3 <= 16'hed5e;
        src4 <= 16'h2ed9;
        src5 <= 16'hc00b;
        src6 <= 16'h9d5f;
        src7 <= 16'h2f5b;
        src8 <= 16'h4d46;
        src9 <= 16'h48ed;
        src10 <= 16'hcfaa;
        src11 <= 16'h4c67;
        src12 <= 16'h7527;
        src13 <= 16'hfc43;
        src14 <= 16'hd5b7;
        src15 <= 16'hc36e;
        src16 <= 16'h2ffb;
        src17 <= 16'h1fe4;
        src18 <= 16'hfd4b;
        src19 <= 16'hc866;
        src20 <= 16'h7935;
        src21 <= 16'h72b1;
        src22 <= 16'h26eb;
        src23 <= 16'hdc86;
        src24 <= 16'hd851;
        src25 <= 16'h2c79;
        src26 <= 16'h9a77;
        src27 <= 16'hce8d;
        src28 <= 16'h4a10;
        src29 <= 16'h850f;
        src30 <= 16'h3233;
        src31 <= 16'ha927;
        src32 <= 16'he088;
        src33 <= 16'hf0c2;
        src34 <= 16'h9c80;
        src35 <= 16'h6c3a;
        src36 <= 16'h4b74;
        src37 <= 16'he840;
        src38 <= 16'h21fa;
        src39 <= 16'hf886;
        src40 <= 16'h6b8;
        src41 <= 16'hada5;
        src42 <= 16'hc837;
        src43 <= 16'hea11;
        src44 <= 16'hb35d;
        src45 <= 16'h72f9;
        src46 <= 16'h7f2a;
        src47 <= 16'he367;
        src48 <= 16'hd825;
        src49 <= 16'h9c5;
        src50 <= 16'h3a1f;
        src51 <= 16'hb4e8;
        src52 <= 16'haa4c;
        src53 <= 16'h2586;
        exp <= 22'h1def36;
        #1
        src0 <= 16'h597e;
        src1 <= 16'hbd09;
        src2 <= 16'h4b4d;
        src3 <= 16'h8e23;
        src4 <= 16'h2245;
        src5 <= 16'h9e1f;
        src6 <= 16'hf492;
        src7 <= 16'ha0c0;
        src8 <= 16'ha6ef;
        src9 <= 16'h8097;
        src10 <= 16'h693;
        src11 <= 16'hc2f0;
        src12 <= 16'h9955;
        src13 <= 16'hc746;
        src14 <= 16'h32e0;
        src15 <= 16'h244;
        src16 <= 16'h29b7;
        src17 <= 16'h5059;
        src18 <= 16'h10a5;
        src19 <= 16'h899;
        src20 <= 16'hb50b;
        src21 <= 16'hbd46;
        src22 <= 16'h1d44;
        src23 <= 16'h19f7;
        src24 <= 16'hc095;
        src25 <= 16'h769f;
        src26 <= 16'hc8c9;
        src27 <= 16'h5d78;
        src28 <= 16'h38ec;
        src29 <= 16'h216b;
        src30 <= 16'hd850;
        src31 <= 16'he61c;
        src32 <= 16'h4b58;
        src33 <= 16'ha045;
        src34 <= 16'heab7;
        src35 <= 16'hd359;
        src36 <= 16'hbaad;
        src37 <= 16'h6924;
        src38 <= 16'hb7c6;
        src39 <= 16'h357a;
        src40 <= 16'h5c2e;
        src41 <= 16'h3595;
        src42 <= 16'h7597;
        src43 <= 16'hdb63;
        src44 <= 16'h5c0;
        src45 <= 16'h1416;
        src46 <= 16'h29af;
        src47 <= 16'hedec;
        src48 <= 16'hddb8;
        src49 <= 16'h8df1;
        src50 <= 16'hdb01;
        src51 <= 16'h4030;
        src52 <= 16'h2000;
        src53 <= 16'h139f;
        exp <= 22'h1908ec;
        #1
        src0 <= 16'h47c2;
        src1 <= 16'h431c;
        src2 <= 16'h741b;
        src3 <= 16'h6f36;
        src4 <= 16'h7c7e;
        src5 <= 16'ha3c5;
        src6 <= 16'h2a0d;
        src7 <= 16'h9b4c;
        src8 <= 16'h8912;
        src9 <= 16'h4621;
        src10 <= 16'ha928;
        src11 <= 16'h6458;
        src12 <= 16'h261c;
        src13 <= 16'h4b44;
        src14 <= 16'hb246;
        src15 <= 16'hf7ef;
        src16 <= 16'h6e40;
        src17 <= 16'hf9ef;
        src18 <= 16'h5d77;
        src19 <= 16'h6814;
        src20 <= 16'hf8ca;
        src21 <= 16'h5543;
        src22 <= 16'h47bd;
        src23 <= 16'hadce;
        src24 <= 16'h6c6c;
        src25 <= 16'h4408;
        src26 <= 16'hfd92;
        src27 <= 16'h1542;
        src28 <= 16'he029;
        src29 <= 16'hcd03;
        src30 <= 16'h6444;
        src31 <= 16'hf240;
        src32 <= 16'h155f;
        src33 <= 16'h178;
        src34 <= 16'h58d6;
        src35 <= 16'h600a;
        src36 <= 16'hc78f;
        src37 <= 16'h22e6;
        src38 <= 16'h6163;
        src39 <= 16'h1744;
        src40 <= 16'h6bc4;
        src41 <= 16'hca77;
        src42 <= 16'h26a6;
        src43 <= 16'hd42b;
        src44 <= 16'hea38;
        src45 <= 16'h83b3;
        src46 <= 16'hb56f;
        src47 <= 16'had9;
        src48 <= 16'hb651;
        src49 <= 16'h73b8;
        src50 <= 16'h7243;
        src51 <= 16'h3be8;
        src52 <= 16'ha56;
        src53 <= 16'h6c76;
        exp <= 22'h19656f;
        #1
        src0 <= 16'h7ddc;
        src1 <= 16'h2473;
        src2 <= 16'h99a;
        src3 <= 16'h4095;
        src4 <= 16'h8bd9;
        src5 <= 16'h3875;
        src6 <= 16'hd1e2;
        src7 <= 16'h1a8e;
        src8 <= 16'h6dc8;
        src9 <= 16'ha5aa;
        src10 <= 16'hc368;
        src11 <= 16'h7f34;
        src12 <= 16'h8ca0;
        src13 <= 16'h17e3;
        src14 <= 16'ha981;
        src15 <= 16'h9df2;
        src16 <= 16'hf0a;
        src17 <= 16'ha8e3;
        src18 <= 16'h786c;
        src19 <= 16'h79c2;
        src20 <= 16'h7692;
        src21 <= 16'h8d89;
        src22 <= 16'hf8b9;
        src23 <= 16'hef14;
        src24 <= 16'h9da0;
        src25 <= 16'hd2dd;
        src26 <= 16'hf1fc;
        src27 <= 16'h5a97;
        src28 <= 16'heee0;
        src29 <= 16'h5440;
        src30 <= 16'hff6d;
        src31 <= 16'h8690;
        src32 <= 16'hc2b6;
        src33 <= 16'h1e74;
        src34 <= 16'hc2f;
        src35 <= 16'h5078;
        src36 <= 16'h6ad8;
        src37 <= 16'h9863;
        src38 <= 16'h7afa;
        src39 <= 16'h689d;
        src40 <= 16'h7f9e;
        src41 <= 16'hff87;
        src42 <= 16'h8e24;
        src43 <= 16'h4dec;
        src44 <= 16'h5668;
        src45 <= 16'h311b;
        src46 <= 16'h1bc6;
        src47 <= 16'h9194;
        src48 <= 16'h73e8;
        src49 <= 16'h31ae;
        src50 <= 16'h9a17;
        src51 <= 16'h718e;
        src52 <= 16'h5db9;
        src53 <= 16'hdebb;
        exp <= 22'h1a9dd4;
        #1
        src0 <= 16'he8ae;
        src1 <= 16'h4b2a;
        src2 <= 16'hd868;
        src3 <= 16'ha4cc;
        src4 <= 16'heb1e;
        src5 <= 16'ha847;
        src6 <= 16'hd3ae;
        src7 <= 16'h4fbc;
        src8 <= 16'h38ef;
        src9 <= 16'h75b5;
        src10 <= 16'h3042;
        src11 <= 16'haa9c;
        src12 <= 16'hbf67;
        src13 <= 16'h2db7;
        src14 <= 16'h6267;
        src15 <= 16'h5316;
        src16 <= 16'hfe01;
        src17 <= 16'h26e9;
        src18 <= 16'h4671;
        src19 <= 16'h3732;
        src20 <= 16'hac42;
        src21 <= 16'h4495;
        src22 <= 16'h7798;
        src23 <= 16'hcd1d;
        src24 <= 16'h434f;
        src25 <= 16'h3af4;
        src26 <= 16'h4628;
        src27 <= 16'ha09b;
        src28 <= 16'h9b9a;
        src29 <= 16'h4110;
        src30 <= 16'h81bf;
        src31 <= 16'h3020;
        src32 <= 16'h4917;
        src33 <= 16'h42c3;
        src34 <= 16'hc191;
        src35 <= 16'h87ef;
        src36 <= 16'ha326;
        src37 <= 16'hd082;
        src38 <= 16'h37ed;
        src39 <= 16'h5fab;
        src40 <= 16'hb40d;
        src41 <= 16'h32ab;
        src42 <= 16'h1e67;
        src43 <= 16'h6302;
        src44 <= 16'hfe0d;
        src45 <= 16'ha6e2;
        src46 <= 16'hebe6;
        src47 <= 16'h7ddd;
        src48 <= 16'h33b9;
        src49 <= 16'he5ec;
        src50 <= 16'h6f3e;
        src51 <= 16'h7047;
        src52 <= 16'h3a11;
        src53 <= 16'hdec7;
        exp <= 22'h1ac90f;
        #1
        src0 <= 16'h281b;
        src1 <= 16'hd93;
        src2 <= 16'h195c;
        src3 <= 16'h421d;
        src4 <= 16'h29bb;
        src5 <= 16'h755e;
        src6 <= 16'h69af;
        src7 <= 16'h4dc3;
        src8 <= 16'hdbe;
        src9 <= 16'h808a;
        src10 <= 16'h3d16;
        src11 <= 16'hd40a;
        src12 <= 16'hbc08;
        src13 <= 16'hf64d;
        src14 <= 16'hd663;
        src15 <= 16'he7e8;
        src16 <= 16'h2974;
        src17 <= 16'h301;
        src18 <= 16'h71d1;
        src19 <= 16'h5799;
        src20 <= 16'hec01;
        src21 <= 16'he533;
        src22 <= 16'h593a;
        src23 <= 16'hc900;
        src24 <= 16'h8135;
        src25 <= 16'hd41e;
        src26 <= 16'h12c2;
        src27 <= 16'hfb1e;
        src28 <= 16'h565d;
        src29 <= 16'h742e;
        src30 <= 16'hd61b;
        src31 <= 16'hd80a;
        src32 <= 16'h8169;
        src33 <= 16'h4f28;
        src34 <= 16'h79b2;
        src35 <= 16'hcb06;
        src36 <= 16'h8a05;
        src37 <= 16'h602c;
        src38 <= 16'h2232;
        src39 <= 16'h7cd9;
        src40 <= 16'h26e8;
        src41 <= 16'hb74f;
        src42 <= 16'hc2d8;
        src43 <= 16'heb0;
        src44 <= 16'hc6d4;
        src45 <= 16'h4dde;
        src46 <= 16'h5116;
        src47 <= 16'hd6fd;
        src48 <= 16'hea23;
        src49 <= 16'h8721;
        src50 <= 16'h88a1;
        src51 <= 16'hcb2e;
        src52 <= 16'hd2ef;
        src53 <= 16'h3c5d;
        exp <= 22'h1b1c52;
        #1
        src0 <= 16'h6ca1;
        src1 <= 16'h71ee;
        src2 <= 16'hc945;
        src3 <= 16'h715e;
        src4 <= 16'h8e51;
        src5 <= 16'h362f;
        src6 <= 16'ha5ae;
        src7 <= 16'h245e;
        src8 <= 16'h1f5c;
        src9 <= 16'hc0b6;
        src10 <= 16'h7c85;
        src11 <= 16'h63af;
        src12 <= 16'h1df8;
        src13 <= 16'h7546;
        src14 <= 16'h7001;
        src15 <= 16'h52fb;
        src16 <= 16'h9756;
        src17 <= 16'h3554;
        src18 <= 16'h40cc;
        src19 <= 16'ha66c;
        src20 <= 16'h34ce;
        src21 <= 16'hfe48;
        src22 <= 16'h6992;
        src23 <= 16'h2fb9;
        src24 <= 16'h4fc;
        src25 <= 16'h8e04;
        src26 <= 16'hbb58;
        src27 <= 16'hca6e;
        src28 <= 16'hf6f9;
        src29 <= 16'hcce0;
        src30 <= 16'h5f83;
        src31 <= 16'h1452;
        src32 <= 16'h3aef;
        src33 <= 16'hf536;
        src34 <= 16'h2dd1;
        src35 <= 16'hcd8c;
        src36 <= 16'h650f;
        src37 <= 16'h2cd9;
        src38 <= 16'hbaab;
        src39 <= 16'h9feb;
        src40 <= 16'heedf;
        src41 <= 16'h82e8;
        src42 <= 16'h46e2;
        src43 <= 16'h4c45;
        src44 <= 16'hf24a;
        src45 <= 16'hbde6;
        src46 <= 16'h1f3c;
        src47 <= 16'hb90d;
        src48 <= 16'he7f0;
        src49 <= 16'h475f;
        src50 <= 16'h7d6f;
        src51 <= 16'he06f;
        src52 <= 16'h818a;
        src53 <= 16'hb52c;
        exp <= 22'h1af83f;
        #1
        src0 <= 16'h7f85;
        src1 <= 16'hefdd;
        src2 <= 16'h747a;
        src3 <= 16'hc1c6;
        src4 <= 16'h2d57;
        src5 <= 16'h6c43;
        src6 <= 16'h57c9;
        src7 <= 16'he3d0;
        src8 <= 16'h2ad5;
        src9 <= 16'hdbbc;
        src10 <= 16'h509b;
        src11 <= 16'h603d;
        src12 <= 16'h9ea9;
        src13 <= 16'h7311;
        src14 <= 16'h88fd;
        src15 <= 16'h907d;
        src16 <= 16'h516c;
        src17 <= 16'hd1b5;
        src18 <= 16'hefcc;
        src19 <= 16'hb8dc;
        src20 <= 16'h71e4;
        src21 <= 16'h434c;
        src22 <= 16'hf30d;
        src23 <= 16'h2619;
        src24 <= 16'hec8d;
        src25 <= 16'h8d49;
        src26 <= 16'h1d37;
        src27 <= 16'h9462;
        src28 <= 16'hee09;
        src29 <= 16'h8dd1;
        src30 <= 16'h4477;
        src31 <= 16'hefed;
        src32 <= 16'h4dee;
        src33 <= 16'h19f;
        src34 <= 16'h6b26;
        src35 <= 16'hd0f0;
        src36 <= 16'hb016;
        src37 <= 16'he9c6;
        src38 <= 16'h35b2;
        src39 <= 16'h93c3;
        src40 <= 16'h9a38;
        src41 <= 16'h9292;
        src42 <= 16'h101;
        src43 <= 16'hfe4f;
        src44 <= 16'h486e;
        src45 <= 16'hc96;
        src46 <= 16'h734b;
        src47 <= 16'hd579;
        src48 <= 16'hcec4;
        src49 <= 16'h778c;
        src50 <= 16'h2814;
        src51 <= 16'h50c0;
        src52 <= 16'h54bc;
        src53 <= 16'h3566;
        exp <= 22'h1bd55a;
        #1
        src0 <= 16'hec73;
        src1 <= 16'h4f06;
        src2 <= 16'h1c96;
        src3 <= 16'hb0b9;
        src4 <= 16'h487;
        src5 <= 16'hce48;
        src6 <= 16'ha3cb;
        src7 <= 16'hc21b;
        src8 <= 16'h7495;
        src9 <= 16'h713c;
        src10 <= 16'hd8df;
        src11 <= 16'h233a;
        src12 <= 16'h4e7a;
        src13 <= 16'h50d7;
        src14 <= 16'h6752;
        src15 <= 16'h3632;
        src16 <= 16'h74b7;
        src17 <= 16'h5a1;
        src18 <= 16'hf12e;
        src19 <= 16'h4913;
        src20 <= 16'h68a3;
        src21 <= 16'he946;
        src22 <= 16'h223a;
        src23 <= 16'h190a;
        src24 <= 16'h53f4;
        src25 <= 16'h1641;
        src26 <= 16'h4bff;
        src27 <= 16'h82d0;
        src28 <= 16'hd1c5;
        src29 <= 16'hf739;
        src30 <= 16'h1373;
        src31 <= 16'h822f;
        src32 <= 16'heaaa;
        src33 <= 16'hc6a;
        src34 <= 16'h9f2f;
        src35 <= 16'hbf38;
        src36 <= 16'h5a97;
        src37 <= 16'h695f;
        src38 <= 16'h101a;
        src39 <= 16'h9e16;
        src40 <= 16'h8a97;
        src41 <= 16'h1d81;
        src42 <= 16'head3;
        src43 <= 16'h4f49;
        src44 <= 16'h4359;
        src45 <= 16'h136c;
        src46 <= 16'h3815;
        src47 <= 16'h2887;
        src48 <= 16'ha6d9;
        src49 <= 16'hb407;
        src50 <= 16'h40b9;
        src51 <= 16'hcbf2;
        src52 <= 16'h1979;
        src53 <= 16'h8c24;
        exp <= 22'h17a804;
        #1
        src0 <= 16'h3a41;
        src1 <= 16'h43d0;
        src2 <= 16'hf69c;
        src3 <= 16'hdb1c;
        src4 <= 16'h39c7;
        src5 <= 16'h23ef;
        src6 <= 16'h8f43;
        src7 <= 16'head2;
        src8 <= 16'he2c9;
        src9 <= 16'hfab5;
        src10 <= 16'hb610;
        src11 <= 16'h4008;
        src12 <= 16'hac13;
        src13 <= 16'hcd61;
        src14 <= 16'hcae0;
        src15 <= 16'hf9e9;
        src16 <= 16'h19ed;
        src17 <= 16'h70c2;
        src18 <= 16'heb4f;
        src19 <= 16'hcacb;
        src20 <= 16'h1702;
        src21 <= 16'h4290;
        src22 <= 16'h459c;
        src23 <= 16'h516c;
        src24 <= 16'h4080;
        src25 <= 16'h2ad7;
        src26 <= 16'h6ac4;
        src27 <= 16'h4c9c;
        src28 <= 16'h4234;
        src29 <= 16'he1f6;
        src30 <= 16'hbf9f;
        src31 <= 16'hc094;
        src32 <= 16'hee40;
        src33 <= 16'hfbc8;
        src34 <= 16'h8650;
        src35 <= 16'h39a3;
        src36 <= 16'h73ba;
        src37 <= 16'h8850;
        src38 <= 16'hb4b8;
        src39 <= 16'h6cfa;
        src40 <= 16'hb3a1;
        src41 <= 16'h7c87;
        src42 <= 16'hd1c;
        src43 <= 16'h27df;
        src44 <= 16'hbc41;
        src45 <= 16'h1d0b;
        src46 <= 16'h8de;
        src47 <= 16'hadc2;
        src48 <= 16'hdeb3;
        src49 <= 16'h9693;
        src50 <= 16'h3099;
        src51 <= 16'h5cf;
        src52 <= 16'he469;
        src53 <= 16'hd5df;
        exp <= 22'h1c549a;
        #1
        src0 <= 16'hbcf6;
        src1 <= 16'h2d27;
        src2 <= 16'he9d5;
        src3 <= 16'h6f06;
        src4 <= 16'had90;
        src5 <= 16'h42c9;
        src6 <= 16'hdc78;
        src7 <= 16'h4cf6;
        src8 <= 16'h6ca8;
        src9 <= 16'hcee5;
        src10 <= 16'h2e9f;
        src11 <= 16'h4db7;
        src12 <= 16'he81a;
        src13 <= 16'h9bb6;
        src14 <= 16'h173c;
        src15 <= 16'hbf5c;
        src16 <= 16'he57;
        src17 <= 16'haff1;
        src18 <= 16'h8db;
        src19 <= 16'h3bc5;
        src20 <= 16'hab22;
        src21 <= 16'h92c;
        src22 <= 16'hc80e;
        src23 <= 16'hbdc8;
        src24 <= 16'ha083;
        src25 <= 16'h5ebe;
        src26 <= 16'ha7e;
        src27 <= 16'h85e6;
        src28 <= 16'h3057;
        src29 <= 16'h2de2;
        src30 <= 16'h3544;
        src31 <= 16'h5a34;
        src32 <= 16'hdbe5;
        src33 <= 16'h789c;
        src34 <= 16'h61b8;
        src35 <= 16'h7935;
        src36 <= 16'h3dd5;
        src37 <= 16'ha752;
        src38 <= 16'h22f9;
        src39 <= 16'h943;
        src40 <= 16'h679f;
        src41 <= 16'hbb9a;
        src42 <= 16'h6f93;
        src43 <= 16'h6ee7;
        src44 <= 16'h33fe;
        src45 <= 16'hb568;
        src46 <= 16'h2ce8;
        src47 <= 16'h3286;
        src48 <= 16'h736;
        src49 <= 16'hf00b;
        src50 <= 16'hc444;
        src51 <= 16'hda9;
        src52 <= 16'h603f;
        src53 <= 16'hee;
        exp <= 22'h16df1f;
        #1
        src0 <= 16'h4a4a;
        src1 <= 16'h6a15;
        src2 <= 16'h7fca;
        src3 <= 16'h61be;
        src4 <= 16'hd4fb;
        src5 <= 16'h5f6;
        src6 <= 16'h4da8;
        src7 <= 16'ha42e;
        src8 <= 16'h7a38;
        src9 <= 16'h9a82;
        src10 <= 16'he690;
        src11 <= 16'hf6aa;
        src12 <= 16'he9c8;
        src13 <= 16'hfb57;
        src14 <= 16'h6068;
        src15 <= 16'h2557;
        src16 <= 16'hd22d;
        src17 <= 16'h1aaf;
        src18 <= 16'h57c0;
        src19 <= 16'h4990;
        src20 <= 16'h3f34;
        src21 <= 16'he893;
        src22 <= 16'ha612;
        src23 <= 16'hb279;
        src24 <= 16'hdbc3;
        src25 <= 16'h49e0;
        src26 <= 16'h820c;
        src27 <= 16'hf41e;
        src28 <= 16'hb48b;
        src29 <= 16'h780;
        src30 <= 16'h7049;
        src31 <= 16'h3d0b;
        src32 <= 16'h65a5;
        src33 <= 16'h9021;
        src34 <= 16'ha043;
        src35 <= 16'hc2e8;
        src36 <= 16'h27af;
        src37 <= 16'h8ff;
        src38 <= 16'hc135;
        src39 <= 16'hb8d9;
        src40 <= 16'h39b9;
        src41 <= 16'h2547;
        src42 <= 16'h1443;
        src43 <= 16'h313a;
        src44 <= 16'hfd4c;
        src45 <= 16'haabf;
        src46 <= 16'h936e;
        src47 <= 16'h356b;
        src48 <= 16'h2c3a;
        src49 <= 16'h8f27;
        src50 <= 16'h17c4;
        src51 <= 16'h646d;
        src52 <= 16'hf3f2;
        src53 <= 16'hd4c8;
        exp <= 22'h1aec84;
        #1
        src0 <= 16'h169b;
        src1 <= 16'ha608;
        src2 <= 16'h470b;
        src3 <= 16'h153f;
        src4 <= 16'h97d9;
        src5 <= 16'h1418;
        src6 <= 16'hb18a;
        src7 <= 16'hb925;
        src8 <= 16'hc177;
        src9 <= 16'hea5d;
        src10 <= 16'hfe60;
        src11 <= 16'h74ce;
        src12 <= 16'hcf02;
        src13 <= 16'he11c;
        src14 <= 16'h5e02;
        src15 <= 16'h696d;
        src16 <= 16'h50da;
        src17 <= 16'hfb63;
        src18 <= 16'h8ce0;
        src19 <= 16'h6ef9;
        src20 <= 16'h30ad;
        src21 <= 16'h1e4f;
        src22 <= 16'hcf3b;
        src23 <= 16'heb98;
        src24 <= 16'h54e3;
        src25 <= 16'h529c;
        src26 <= 16'h4219;
        src27 <= 16'h69a3;
        src28 <= 16'hfb47;
        src29 <= 16'h8b37;
        src30 <= 16'h9901;
        src31 <= 16'h8482;
        src32 <= 16'h687a;
        src33 <= 16'h40d9;
        src34 <= 16'hef19;
        src35 <= 16'h944d;
        src36 <= 16'h7a00;
        src37 <= 16'h3316;
        src38 <= 16'hb783;
        src39 <= 16'h9f29;
        src40 <= 16'h94cf;
        src41 <= 16'h5755;
        src42 <= 16'hc86a;
        src43 <= 16'h3a8e;
        src44 <= 16'h3af;
        src45 <= 16'h33e;
        src46 <= 16'ha877;
        src47 <= 16'h509d;
        src48 <= 16'h599c;
        src49 <= 16'heed0;
        src50 <= 16'hc13e;
        src51 <= 16'h2b43;
        src52 <= 16'h1fa5;
        src53 <= 16'hf154;
        exp <= 22'h1b74bb;
        #1
        src0 <= 16'h4219;
        src1 <= 16'h9997;
        src2 <= 16'h1eae;
        src3 <= 16'h95ea;
        src4 <= 16'hd183;
        src5 <= 16'he077;
        src6 <= 16'hdf13;
        src7 <= 16'he026;
        src8 <= 16'h8752;
        src9 <= 16'hab47;
        src10 <= 16'h27da;
        src11 <= 16'h9ce8;
        src12 <= 16'hc26f;
        src13 <= 16'hdba0;
        src14 <= 16'h76f6;
        src15 <= 16'h685f;
        src16 <= 16'he205;
        src17 <= 16'h7315;
        src18 <= 16'h4259;
        src19 <= 16'h1c83;
        src20 <= 16'h7b31;
        src21 <= 16'h5149;
        src22 <= 16'he70c;
        src23 <= 16'ha920;
        src24 <= 16'h749a;
        src25 <= 16'haf18;
        src26 <= 16'hd99;
        src27 <= 16'h58b5;
        src28 <= 16'h5672;
        src29 <= 16'hdd1d;
        src30 <= 16'hff93;
        src31 <= 16'h9706;
        src32 <= 16'h3de9;
        src33 <= 16'h47eb;
        src34 <= 16'h90b5;
        src35 <= 16'h1ec7;
        src36 <= 16'h3f87;
        src37 <= 16'ha345;
        src38 <= 16'ha00b;
        src39 <= 16'h9d8d;
        src40 <= 16'h8c6c;
        src41 <= 16'h2097;
        src42 <= 16'h20d5;
        src43 <= 16'hb41f;
        src44 <= 16'he1f1;
        src45 <= 16'hc469;
        src46 <= 16'hbca7;
        src47 <= 16'hd1c;
        src48 <= 16'h454e;
        src49 <= 16'hc4b5;
        src50 <= 16'h1f41;
        src51 <= 16'hb4;
        src52 <= 16'hd6c2;
        src53 <= 16'hbc85;
        exp <= 22'h1be005;
        #1
        src0 <= 16'h59be;
        src1 <= 16'h77b1;
        src2 <= 16'h4ad3;
        src3 <= 16'h2290;
        src4 <= 16'h90da;
        src5 <= 16'h888;
        src6 <= 16'h8af4;
        src7 <= 16'hc79a;
        src8 <= 16'hf1de;
        src9 <= 16'h8ed3;
        src10 <= 16'h4ba1;
        src11 <= 16'hb5e6;
        src12 <= 16'h18de;
        src13 <= 16'h87d0;
        src14 <= 16'h92c4;
        src15 <= 16'h8442;
        src16 <= 16'hda51;
        src17 <= 16'h4810;
        src18 <= 16'hef53;
        src19 <= 16'h2330;
        src20 <= 16'h958a;
        src21 <= 16'hb746;
        src22 <= 16'h8912;
        src23 <= 16'h2bbe;
        src24 <= 16'hdfb6;
        src25 <= 16'h121e;
        src26 <= 16'h8d54;
        src27 <= 16'hc25c;
        src28 <= 16'h96ca;
        src29 <= 16'h8ca4;
        src30 <= 16'h6a8c;
        src31 <= 16'hca03;
        src32 <= 16'h821b;
        src33 <= 16'h176b;
        src34 <= 16'h58cf;
        src35 <= 16'h1b0f;
        src36 <= 16'hb0e5;
        src37 <= 16'h5a17;
        src38 <= 16'ha906;
        src39 <= 16'habc9;
        src40 <= 16'h7f66;
        src41 <= 16'h4446;
        src42 <= 16'h246;
        src43 <= 16'h407a;
        src44 <= 16'he9d3;
        src45 <= 16'hcbb6;
        src46 <= 16'h7d2e;
        src47 <= 16'hb0c3;
        src48 <= 16'h3511;
        src49 <= 16'h8fec;
        src50 <= 16'hc9db;
        src51 <= 16'h4d55;
        src52 <= 16'ha66e;
        src53 <= 16'hd732;
        exp <= 22'h1ae595;
        #1
        src0 <= 16'he107;
        src1 <= 16'hbb6e;
        src2 <= 16'h35aa;
        src3 <= 16'h285c;
        src4 <= 16'hd2a8;
        src5 <= 16'h9c06;
        src6 <= 16'h46ac;
        src7 <= 16'h9327;
        src8 <= 16'hf84;
        src9 <= 16'hf074;
        src10 <= 16'h40a2;
        src11 <= 16'h24e6;
        src12 <= 16'h180d;
        src13 <= 16'hb26a;
        src14 <= 16'h9556;
        src15 <= 16'h8fe5;
        src16 <= 16'hd34a;
        src17 <= 16'hdb4e;
        src18 <= 16'hb78b;
        src19 <= 16'hf507;
        src20 <= 16'ha1ed;
        src21 <= 16'h229b;
        src22 <= 16'h54b7;
        src23 <= 16'h7195;
        src24 <= 16'haaff;
        src25 <= 16'h46c4;
        src26 <= 16'h521c;
        src27 <= 16'hbf9e;
        src28 <= 16'h9460;
        src29 <= 16'h8abe;
        src30 <= 16'h66ff;
        src31 <= 16'ha28e;
        src32 <= 16'h173c;
        src33 <= 16'h615a;
        src34 <= 16'hc3f9;
        src35 <= 16'hd1bd;
        src36 <= 16'hf731;
        src37 <= 16'h6b9e;
        src38 <= 16'h743;
        src39 <= 16'h686d;
        src40 <= 16'h99e9;
        src41 <= 16'h96e6;
        src42 <= 16'he0f1;
        src43 <= 16'h20bd;
        src44 <= 16'hd9f8;
        src45 <= 16'h3f8;
        src46 <= 16'hbca3;
        src47 <= 16'ha66e;
        src48 <= 16'h1a7a;
        src49 <= 16'hca2;
        src50 <= 16'hd253;
        src51 <= 16'h6fb4;
        src52 <= 16'h1858;
        src53 <= 16'h7d89;
        exp <= 22'h1afda1;
        #1
        src0 <= 16'hdd48;
        src1 <= 16'h6220;
        src2 <= 16'h8a97;
        src3 <= 16'h961e;
        src4 <= 16'heb2d;
        src5 <= 16'h5dad;
        src6 <= 16'hbd3b;
        src7 <= 16'hc0bf;
        src8 <= 16'h96d3;
        src9 <= 16'h597f;
        src10 <= 16'hf144;
        src11 <= 16'hd888;
        src12 <= 16'h1a77;
        src13 <= 16'h5774;
        src14 <= 16'h4efb;
        src15 <= 16'h3497;
        src16 <= 16'h7d07;
        src17 <= 16'h79c2;
        src18 <= 16'hcc2f;
        src19 <= 16'hae8;
        src20 <= 16'hbbf8;
        src21 <= 16'h1b2b;
        src22 <= 16'h240a;
        src23 <= 16'hcfe0;
        src24 <= 16'h9ad4;
        src25 <= 16'h963c;
        src26 <= 16'h2a4b;
        src27 <= 16'h9919;
        src28 <= 16'hb500;
        src29 <= 16'hd3a6;
        src30 <= 16'hb1b5;
        src31 <= 16'hde23;
        src32 <= 16'h7ddb;
        src33 <= 16'h3658;
        src34 <= 16'h1ecd;
        src35 <= 16'h6557;
        src36 <= 16'hb13c;
        src37 <= 16'h135a;
        src38 <= 16'h615c;
        src39 <= 16'hf8dc;
        src40 <= 16'hd1fe;
        src41 <= 16'hc3c2;
        src42 <= 16'h2f2d;
        src43 <= 16'hec98;
        src44 <= 16'hcda;
        src45 <= 16'hb106;
        src46 <= 16'ha3af;
        src47 <= 16'h8d7;
        src48 <= 16'h6b9d;
        src49 <= 16'h1648;
        src50 <= 16'h2575;
        src51 <= 16'hbb43;
        src52 <= 16'he85c;
        src53 <= 16'h4e45;
        exp <= 22'h1b88b9;
        #1
        src0 <= 16'hf7ad;
        src1 <= 16'hdfe0;
        src2 <= 16'hb657;
        src3 <= 16'h2930;
        src4 <= 16'h834f;
        src5 <= 16'he736;
        src6 <= 16'hef79;
        src7 <= 16'h756d;
        src8 <= 16'hba52;
        src9 <= 16'h739d;
        src10 <= 16'h4f27;
        src11 <= 16'h2ccb;
        src12 <= 16'h47e4;
        src13 <= 16'hb5df;
        src14 <= 16'hcea6;
        src15 <= 16'hce9c;
        src16 <= 16'h1e2e;
        src17 <= 16'h4fda;
        src18 <= 16'h1635;
        src19 <= 16'hf92f;
        src20 <= 16'h9a67;
        src21 <= 16'h4346;
        src22 <= 16'h4be8;
        src23 <= 16'h449;
        src24 <= 16'hbb5c;
        src25 <= 16'hfc08;
        src26 <= 16'h2737;
        src27 <= 16'hf2e4;
        src28 <= 16'h5f93;
        src29 <= 16'h70c4;
        src30 <= 16'hf520;
        src31 <= 16'h1968;
        src32 <= 16'h15d6;
        src33 <= 16'h6319;
        src34 <= 16'h3316;
        src35 <= 16'h5e8f;
        src36 <= 16'hd841;
        src37 <= 16'h1d47;
        src38 <= 16'h4504;
        src39 <= 16'h8bf7;
        src40 <= 16'h9ee4;
        src41 <= 16'h3495;
        src42 <= 16'hbf26;
        src43 <= 16'ha2ce;
        src44 <= 16'hee39;
        src45 <= 16'he0f7;
        src46 <= 16'h3a78;
        src47 <= 16'ha1ef;
        src48 <= 16'h16dd;
        src49 <= 16'hc88b;
        src50 <= 16'h29b9;
        src51 <= 16'hc918;
        src52 <= 16'h8b00;
        src53 <= 16'h3e81;
        exp <= 22'h1b74e2;
        #1
        src0 <= 16'h9aa4;
        src1 <= 16'h993b;
        src2 <= 16'hae66;
        src3 <= 16'h8c5a;
        src4 <= 16'h7a40;
        src5 <= 16'h8e5e;
        src6 <= 16'h103b;
        src7 <= 16'hfb43;
        src8 <= 16'ha748;
        src9 <= 16'h5ae4;
        src10 <= 16'h2e18;
        src11 <= 16'h6b7b;
        src12 <= 16'h4d50;
        src13 <= 16'h9c26;
        src14 <= 16'h68cf;
        src15 <= 16'hedf7;
        src16 <= 16'h8a0e;
        src17 <= 16'hd0;
        src18 <= 16'hdde8;
        src19 <= 16'h4c9b;
        src20 <= 16'h8952;
        src21 <= 16'h45c8;
        src22 <= 16'h81a5;
        src23 <= 16'h671d;
        src24 <= 16'hf33d;
        src25 <= 16'h205a;
        src26 <= 16'hba46;
        src27 <= 16'hf5b;
        src28 <= 16'hd046;
        src29 <= 16'h583d;
        src30 <= 16'ha711;
        src31 <= 16'h7849;
        src32 <= 16'hb97d;
        src33 <= 16'h37fe;
        src34 <= 16'h9971;
        src35 <= 16'h8de6;
        src36 <= 16'hc036;
        src37 <= 16'h1839;
        src38 <= 16'h5bfd;
        src39 <= 16'h2a7b;
        src40 <= 16'h9050;
        src41 <= 16'h606a;
        src42 <= 16'h66b1;
        src43 <= 16'h98c1;
        src44 <= 16'hd75f;
        src45 <= 16'h6dd1;
        src46 <= 16'hcdf3;
        src47 <= 16'hd846;
        src48 <= 16'h5030;
        src49 <= 16'habfd;
        src50 <= 16'hdc46;
        src51 <= 16'hf3da;
        src52 <= 16'hbe5e;
        src53 <= 16'h6b0d;
        exp <= 22'h1c3a0e;
        #1
        src0 <= 16'h3f8d;
        src1 <= 16'hd117;
        src2 <= 16'h458d;
        src3 <= 16'h6bac;
        src4 <= 16'h5229;
        src5 <= 16'h4e3b;
        src6 <= 16'hca9f;
        src7 <= 16'h2d64;
        src8 <= 16'hff5c;
        src9 <= 16'h252c;
        src10 <= 16'hb7dc;
        src11 <= 16'h7019;
        src12 <= 16'hfe8f;
        src13 <= 16'h5e66;
        src14 <= 16'hd3ad;
        src15 <= 16'h8b62;
        src16 <= 16'h1270;
        src17 <= 16'h4c36;
        src18 <= 16'hef3e;
        src19 <= 16'h4703;
        src20 <= 16'he74;
        src21 <= 16'h3fb3;
        src22 <= 16'hf67d;
        src23 <= 16'heaf3;
        src24 <= 16'ha0b6;
        src25 <= 16'h4728;
        src26 <= 16'heb73;
        src27 <= 16'h3ce6;
        src28 <= 16'h3459;
        src29 <= 16'hd6b8;
        src30 <= 16'h9531;
        src31 <= 16'h2d2d;
        src32 <= 16'h2ff;
        src33 <= 16'h5f79;
        src34 <= 16'h1fdc;
        src35 <= 16'hc53a;
        src36 <= 16'h6af8;
        src37 <= 16'hd965;
        src38 <= 16'hd3f5;
        src39 <= 16'ha991;
        src40 <= 16'h3e86;
        src41 <= 16'h548b;
        src42 <= 16'hbebb;
        src43 <= 16'h1096;
        src44 <= 16'h3af0;
        src45 <= 16'h2c06;
        src46 <= 16'hcc30;
        src47 <= 16'h363a;
        src48 <= 16'h7d59;
        src49 <= 16'h1bb6;
        src50 <= 16'h24c4;
        src51 <= 16'hd8bd;
        src52 <= 16'h4e21;
        src53 <= 16'h154;
        exp <= 22'h18c021;
        #1
        src0 <= 16'h6b42;
        src1 <= 16'h4b0f;
        src2 <= 16'h9e62;
        src3 <= 16'hb6dd;
        src4 <= 16'h43d1;
        src5 <= 16'h520e;
        src6 <= 16'h8adc;
        src7 <= 16'h8eca;
        src8 <= 16'hd7c0;
        src9 <= 16'hd838;
        src10 <= 16'h9fa6;
        src11 <= 16'hd668;
        src12 <= 16'hde2c;
        src13 <= 16'hee52;
        src14 <= 16'h9a42;
        src15 <= 16'hb913;
        src16 <= 16'hb87c;
        src17 <= 16'hf4dc;
        src18 <= 16'he4e2;
        src19 <= 16'h972e;
        src20 <= 16'h6f8;
        src21 <= 16'h14f9;
        src22 <= 16'he0f;
        src23 <= 16'hcc9a;
        src24 <= 16'h49c2;
        src25 <= 16'h3316;
        src26 <= 16'hde1f;
        src27 <= 16'ha94b;
        src28 <= 16'h3e37;
        src29 <= 16'h897b;
        src30 <= 16'h84ad;
        src31 <= 16'h74c7;
        src32 <= 16'h1e8f;
        src33 <= 16'h8fc9;
        src34 <= 16'h6ad4;
        src35 <= 16'hf883;
        src36 <= 16'hba93;
        src37 <= 16'h65fd;
        src38 <= 16'h9602;
        src39 <= 16'h3d11;
        src40 <= 16'h2981;
        src41 <= 16'hbaed;
        src42 <= 16'h129b;
        src43 <= 16'h2f8b;
        src44 <= 16'h78e0;
        src45 <= 16'h6894;
        src46 <= 16'ha5f7;
        src47 <= 16'h53a6;
        src48 <= 16'h4912;
        src49 <= 16'hb79a;
        src50 <= 16'h5a0;
        src51 <= 16'h6a2;
        src52 <= 16'h3b1d;
        src53 <= 16'ha81e;
        exp <= 22'h1add78;
        #1
        src0 <= 16'h3736;
        src1 <= 16'ha487;
        src2 <= 16'h1fd2;
        src3 <= 16'h978c;
        src4 <= 16'ha517;
        src5 <= 16'h981d;
        src6 <= 16'hd64f;
        src7 <= 16'he576;
        src8 <= 16'hbb01;
        src9 <= 16'hb79a;
        src10 <= 16'h762a;
        src11 <= 16'h9393;
        src12 <= 16'h7ddd;
        src13 <= 16'hbdf0;
        src14 <= 16'hc476;
        src15 <= 16'hde52;
        src16 <= 16'h4afd;
        src17 <= 16'h4000;
        src18 <= 16'ha4de;
        src19 <= 16'hbca7;
        src20 <= 16'h771a;
        src21 <= 16'h41c0;
        src22 <= 16'h8cc0;
        src23 <= 16'h420a;
        src24 <= 16'hfdce;
        src25 <= 16'h32be;
        src26 <= 16'hc668;
        src27 <= 16'h498b;
        src28 <= 16'h18e3;
        src29 <= 16'h95b;
        src30 <= 16'hc96;
        src31 <= 16'h9f75;
        src32 <= 16'h8ee7;
        src33 <= 16'h507a;
        src34 <= 16'h5a8f;
        src35 <= 16'hd08b;
        src36 <= 16'h3e73;
        src37 <= 16'h985e;
        src38 <= 16'h8e9e;
        src39 <= 16'h5a39;
        src40 <= 16'hd26c;
        src41 <= 16'haf14;
        src42 <= 16'hab93;
        src43 <= 16'h7ba9;
        src44 <= 16'h2e22;
        src45 <= 16'hc72a;
        src46 <= 16'h5932;
        src47 <= 16'h6be0;
        src48 <= 16'hcf3a;
        src49 <= 16'ha597;
        src50 <= 16'hcade;
        src51 <= 16'h8697;
        src52 <= 16'h4b36;
        src53 <= 16'hd05d;
        exp <= 22'h1c7905;
        #1
        src0 <= 16'hb910;
        src1 <= 16'h9d80;
        src2 <= 16'he21c;
        src3 <= 16'h12aa;
        src4 <= 16'h58d3;
        src5 <= 16'h3ac2;
        src6 <= 16'h57a7;
        src7 <= 16'h742f;
        src8 <= 16'hb21c;
        src9 <= 16'h5cea;
        src10 <= 16'hdf7e;
        src11 <= 16'h937c;
        src12 <= 16'h9717;
        src13 <= 16'h8184;
        src14 <= 16'hb01d;
        src15 <= 16'h84a3;
        src16 <= 16'h6caf;
        src17 <= 16'hdda5;
        src18 <= 16'hf067;
        src19 <= 16'h5d05;
        src20 <= 16'he855;
        src21 <= 16'hb25b;
        src22 <= 16'h4211;
        src23 <= 16'h8dd9;
        src24 <= 16'h3e27;
        src25 <= 16'hfe46;
        src26 <= 16'h6e56;
        src27 <= 16'h68fa;
        src28 <= 16'hcd87;
        src29 <= 16'h2c5b;
        src30 <= 16'h3f82;
        src31 <= 16'hb280;
        src32 <= 16'h66b;
        src33 <= 16'h5c75;
        src34 <= 16'he7c0;
        src35 <= 16'heb46;
        src36 <= 16'he638;
        src37 <= 16'h76be;
        src38 <= 16'haa9f;
        src39 <= 16'hcaf0;
        src40 <= 16'hdb70;
        src41 <= 16'h9c23;
        src42 <= 16'h3571;
        src43 <= 16'hb1d0;
        src44 <= 16'h1b10;
        src45 <= 16'h4165;
        src46 <= 16'h5eeb;
        src47 <= 16'h2ff6;
        src48 <= 16'he021;
        src49 <= 16'h7b7e;
        src50 <= 16'h2fa;
        src51 <= 16'h86c9;
        src52 <= 16'hda86;
        src53 <= 16'h1eee;
        exp <= 22'h1cad82;
        #1
        src0 <= 16'h7481;
        src1 <= 16'hef6f;
        src2 <= 16'ha89d;
        src3 <= 16'ha9ca;
        src4 <= 16'hfab0;
        src5 <= 16'hfaf;
        src6 <= 16'h76ad;
        src7 <= 16'h9e32;
        src8 <= 16'h1353;
        src9 <= 16'h87db;
        src10 <= 16'hbe80;
        src11 <= 16'h8e20;
        src12 <= 16'h87a1;
        src13 <= 16'h7506;
        src14 <= 16'h73ad;
        src15 <= 16'hcacd;
        src16 <= 16'h6d9;
        src17 <= 16'hd6a0;
        src18 <= 16'h5073;
        src19 <= 16'h170b;
        src20 <= 16'hfccd;
        src21 <= 16'h6986;
        src22 <= 16'hb412;
        src23 <= 16'h1e42;
        src24 <= 16'hc4f6;
        src25 <= 16'h2e61;
        src26 <= 16'hcc3a;
        src27 <= 16'hafe;
        src28 <= 16'h3137;
        src29 <= 16'hb9f9;
        src30 <= 16'h9cae;
        src31 <= 16'ha2cd;
        src32 <= 16'hb0a7;
        src33 <= 16'h5010;
        src34 <= 16'h5228;
        src35 <= 16'h3fcf;
        src36 <= 16'hf447;
        src37 <= 16'h6a5d;
        src38 <= 16'h3e76;
        src39 <= 16'ha6ff;
        src40 <= 16'h360c;
        src41 <= 16'h34cb;
        src42 <= 16'hd069;
        src43 <= 16'hc52a;
        src44 <= 16'h52ef;
        src45 <= 16'h81ea;
        src46 <= 16'h6953;
        src47 <= 16'h65d6;
        src48 <= 16'hd7bb;
        src49 <= 16'h8928;
        src50 <= 16'hd3a0;
        src51 <= 16'h1d18;
        src52 <= 16'h29db;
        src53 <= 16'h5dac;
        exp <= 22'h1abfb1;
        #1
        src0 <= 16'h1aaa;
        src1 <= 16'h86f5;
        src2 <= 16'h62a0;
        src3 <= 16'hd087;
        src4 <= 16'h682d;
        src5 <= 16'h6807;
        src6 <= 16'hb12d;
        src7 <= 16'hee62;
        src8 <= 16'hd37d;
        src9 <= 16'h1758;
        src10 <= 16'hc6ef;
        src11 <= 16'hc9d3;
        src12 <= 16'ha3dd;
        src13 <= 16'h8e42;
        src14 <= 16'hfbd8;
        src15 <= 16'h1e06;
        src16 <= 16'h6c50;
        src17 <= 16'h571b;
        src18 <= 16'h1c1b;
        src19 <= 16'h6913;
        src20 <= 16'hba36;
        src21 <= 16'h3ac8;
        src22 <= 16'h3c37;
        src23 <= 16'hd1ca;
        src24 <= 16'hde7f;
        src25 <= 16'ha609;
        src26 <= 16'haef5;
        src27 <= 16'hff1e;
        src28 <= 16'h79d4;
        src29 <= 16'h56bc;
        src30 <= 16'h5fe1;
        src31 <= 16'h3ccb;
        src32 <= 16'ha5cd;
        src33 <= 16'h396a;
        src34 <= 16'ha8a5;
        src35 <= 16'h5639;
        src36 <= 16'ha9d;
        src37 <= 16'h2882;
        src38 <= 16'h6973;
        src39 <= 16'h5edc;
        src40 <= 16'h57b9;
        src41 <= 16'he657;
        src42 <= 16'h288d;
        src43 <= 16'h7519;
        src44 <= 16'hefb5;
        src45 <= 16'h7596;
        src46 <= 16'ha1c1;
        src47 <= 16'ha573;
        src48 <= 16'h31c4;
        src49 <= 16'h3a9b;
        src50 <= 16'ha2db;
        src51 <= 16'h10ec;
        src52 <= 16'h5404;
        src53 <= 16'hf1f1;
        exp <= 22'h1abf5f;
        #1
        src0 <= 16'h6b10;
        src1 <= 16'hb7ff;
        src2 <= 16'h2251;
        src3 <= 16'h49bb;
        src4 <= 16'h5992;
        src5 <= 16'hae03;
        src6 <= 16'h75aa;
        src7 <= 16'h8427;
        src8 <= 16'h4154;
        src9 <= 16'h2f89;
        src10 <= 16'h40e5;
        src11 <= 16'h9e1d;
        src12 <= 16'h4d7;
        src13 <= 16'had3;
        src14 <= 16'h4107;
        src15 <= 16'he394;
        src16 <= 16'he047;
        src17 <= 16'h5d3a;
        src18 <= 16'h78cd;
        src19 <= 16'h9d78;
        src20 <= 16'hef41;
        src21 <= 16'hb212;
        src22 <= 16'h8efe;
        src23 <= 16'hb04c;
        src24 <= 16'hc825;
        src25 <= 16'he681;
        src26 <= 16'h9ade;
        src27 <= 16'h775c;
        src28 <= 16'h3b1c;
        src29 <= 16'h9c07;
        src30 <= 16'hbc6f;
        src31 <= 16'hc920;
        src32 <= 16'h9cc6;
        src33 <= 16'h72c6;
        src34 <= 16'haf1a;
        src35 <= 16'h5bdb;
        src36 <= 16'hbd4e;
        src37 <= 16'had64;
        src38 <= 16'he510;
        src39 <= 16'h8e3d;
        src40 <= 16'hab2e;
        src41 <= 16'he35b;
        src42 <= 16'he11a;
        src43 <= 16'h8b8c;
        src44 <= 16'h8315;
        src45 <= 16'h70a0;
        src46 <= 16'h8c26;
        src47 <= 16'ha434;
        src48 <= 16'hde22;
        src49 <= 16'h4dae;
        src50 <= 16'hcea2;
        src51 <= 16'hd90b;
        src52 <= 16'h5532;
        src53 <= 16'hda71;
        exp <= 22'h1e8178;
        #1
        src0 <= 16'hacd3;
        src1 <= 16'ha26b;
        src2 <= 16'ha743;
        src3 <= 16'he012;
        src4 <= 16'h4377;
        src5 <= 16'h7bf0;
        src6 <= 16'hef20;
        src7 <= 16'h4f8b;
        src8 <= 16'h4fee;
        src9 <= 16'he7f7;
        src10 <= 16'h7a94;
        src11 <= 16'hb2ed;
        src12 <= 16'h40cf;
        src13 <= 16'hff48;
        src14 <= 16'h2466;
        src15 <= 16'h8a41;
        src16 <= 16'hea89;
        src17 <= 16'h7a89;
        src18 <= 16'hc815;
        src19 <= 16'hc56d;
        src20 <= 16'had01;
        src21 <= 16'h3ad1;
        src22 <= 16'h1aa6;
        src23 <= 16'hba3e;
        src24 <= 16'h2399;
        src25 <= 16'h4693;
        src26 <= 16'h513b;
        src27 <= 16'h2e85;
        src28 <= 16'hf4f3;
        src29 <= 16'h85e0;
        src30 <= 16'h7af5;
        src31 <= 16'ha2b3;
        src32 <= 16'hfb86;
        src33 <= 16'hd0d5;
        src34 <= 16'h6551;
        src35 <= 16'hac4f;
        src36 <= 16'hdcdb;
        src37 <= 16'hfc87;
        src38 <= 16'hdadf;
        src39 <= 16'hc2c4;
        src40 <= 16'h86de;
        src41 <= 16'hc04c;
        src42 <= 16'ha1d3;
        src43 <= 16'h4c87;
        src44 <= 16'hf483;
        src45 <= 16'h88e9;
        src46 <= 16'h3410;
        src47 <= 16'h2166;
        src48 <= 16'h40ac;
        src49 <= 16'he0ce;
        src50 <= 16'h9b23;
        src51 <= 16'hf8c;
        src52 <= 16'h9b85;
        src53 <= 16'hf037;
        exp <= 22'h1f0fc5;
        #1
        src0 <= 16'h2ba3;
        src1 <= 16'h383a;
        src2 <= 16'hadc3;
        src3 <= 16'haaad;
        src4 <= 16'h7bab;
        src5 <= 16'ha8cd;
        src6 <= 16'hef3;
        src7 <= 16'hb73;
        src8 <= 16'hf773;
        src9 <= 16'h2e27;
        src10 <= 16'h5c2d;
        src11 <= 16'h6775;
        src12 <= 16'h2182;
        src13 <= 16'hd909;
        src14 <= 16'h1363;
        src15 <= 16'he724;
        src16 <= 16'h528c;
        src17 <= 16'h5a1;
        src18 <= 16'hd479;
        src19 <= 16'haaef;
        src20 <= 16'h477d;
        src21 <= 16'h8530;
        src22 <= 16'hc281;
        src23 <= 16'hdb76;
        src24 <= 16'h3c1c;
        src25 <= 16'h2b82;
        src26 <= 16'h61cd;
        src27 <= 16'h735e;
        src28 <= 16'h4d53;
        src29 <= 16'h17f5;
        src30 <= 16'h82fe;
        src31 <= 16'h369a;
        src32 <= 16'ha513;
        src33 <= 16'hd27d;
        src34 <= 16'hf52f;
        src35 <= 16'he9af;
        src36 <= 16'h9e30;
        src37 <= 16'ha338;
        src38 <= 16'h33f8;
        src39 <= 16'hdfe7;
        src40 <= 16'h3961;
        src41 <= 16'h7a5;
        src42 <= 16'he6bd;
        src43 <= 16'hd62a;
        src44 <= 16'h8b16;
        src45 <= 16'hc714;
        src46 <= 16'hde04;
        src47 <= 16'h23dc;
        src48 <= 16'h1a85;
        src49 <= 16'hdbac;
        src50 <= 16'hb728;
        src51 <= 16'h170c;
        src52 <= 16'h342b;
        src53 <= 16'hdb7c;
        exp <= 22'h1a4913;
        #1
        src0 <= 16'h2159;
        src1 <= 16'h5320;
        src2 <= 16'hf683;
        src3 <= 16'h2495;
        src4 <= 16'h744c;
        src5 <= 16'he5e;
        src6 <= 16'h9ff8;
        src7 <= 16'h9e54;
        src8 <= 16'h8ee;
        src9 <= 16'h68d4;
        src10 <= 16'hd006;
        src11 <= 16'hf7c9;
        src12 <= 16'h3e5a;
        src13 <= 16'hce64;
        src14 <= 16'h545;
        src15 <= 16'hc0bd;
        src16 <= 16'h923c;
        src17 <= 16'hf853;
        src18 <= 16'h492b;
        src19 <= 16'h7975;
        src20 <= 16'h84a4;
        src21 <= 16'h4d23;
        src22 <= 16'hd54e;
        src23 <= 16'hd605;
        src24 <= 16'h74ab;
        src25 <= 16'h7ae8;
        src26 <= 16'hd603;
        src27 <= 16'he4;
        src28 <= 16'hafaf;
        src29 <= 16'h636c;
        src30 <= 16'h41a4;
        src31 <= 16'h9edf;
        src32 <= 16'hddf1;
        src33 <= 16'hf41c;
        src34 <= 16'hae2b;
        src35 <= 16'hb4f2;
        src36 <= 16'h82a7;
        src37 <= 16'h9182;
        src38 <= 16'h2185;
        src39 <= 16'hf12;
        src40 <= 16'hb623;
        src41 <= 16'h26fe;
        src42 <= 16'he071;
        src43 <= 16'h192b;
        src44 <= 16'habd;
        src45 <= 16'h4455;
        src46 <= 16'hd579;
        src47 <= 16'hce93;
        src48 <= 16'h4f46;
        src49 <= 16'hbacf;
        src50 <= 16'hde7;
        src51 <= 16'hc08e;
        src52 <= 16'h38a3;
        src53 <= 16'h781a;
        exp <= 22'h1aae45;
        #1
        src0 <= 16'h45fe;
        src1 <= 16'hd956;
        src2 <= 16'hf29f;
        src3 <= 16'h1c48;
        src4 <= 16'he96e;
        src5 <= 16'ha310;
        src6 <= 16'h4ebd;
        src7 <= 16'hc6be;
        src8 <= 16'h5710;
        src9 <= 16'hd5b8;
        src10 <= 16'he325;
        src11 <= 16'hfa50;
        src12 <= 16'h5263;
        src13 <= 16'h5870;
        src14 <= 16'haf4e;
        src15 <= 16'h266e;
        src16 <= 16'hde53;
        src17 <= 16'h3ca3;
        src18 <= 16'hbf53;
        src19 <= 16'hfb51;
        src20 <= 16'he3f8;
        src21 <= 16'h5d08;
        src22 <= 16'hcb51;
        src23 <= 16'h8dd2;
        src24 <= 16'hb528;
        src25 <= 16'he80a;
        src26 <= 16'h5bc3;
        src27 <= 16'h97d;
        src28 <= 16'h9a8;
        src29 <= 16'hbaad;
        src30 <= 16'h5022;
        src31 <= 16'h9a95;
        src32 <= 16'h8284;
        src33 <= 16'hf9b2;
        src34 <= 16'h7a89;
        src35 <= 16'h834e;
        src36 <= 16'h97b1;
        src37 <= 16'hb27d;
        src38 <= 16'h6f94;
        src39 <= 16'he1f8;
        src40 <= 16'habee;
        src41 <= 16'h1d31;
        src42 <= 16'hc10;
        src43 <= 16'hb17f;
        src44 <= 16'ha326;
        src45 <= 16'ha610;
        src46 <= 16'h1d99;
        src47 <= 16'hdf67;
        src48 <= 16'hd02;
        src49 <= 16'h4092;
        src50 <= 16'hf9ec;
        src51 <= 16'hef95;
        src52 <= 16'h79bd;
        src53 <= 16'h103a;
        exp <= 22'h1e1ff2;
        #1
        src0 <= 16'h9206;
        src1 <= 16'h74a0;
        src2 <= 16'h13bd;
        src3 <= 16'h4e60;
        src4 <= 16'h9949;
        src5 <= 16'h7ed0;
        src6 <= 16'h78d4;
        src7 <= 16'hb926;
        src8 <= 16'h80a6;
        src9 <= 16'hf7a2;
        src10 <= 16'hb8ec;
        src11 <= 16'hda5d;
        src12 <= 16'hbe4a;
        src13 <= 16'h8901;
        src14 <= 16'h2860;
        src15 <= 16'h6858;
        src16 <= 16'h4d5a;
        src17 <= 16'h7136;
        src18 <= 16'hb08a;
        src19 <= 16'hea3d;
        src20 <= 16'hf5b2;
        src21 <= 16'h4d1;
        src22 <= 16'h5f83;
        src23 <= 16'h6a0b;
        src24 <= 16'hc056;
        src25 <= 16'h27f9;
        src26 <= 16'h4026;
        src27 <= 16'h9fc9;
        src28 <= 16'h8039;
        src29 <= 16'h2a87;
        src30 <= 16'h1c3c;
        src31 <= 16'h8b96;
        src32 <= 16'hb908;
        src33 <= 16'h32c7;
        src34 <= 16'he0b1;
        src35 <= 16'hcebc;
        src36 <= 16'h46f1;
        src37 <= 16'h413f;
        src38 <= 16'hb8ff;
        src39 <= 16'h461e;
        src40 <= 16'h208c;
        src41 <= 16'h6d40;
        src42 <= 16'hbdc7;
        src43 <= 16'h2410;
        src44 <= 16'h7c83;
        src45 <= 16'h370c;
        src46 <= 16'h3c2b;
        src47 <= 16'hed15;
        src48 <= 16'hea3a;
        src49 <= 16'hb418;
        src50 <= 16'hd633;
        src51 <= 16'heff1;
        src52 <= 16'h49a7;
        src53 <= 16'h50ee;
        exp <= 22'h1b3ca8;
        #1
        src0 <= 16'hea26;
        src1 <= 16'h4b25;
        src2 <= 16'hc45a;
        src3 <= 16'h5f05;
        src4 <= 16'hcc88;
        src5 <= 16'he626;
        src6 <= 16'h5487;
        src7 <= 16'h5378;
        src8 <= 16'hd740;
        src9 <= 16'h19e5;
        src10 <= 16'h6480;
        src11 <= 16'h85c2;
        src12 <= 16'hcbbc;
        src13 <= 16'hc144;
        src14 <= 16'hc0d1;
        src15 <= 16'h3be8;
        src16 <= 16'h2f71;
        src17 <= 16'h2def;
        src18 <= 16'h5941;
        src19 <= 16'hbce0;
        src20 <= 16'h5e9b;
        src21 <= 16'h72d6;
        src22 <= 16'h9cfb;
        src23 <= 16'h541a;
        src24 <= 16'h4d38;
        src25 <= 16'h9f55;
        src26 <= 16'h9dda;
        src27 <= 16'he133;
        src28 <= 16'hdd43;
        src29 <= 16'h2851;
        src30 <= 16'hc988;
        src31 <= 16'hb6c8;
        src32 <= 16'hb129;
        src33 <= 16'ha82e;
        src34 <= 16'he6ed;
        src35 <= 16'hc34b;
        src36 <= 16'h9a98;
        src37 <= 16'hc561;
        src38 <= 16'hdf9c;
        src39 <= 16'h7411;
        src40 <= 16'h3523;
        src41 <= 16'hf8c7;
        src42 <= 16'h8d4b;
        src43 <= 16'h1858;
        src44 <= 16'h28de;
        src45 <= 16'h8894;
        src46 <= 16'hae46;
        src47 <= 16'h8a68;
        src48 <= 16'hc218;
        src49 <= 16'h7c4e;
        src50 <= 16'hd6c7;
        src51 <= 16'h417a;
        src52 <= 16'h566;
        src53 <= 16'he60e;
        exp <= 22'h1df6f9;
        #1
        src0 <= 16'h2f2b;
        src1 <= 16'h5220;
        src2 <= 16'h8b55;
        src3 <= 16'he63f;
        src4 <= 16'hedeb;
        src5 <= 16'h7c2f;
        src6 <= 16'h250f;
        src7 <= 16'h7b3c;
        src8 <= 16'h1e99;
        src9 <= 16'h4e73;
        src10 <= 16'h1482;
        src11 <= 16'h8e4d;
        src12 <= 16'hd96b;
        src13 <= 16'h604b;
        src14 <= 16'hba15;
        src15 <= 16'h4012;
        src16 <= 16'h448b;
        src17 <= 16'hce0c;
        src18 <= 16'h28ee;
        src19 <= 16'h8164;
        src20 <= 16'h5505;
        src21 <= 16'hf8d3;
        src22 <= 16'h8cac;
        src23 <= 16'hd99c;
        src24 <= 16'h9767;
        src25 <= 16'hd8ce;
        src26 <= 16'h3650;
        src27 <= 16'h4b05;
        src28 <= 16'h6ac5;
        src29 <= 16'hea5c;
        src30 <= 16'h8c5a;
        src31 <= 16'h578b;
        src32 <= 16'hfb8f;
        src33 <= 16'h2d38;
        src34 <= 16'h4153;
        src35 <= 16'ha554;
        src36 <= 16'hcd21;
        src37 <= 16'h9022;
        src38 <= 16'hb2aa;
        src39 <= 16'h5a1b;
        src40 <= 16'hbba2;
        src41 <= 16'h9611;
        src42 <= 16'h5154;
        src43 <= 16'hd18d;
        src44 <= 16'h2dbb;
        src45 <= 16'h88a1;
        src46 <= 16'h649c;
        src47 <= 16'h9cbe;
        src48 <= 16'hf087;
        src49 <= 16'hb608;
        src50 <= 16'hc33b;
        src51 <= 16'hf12a;
        src52 <= 16'hdd2b;
        src53 <= 16'h85f7;
        exp <= 22'h1d406b;
        #1
        src0 <= 16'hedd;
        src1 <= 16'hb25f;
        src2 <= 16'hc7fa;
        src3 <= 16'h8775;
        src4 <= 16'ha3f0;
        src5 <= 16'ha81;
        src6 <= 16'hda92;
        src7 <= 16'he7de;
        src8 <= 16'h7033;
        src9 <= 16'hb814;
        src10 <= 16'h5ee1;
        src11 <= 16'hc63e;
        src12 <= 16'hcfa1;
        src13 <= 16'hdc8c;
        src14 <= 16'hb856;
        src15 <= 16'h6f81;
        src16 <= 16'hf9e4;
        src17 <= 16'h9e95;
        src18 <= 16'ha451;
        src19 <= 16'hbb02;
        src20 <= 16'h9bc6;
        src21 <= 16'h27b3;
        src22 <= 16'h4c6e;
        src23 <= 16'hd0e0;
        src24 <= 16'h847d;
        src25 <= 16'h4b25;
        src26 <= 16'h1c45;
        src27 <= 16'h8622;
        src28 <= 16'h2de8;
        src29 <= 16'h2a42;
        src30 <= 16'h9017;
        src31 <= 16'he4e5;
        src32 <= 16'h7bcf;
        src33 <= 16'h58ee;
        src34 <= 16'h6aed;
        src35 <= 16'hdcaf;
        src36 <= 16'h9feb;
        src37 <= 16'hddb4;
        src38 <= 16'h2366;
        src39 <= 16'h3bc3;
        src40 <= 16'he0f0;
        src41 <= 16'h1fd8;
        src42 <= 16'h9e44;
        src43 <= 16'hb672;
        src44 <= 16'h590c;
        src45 <= 16'h10a7;
        src46 <= 16'h224d;
        src47 <= 16'hc9ec;
        src48 <= 16'h8f28;
        src49 <= 16'h4691;
        src50 <= 16'h77d6;
        src51 <= 16'ha70d;
        src52 <= 16'hecda;
        src53 <= 16'hd395;
        exp <= 22'h1d144e;
        #1
        src0 <= 16'h9cb7;
        src1 <= 16'h33ae;
        src2 <= 16'h991c;
        src3 <= 16'h9e37;
        src4 <= 16'hf294;
        src5 <= 16'h7767;
        src6 <= 16'h4e79;
        src7 <= 16'hdc95;
        src8 <= 16'h21d7;
        src9 <= 16'he774;
        src10 <= 16'h8797;
        src11 <= 16'h3ed2;
        src12 <= 16'hb57;
        src13 <= 16'h62df;
        src14 <= 16'h4827;
        src15 <= 16'h48a8;
        src16 <= 16'h9369;
        src17 <= 16'hb72b;
        src18 <= 16'h56a;
        src19 <= 16'he24a;
        src20 <= 16'h554a;
        src21 <= 16'hbfd2;
        src22 <= 16'hbb3f;
        src23 <= 16'he6c2;
        src24 <= 16'hcca9;
        src25 <= 16'h5b81;
        src26 <= 16'hdaea;
        src27 <= 16'hbf71;
        src28 <= 16'hd259;
        src29 <= 16'hf755;
        src30 <= 16'h50cc;
        src31 <= 16'hda99;
        src32 <= 16'hbe4a;
        src33 <= 16'he885;
        src34 <= 16'h4810;
        src35 <= 16'h930;
        src36 <= 16'h7339;
        src37 <= 16'h8e48;
        src38 <= 16'h8d82;
        src39 <= 16'h96ba;
        src40 <= 16'h7e1e;
        src41 <= 16'he26f;
        src42 <= 16'h6722;
        src43 <= 16'h2f7;
        src44 <= 16'h517d;
        src45 <= 16'hfb87;
        src46 <= 16'hf2ae;
        src47 <= 16'hc3e5;
        src48 <= 16'h7292;
        src49 <= 16'hbcbd;
        src50 <= 16'hbe6;
        src51 <= 16'hde24;
        src52 <= 16'ha84b;
        src53 <= 16'h7a06;
        exp <= 22'h1e342a;
        #1
        src0 <= 16'hf45f;
        src1 <= 16'h77ef;
        src2 <= 16'ha5ba;
        src3 <= 16'hc8af;
        src4 <= 16'h9d42;
        src5 <= 16'h9a;
        src6 <= 16'h66ef;
        src7 <= 16'h7797;
        src8 <= 16'h8374;
        src9 <= 16'hdb8e;
        src10 <= 16'hdec9;
        src11 <= 16'hd060;
        src12 <= 16'ha8dc;
        src13 <= 16'h9d2;
        src14 <= 16'h2bda;
        src15 <= 16'h430;
        src16 <= 16'he0a2;
        src17 <= 16'h5a69;
        src18 <= 16'h22c;
        src19 <= 16'h7837;
        src20 <= 16'h4e7;
        src21 <= 16'ha46b;
        src22 <= 16'h249f;
        src23 <= 16'hf250;
        src24 <= 16'h3964;
        src25 <= 16'hacb8;
        src26 <= 16'h790;
        src27 <= 16'h38dc;
        src28 <= 16'h1b88;
        src29 <= 16'hbde8;
        src30 <= 16'he654;
        src31 <= 16'h4955;
        src32 <= 16'hd5c;
        src33 <= 16'h74d4;
        src34 <= 16'h7ce3;
        src35 <= 16'h343b;
        src36 <= 16'h6abc;
        src37 <= 16'hb5c4;
        src38 <= 16'h6d75;
        src39 <= 16'h8713;
        src40 <= 16'h3b56;
        src41 <= 16'he16c;
        src42 <= 16'hbe3;
        src43 <= 16'h992;
        src44 <= 16'h3216;
        src45 <= 16'h1bc4;
        src46 <= 16'h2727;
        src47 <= 16'hc117;
        src48 <= 16'he5b5;
        src49 <= 16'h95cb;
        src50 <= 16'h7d08;
        src51 <= 16'h6558;
        src52 <= 16'h677e;
        src53 <= 16'hbd70;
        exp <= 22'h1820bf;
        #1
        src0 <= 16'hf916;
        src1 <= 16'hbf9;
        src2 <= 16'h9f94;
        src3 <= 16'h566e;
        src4 <= 16'he916;
        src5 <= 16'h82fd;
        src6 <= 16'h362e;
        src7 <= 16'h8e5a;
        src8 <= 16'hd965;
        src9 <= 16'h5379;
        src10 <= 16'h95b2;
        src11 <= 16'h191a;
        src12 <= 16'h6453;
        src13 <= 16'hd9ae;
        src14 <= 16'hf8b2;
        src15 <= 16'hd93c;
        src16 <= 16'h71c5;
        src17 <= 16'h675a;
        src18 <= 16'h1db9;
        src19 <= 16'h9ff4;
        src20 <= 16'hfc4a;
        src21 <= 16'h79b0;
        src22 <= 16'h611d;
        src23 <= 16'h6585;
        src24 <= 16'h2a49;
        src25 <= 16'h2b93;
        src26 <= 16'hc7e7;
        src27 <= 16'h60e9;
        src28 <= 16'hcff5;
        src29 <= 16'hf0d2;
        src30 <= 16'hb9db;
        src31 <= 16'hb3cb;
        src32 <= 16'hd62;
        src33 <= 16'h3f46;
        src34 <= 16'h5081;
        src35 <= 16'h105f;
        src36 <= 16'hc3dd;
        src37 <= 16'h1697;
        src38 <= 16'h5107;
        src39 <= 16'h229a;
        src40 <= 16'ha237;
        src41 <= 16'h5941;
        src42 <= 16'hc7ab;
        src43 <= 16'h3a50;
        src44 <= 16'h3f4d;
        src45 <= 16'h3db7;
        src46 <= 16'hcaab;
        src47 <= 16'h3be0;
        src48 <= 16'h3201;
        src49 <= 16'hc258;
        src50 <= 16'h9ae4;
        src51 <= 16'h8671;
        src52 <= 16'h198;
        src53 <= 16'hb111;
        exp <= 22'h19dcbc;
        #1
        src0 <= 16'h69ad;
        src1 <= 16'h18d;
        src2 <= 16'he10;
        src3 <= 16'h3a63;
        src4 <= 16'ha544;
        src5 <= 16'h5481;
        src6 <= 16'h6e59;
        src7 <= 16'h3765;
        src8 <= 16'h9408;
        src9 <= 16'h9f92;
        src10 <= 16'h7970;
        src11 <= 16'h2ee8;
        src12 <= 16'h2179;
        src13 <= 16'he2b4;
        src14 <= 16'hff85;
        src15 <= 16'he86e;
        src16 <= 16'ha89d;
        src17 <= 16'h2532;
        src18 <= 16'h8c4a;
        src19 <= 16'h8b11;
        src20 <= 16'h6b9;
        src21 <= 16'hf074;
        src22 <= 16'hc00;
        src23 <= 16'h8a3b;
        src24 <= 16'h56b6;
        src25 <= 16'h56ae;
        src26 <= 16'h72ab;
        src27 <= 16'h7723;
        src28 <= 16'hd93e;
        src29 <= 16'h20d6;
        src30 <= 16'h2e66;
        src31 <= 16'h5f39;
        src32 <= 16'h6594;
        src33 <= 16'h84ce;
        src34 <= 16'hd890;
        src35 <= 16'h4103;
        src36 <= 16'h2775;
        src37 <= 16'h9528;
        src38 <= 16'h460e;
        src39 <= 16'h1d83;
        src40 <= 16'ha0d7;
        src41 <= 16'hbe91;
        src42 <= 16'h32f5;
        src43 <= 16'h451b;
        src44 <= 16'h6990;
        src45 <= 16'h9284;
        src46 <= 16'hfd3a;
        src47 <= 16'hc0ef;
        src48 <= 16'hcd12;
        src49 <= 16'he810;
        src50 <= 16'h9ed6;
        src51 <= 16'h75a9;
        src52 <= 16'hc743;
        src53 <= 16'h38e4;
        exp <= 22'h192c59;
        #1
        src0 <= 16'h9fe6;
        src1 <= 16'hd802;
        src2 <= 16'h259;
        src3 <= 16'h6883;
        src4 <= 16'h2cf0;
        src5 <= 16'h2229;
        src6 <= 16'hb51e;
        src7 <= 16'he40d;
        src8 <= 16'hf0f3;
        src9 <= 16'hd2e0;
        src10 <= 16'h1f75;
        src11 <= 16'h7eca;
        src12 <= 16'heab;
        src13 <= 16'hb714;
        src14 <= 16'h3f71;
        src15 <= 16'hb288;
        src16 <= 16'h2719;
        src17 <= 16'hf937;
        src18 <= 16'h5d05;
        src19 <= 16'hedd0;
        src20 <= 16'hb1e;
        src21 <= 16'ha8ed;
        src22 <= 16'h9197;
        src23 <= 16'hebc5;
        src24 <= 16'h615f;
        src25 <= 16'h8c31;
        src26 <= 16'h5d71;
        src27 <= 16'h2260;
        src28 <= 16'ha76;
        src29 <= 16'h1787;
        src30 <= 16'h5c38;
        src31 <= 16'h2653;
        src32 <= 16'hd843;
        src33 <= 16'hb90f;
        src34 <= 16'hafe;
        src35 <= 16'hde01;
        src36 <= 16'h4857;
        src37 <= 16'h95c0;
        src38 <= 16'h1fda;
        src39 <= 16'h4216;
        src40 <= 16'h840e;
        src41 <= 16'hd79d;
        src42 <= 16'h1d61;
        src43 <= 16'h940b;
        src44 <= 16'h99bb;
        src45 <= 16'hd1cc;
        src46 <= 16'hb8cc;
        src47 <= 16'h888b;
        src48 <= 16'h5e61;
        src49 <= 16'hbb71;
        src50 <= 16'hc2e5;
        src51 <= 16'h8df0;
        src52 <= 16'hb14;
        src53 <= 16'h9d14;
        exp <= 22'h1a1a63;
        #1
        src0 <= 16'h8fef;
        src1 <= 16'h1808;
        src2 <= 16'h1349;
        src3 <= 16'h4d9d;
        src4 <= 16'h8375;
        src5 <= 16'h8282;
        src6 <= 16'hf8ba;
        src7 <= 16'hfc97;
        src8 <= 16'hd114;
        src9 <= 16'h61f9;
        src10 <= 16'h2708;
        src11 <= 16'hcb19;
        src12 <= 16'h307a;
        src13 <= 16'he2de;
        src14 <= 16'hbd72;
        src15 <= 16'h7c61;
        src16 <= 16'h5613;
        src17 <= 16'hb530;
        src18 <= 16'h1db7;
        src19 <= 16'h6063;
        src20 <= 16'he16c;
        src21 <= 16'hb2d6;
        src22 <= 16'h3145;
        src23 <= 16'hc50;
        src24 <= 16'h4e90;
        src25 <= 16'he8d6;
        src26 <= 16'hc3a7;
        src27 <= 16'h6779;
        src28 <= 16'h3305;
        src29 <= 16'hb2e6;
        src30 <= 16'h3b45;
        src31 <= 16'hb069;
        src32 <= 16'hf051;
        src33 <= 16'h5e0e;
        src34 <= 16'hb630;
        src35 <= 16'h6e6b;
        src36 <= 16'h22ba;
        src37 <= 16'h979d;
        src38 <= 16'h8fc;
        src39 <= 16'h4421;
        src40 <= 16'he2fe;
        src41 <= 16'h98e3;
        src42 <= 16'h681;
        src43 <= 16'h3180;
        src44 <= 16'h35e6;
        src45 <= 16'heb3;
        src46 <= 16'h4e5e;
        src47 <= 16'h12c0;
        src48 <= 16'haf23;
        src49 <= 16'h8e4f;
        src50 <= 16'h7e1b;
        src51 <= 16'h836d;
        src52 <= 16'h2915;
        src53 <= 16'h1743;
        exp <= 22'h18592a;
        #1
        src0 <= 16'h6e72;
        src1 <= 16'h59e7;
        src2 <= 16'hb691;
        src3 <= 16'hd1d0;
        src4 <= 16'hf7d6;
        src5 <= 16'hac1e;
        src6 <= 16'hd0f7;
        src7 <= 16'hfa5c;
        src8 <= 16'h5ae;
        src9 <= 16'h5f67;
        src10 <= 16'hb4ab;
        src11 <= 16'h7e1c;
        src12 <= 16'h8c35;
        src13 <= 16'h2bdf;
        src14 <= 16'hdf2a;
        src15 <= 16'hdc07;
        src16 <= 16'h9514;
        src17 <= 16'hb167;
        src18 <= 16'hd3be;
        src19 <= 16'hbc5c;
        src20 <= 16'h7c78;
        src21 <= 16'h23f3;
        src22 <= 16'hadfb;
        src23 <= 16'hdb5;
        src24 <= 16'hf250;
        src25 <= 16'hee68;
        src26 <= 16'hfb9d;
        src27 <= 16'h9f2b;
        src28 <= 16'hd50b;
        src29 <= 16'hcf96;
        src30 <= 16'h4149;
        src31 <= 16'ha7d5;
        src32 <= 16'hcf1c;
        src33 <= 16'hd61d;
        src34 <= 16'h23c;
        src35 <= 16'hfbf4;
        src36 <= 16'h96f4;
        src37 <= 16'h90a5;
        src38 <= 16'hfd0a;
        src39 <= 16'h3e2b;
        src40 <= 16'h95ec;
        src41 <= 16'h6620;
        src42 <= 16'hfbc2;
        src43 <= 16'h4feb;
        src44 <= 16'h5aa;
        src45 <= 16'h93d5;
        src46 <= 16'h8594;
        src47 <= 16'hfb5c;
        src48 <= 16'h7d36;
        src49 <= 16'hb579;
        src50 <= 16'had9f;
        src51 <= 16'hd908;
        src52 <= 16'hf267;
        src53 <= 16'h1577;
        exp <= 22'h2130a4;
        #1
        src0 <= 16'h3ca9;
        src1 <= 16'h3978;
        src2 <= 16'ha58d;
        src3 <= 16'hc789;
        src4 <= 16'h1e4c;
        src5 <= 16'hafbe;
        src6 <= 16'hac97;
        src7 <= 16'h7ba2;
        src8 <= 16'hc85;
        src9 <= 16'h4f1e;
        src10 <= 16'h127b;
        src11 <= 16'h57e0;
        src12 <= 16'he62a;
        src13 <= 16'h9a7c;
        src14 <= 16'h6211;
        src15 <= 16'h2ed1;
        src16 <= 16'h460f;
        src17 <= 16'ha89d;
        src18 <= 16'hbbe6;
        src19 <= 16'hf621;
        src20 <= 16'ha1d;
        src21 <= 16'h834;
        src22 <= 16'h2ba7;
        src23 <= 16'ha198;
        src24 <= 16'hdba9;
        src25 <= 16'h823b;
        src26 <= 16'hbdab;
        src27 <= 16'h3ba8;
        src28 <= 16'h3dcb;
        src29 <= 16'h933c;
        src30 <= 16'had27;
        src31 <= 16'h9f48;
        src32 <= 16'h4c7b;
        src33 <= 16'hff41;
        src34 <= 16'hde45;
        src35 <= 16'h96f9;
        src36 <= 16'h677;
        src37 <= 16'h579d;
        src38 <= 16'hdca7;
        src39 <= 16'hbcc7;
        src40 <= 16'ha6fb;
        src41 <= 16'h552a;
        src42 <= 16'h6404;
        src43 <= 16'hefc0;
        src44 <= 16'he999;
        src45 <= 16'h99a5;
        src46 <= 16'hf5b3;
        src47 <= 16'h4f96;
        src48 <= 16'hdc76;
        src49 <= 16'h126e;
        src50 <= 16'hc002;
        src51 <= 16'h5c47;
        src52 <= 16'h5dc0;
        src53 <= 16'h1704;
        exp <= 22'h1af6cd;
        #1
        src0 <= 16'h4449;
        src1 <= 16'h42cc;
        src2 <= 16'h49d3;
        src3 <= 16'h1d36;
        src4 <= 16'h7b5d;
        src5 <= 16'h1870;
        src6 <= 16'hf5a5;
        src7 <= 16'h58d7;
        src8 <= 16'h8d31;
        src9 <= 16'ha6c6;
        src10 <= 16'h34c6;
        src11 <= 16'h6539;
        src12 <= 16'h4451;
        src13 <= 16'he9e9;
        src14 <= 16'h61d5;
        src15 <= 16'hf666;
        src16 <= 16'hd5e6;
        src17 <= 16'h32b;
        src18 <= 16'hcb38;
        src19 <= 16'h15aa;
        src20 <= 16'hb6a7;
        src21 <= 16'h93fe;
        src22 <= 16'hfd49;
        src23 <= 16'h5e07;
        src24 <= 16'h2573;
        src25 <= 16'hfe9f;
        src26 <= 16'h7a3;
        src27 <= 16'hcca8;
        src28 <= 16'h72c9;
        src29 <= 16'hd5ce;
        src30 <= 16'hae17;
        src31 <= 16'he85b;
        src32 <= 16'h2b62;
        src33 <= 16'hd7a;
        src34 <= 16'hac6c;
        src35 <= 16'h8ef0;
        src36 <= 16'hcdcb;
        src37 <= 16'hceb7;
        src38 <= 16'hce5b;
        src39 <= 16'he6b8;
        src40 <= 16'h2ec9;
        src41 <= 16'hd4c3;
        src42 <= 16'h5d9e;
        src43 <= 16'hb6cc;
        src44 <= 16'h7a58;
        src45 <= 16'hfb66;
        src46 <= 16'h7e6e;
        src47 <= 16'h29fb;
        src48 <= 16'he0c7;
        src49 <= 16'hbdf;
        src50 <= 16'h4965;
        src51 <= 16'h1baa;
        src52 <= 16'hd79;
        src53 <= 16'h2bd9;
        exp <= 22'h1ae311;
        #1
        src0 <= 16'h3c39;
        src1 <= 16'h383f;
        src2 <= 16'hf4ae;
        src3 <= 16'h4f67;
        src4 <= 16'h890d;
        src5 <= 16'h7394;
        src6 <= 16'h4002;
        src7 <= 16'h6002;
        src8 <= 16'hf5d;
        src9 <= 16'ha117;
        src10 <= 16'h93aa;
        src11 <= 16'h62e1;
        src12 <= 16'h9f01;
        src13 <= 16'hb846;
        src14 <= 16'h54c;
        src15 <= 16'hc889;
        src16 <= 16'hdc17;
        src17 <= 16'hf1c4;
        src18 <= 16'h9f93;
        src19 <= 16'h885e;
        src20 <= 16'h6dae;
        src21 <= 16'hf0de;
        src22 <= 16'hbad9;
        src23 <= 16'hcc91;
        src24 <= 16'ha4c2;
        src25 <= 16'h6832;
        src26 <= 16'ha987;
        src27 <= 16'h5c92;
        src28 <= 16'h7948;
        src29 <= 16'h3693;
        src30 <= 16'h7017;
        src31 <= 16'h697;
        src32 <= 16'hcaba;
        src33 <= 16'h8541;
        src34 <= 16'h9072;
        src35 <= 16'h2b93;
        src36 <= 16'hfc99;
        src37 <= 16'h2f9c;
        src38 <= 16'he8e7;
        src39 <= 16'h2142;
        src40 <= 16'h23ee;
        src41 <= 16'hd715;
        src42 <= 16'h53ec;
        src43 <= 16'hf100;
        src44 <= 16'ha6b1;
        src45 <= 16'h2da4;
        src46 <= 16'h8ec0;
        src47 <= 16'h5031;
        src48 <= 16'h6d6e;
        src49 <= 16'hab97;
        src50 <= 16'h472e;
        src51 <= 16'h40b5;
        src52 <= 16'h7b92;
        src53 <= 16'h8c69;
        exp <= 22'h1b151b;
        #1
        src0 <= 16'hdd21;
        src1 <= 16'he3ab;
        src2 <= 16'h9c1;
        src3 <= 16'hc58a;
        src4 <= 16'hc6bb;
        src5 <= 16'h1f51;
        src6 <= 16'h76ac;
        src7 <= 16'h736f;
        src8 <= 16'h466c;
        src9 <= 16'h1a36;
        src10 <= 16'h4ae;
        src11 <= 16'h310c;
        src12 <= 16'h9b42;
        src13 <= 16'h816a;
        src14 <= 16'h4cc1;
        src15 <= 16'h68d;
        src16 <= 16'h9a0e;
        src17 <= 16'haff3;
        src18 <= 16'h39b9;
        src19 <= 16'he7e6;
        src20 <= 16'hba77;
        src21 <= 16'h53f3;
        src22 <= 16'h8ea4;
        src23 <= 16'h2279;
        src24 <= 16'h4547;
        src25 <= 16'h9a0d;
        src26 <= 16'he56d;
        src27 <= 16'ha3de;
        src28 <= 16'heb68;
        src29 <= 16'h6c5d;
        src30 <= 16'h1c43;
        src31 <= 16'h27fe;
        src32 <= 16'hc03d;
        src33 <= 16'hd63f;
        src34 <= 16'h90f0;
        src35 <= 16'hf2a6;
        src36 <= 16'h17d8;
        src37 <= 16'h6b8b;
        src38 <= 16'hae42;
        src39 <= 16'hd1db;
        src40 <= 16'he994;
        src41 <= 16'h877a;
        src42 <= 16'h94be;
        src43 <= 16'h86c4;
        src44 <= 16'h474c;
        src45 <= 16'hb5c0;
        src46 <= 16'h9e57;
        src47 <= 16'h10b9;
        src48 <= 16'h7db2;
        src49 <= 16'hdf3c;
        src50 <= 16'ha648;
        src51 <= 16'h69b1;
        src52 <= 16'h922f;
        src53 <= 16'h215a;
        exp <= 22'h1b0d0e;
        #1
        src0 <= 16'h87fa;
        src1 <= 16'h37d;
        src2 <= 16'hc07f;
        src3 <= 16'hd856;
        src4 <= 16'h13f8;
        src5 <= 16'hd82b;
        src6 <= 16'he61b;
        src7 <= 16'hc5e8;
        src8 <= 16'hb445;
        src9 <= 16'ha292;
        src10 <= 16'h69a3;
        src11 <= 16'hf07;
        src12 <= 16'hb0f8;
        src13 <= 16'h9a78;
        src14 <= 16'hd728;
        src15 <= 16'h385b;
        src16 <= 16'h3ef1;
        src17 <= 16'h1227;
        src18 <= 16'h2fd8;
        src19 <= 16'h5b06;
        src20 <= 16'ha13e;
        src21 <= 16'hd6e0;
        src22 <= 16'h18c;
        src23 <= 16'h8ee7;
        src24 <= 16'h8dcf;
        src25 <= 16'hcf24;
        src26 <= 16'h6867;
        src27 <= 16'h5ed2;
        src28 <= 16'h2b03;
        src29 <= 16'h96a6;
        src30 <= 16'h9db6;
        src31 <= 16'hfa39;
        src32 <= 16'h8984;
        src33 <= 16'h17;
        src34 <= 16'hfd34;
        src35 <= 16'ha126;
        src36 <= 16'h20ee;
        src37 <= 16'h2d43;
        src38 <= 16'h15d3;
        src39 <= 16'h2e17;
        src40 <= 16'hbbce;
        src41 <= 16'h1088;
        src42 <= 16'hbb08;
        src43 <= 16'hc9d8;
        src44 <= 16'h41d3;
        src45 <= 16'h9c3e;
        src46 <= 16'h7a69;
        src47 <= 16'hb907;
        src48 <= 16'ha9fd;
        src49 <= 16'hcbc;
        src50 <= 16'h4f41;
        src51 <= 16'hae04;
        src52 <= 16'hcfd6;
        src53 <= 16'he0a1;
        exp <= 22'h1aca6d;
        #1
        src0 <= 16'h5745;
        src1 <= 16'had12;
        src2 <= 16'hbab6;
        src3 <= 16'h7f16;
        src4 <= 16'haa49;
        src5 <= 16'h6064;
        src6 <= 16'h45b5;
        src7 <= 16'hf6cd;
        src8 <= 16'hece4;
        src9 <= 16'hb833;
        src10 <= 16'h2fd9;
        src11 <= 16'h85af;
        src12 <= 16'h8bc3;
        src13 <= 16'hd20a;
        src14 <= 16'heccf;
        src15 <= 16'h9dba;
        src16 <= 16'h38e9;
        src17 <= 16'h3318;
        src18 <= 16'hc9d5;
        src19 <= 16'hab9c;
        src20 <= 16'h7249;
        src21 <= 16'ha426;
        src22 <= 16'hb55a;
        src23 <= 16'hd403;
        src24 <= 16'hd29c;
        src25 <= 16'h4004;
        src26 <= 16'h76fe;
        src27 <= 16'he88b;
        src28 <= 16'h5ff8;
        src29 <= 16'hd523;
        src30 <= 16'hb6a2;
        src31 <= 16'hba0;
        src32 <= 16'h7f3c;
        src33 <= 16'hf6ac;
        src34 <= 16'h1ff6;
        src35 <= 16'hf7bb;
        src36 <= 16'h9749;
        src37 <= 16'h994d;
        src38 <= 16'hbedc;
        src39 <= 16'h1620;
        src40 <= 16'he867;
        src41 <= 16'hf5cb;
        src42 <= 16'h9020;
        src43 <= 16'ha9eb;
        src44 <= 16'h5935;
        src45 <= 16'h7ab0;
        src46 <= 16'h8cc2;
        src47 <= 16'ha04f;
        src48 <= 16'h2491;
        src49 <= 16'hd6ee;
        src50 <= 16'h61f1;
        src51 <= 16'h31ed;
        src52 <= 16'h8306;
        src53 <= 16'he777;
        exp <= 22'h1f5943;
        #1
        src0 <= 16'hde3c;
        src1 <= 16'hc4d4;
        src2 <= 16'h9394;
        src3 <= 16'h7fbe;
        src4 <= 16'h84ae;
        src5 <= 16'hc00d;
        src6 <= 16'hf17d;
        src7 <= 16'hc4b0;
        src8 <= 16'hbf25;
        src9 <= 16'hb956;
        src10 <= 16'hfb2f;
        src11 <= 16'h975a;
        src12 <= 16'hf9de;
        src13 <= 16'he56d;
        src14 <= 16'h6e6d;
        src15 <= 16'he9de;
        src16 <= 16'h3a94;
        src17 <= 16'h5df0;
        src18 <= 16'hac99;
        src19 <= 16'hf2b;
        src20 <= 16'hb134;
        src21 <= 16'hd8a6;
        src22 <= 16'h1ec8;
        src23 <= 16'h5757;
        src24 <= 16'h368e;
        src25 <= 16'hd476;
        src26 <= 16'ha57f;
        src27 <= 16'h1138;
        src28 <= 16'hbf49;
        src29 <= 16'h6392;
        src30 <= 16'h89b;
        src31 <= 16'h627f;
        src32 <= 16'h626;
        src33 <= 16'h8827;
        src34 <= 16'h867c;
        src35 <= 16'hdf31;
        src36 <= 16'h72df;
        src37 <= 16'ha4d9;
        src38 <= 16'h13c2;
        src39 <= 16'h3aad;
        src40 <= 16'h3faf;
        src41 <= 16'hc7c5;
        src42 <= 16'h4261;
        src43 <= 16'h4ca0;
        src44 <= 16'h879c;
        src45 <= 16'hb510;
        src46 <= 16'h980c;
        src47 <= 16'h4721;
        src48 <= 16'hcae1;
        src49 <= 16'he9b8;
        src50 <= 16'hda43;
        src51 <= 16'h7b30;
        src52 <= 16'h71e9;
        src53 <= 16'h1093;
        exp <= 22'h1d30cc;
        #1
        src0 <= 16'h383;
        src1 <= 16'hc0c5;
        src2 <= 16'hc22;
        src3 <= 16'h74f0;
        src4 <= 16'h1014;
        src5 <= 16'h206b;
        src6 <= 16'h8de9;
        src7 <= 16'h1f59;
        src8 <= 16'hcce;
        src9 <= 16'ha22;
        src10 <= 16'h6ac2;
        src11 <= 16'hf579;
        src12 <= 16'h7eb5;
        src13 <= 16'h5756;
        src14 <= 16'h2a06;
        src15 <= 16'ha54c;
        src16 <= 16'h3832;
        src17 <= 16'hb7b4;
        src18 <= 16'h5025;
        src19 <= 16'h5ab0;
        src20 <= 16'hc194;
        src21 <= 16'hf4c0;
        src22 <= 16'hf84b;
        src23 <= 16'hd59f;
        src24 <= 16'hd2c3;
        src25 <= 16'h83e;
        src26 <= 16'ha7cf;
        src27 <= 16'hb509;
        src28 <= 16'h120b;
        src29 <= 16'h55a3;
        src30 <= 16'he154;
        src31 <= 16'ha85c;
        src32 <= 16'h3fb8;
        src33 <= 16'hca9;
        src34 <= 16'h515a;
        src35 <= 16'hb13d;
        src36 <= 16'h79aa;
        src37 <= 16'h4890;
        src38 <= 16'h433c;
        src39 <= 16'h7737;
        src40 <= 16'h67c3;
        src41 <= 16'ha6b7;
        src42 <= 16'he6ac;
        src43 <= 16'hcb92;
        src44 <= 16'he83f;
        src45 <= 16'hc5be;
        src46 <= 16'h9021;
        src47 <= 16'hfb46;
        src48 <= 16'hfb31;
        src49 <= 16'h179f;
        src50 <= 16'h3da;
        src51 <= 16'h5cee;
        src52 <= 16'hdf46;
        src53 <= 16'h4020;
        exp <= 22'h19e092;
        #1
        src0 <= 16'hb96b;
        src1 <= 16'h3184;
        src2 <= 16'h1b13;
        src3 <= 16'hf85a;
        src4 <= 16'h7ceb;
        src5 <= 16'h8471;
        src6 <= 16'he36a;
        src7 <= 16'h9395;
        src8 <= 16'hc65f;
        src9 <= 16'h8642;
        src10 <= 16'h81ee;
        src11 <= 16'hcd6b;
        src12 <= 16'h5a64;
        src13 <= 16'hd6bc;
        src14 <= 16'h2247;
        src15 <= 16'h3aad;
        src16 <= 16'h1896;
        src17 <= 16'hffb7;
        src18 <= 16'h483;
        src19 <= 16'h58d8;
        src20 <= 16'hfe89;
        src21 <= 16'h4a10;
        src22 <= 16'h441e;
        src23 <= 16'h6eaa;
        src24 <= 16'hab9e;
        src25 <= 16'h2e60;
        src26 <= 16'h3986;
        src27 <= 16'h5500;
        src28 <= 16'hc855;
        src29 <= 16'h2469;
        src30 <= 16'hec21;
        src31 <= 16'h56fc;
        src32 <= 16'hb9de;
        src33 <= 16'h20f4;
        src34 <= 16'h39e0;
        src35 <= 16'h22d8;
        src36 <= 16'h4071;
        src37 <= 16'h58fa;
        src38 <= 16'h7c22;
        src39 <= 16'h7c18;
        src40 <= 16'h75f8;
        src41 <= 16'ha771;
        src42 <= 16'h3727;
        src43 <= 16'ha6d2;
        src44 <= 16'hbc22;
        src45 <= 16'h8e77;
        src46 <= 16'hedaa;
        src47 <= 16'h8a72;
        src48 <= 16'h1e4b;
        src49 <= 16'h1eaa;
        src50 <= 16'h419d;
        src51 <= 16'h8ab2;
        src52 <= 16'hf28e;
        src53 <= 16'ha5cf;
        exp <= 22'h19d314;
        #1
        src0 <= 16'h9130;
        src1 <= 16'hc7f;
        src2 <= 16'hbb08;
        src3 <= 16'hc550;
        src4 <= 16'h1086;
        src5 <= 16'he377;
        src6 <= 16'h288d;
        src7 <= 16'hd354;
        src8 <= 16'hd5a4;
        src9 <= 16'hdc01;
        src10 <= 16'h6012;
        src11 <= 16'he88a;
        src12 <= 16'h5790;
        src13 <= 16'h3781;
        src14 <= 16'h4f83;
        src15 <= 16'hb8ce;
        src16 <= 16'h62a;
        src17 <= 16'h8de6;
        src18 <= 16'heb8c;
        src19 <= 16'h1d4e;
        src20 <= 16'h2061;
        src21 <= 16'hb64a;
        src22 <= 16'h3274;
        src23 <= 16'h761c;
        src24 <= 16'he16;
        src25 <= 16'hae32;
        src26 <= 16'h73dc;
        src27 <= 16'h3db4;
        src28 <= 16'h1d67;
        src29 <= 16'h5066;
        src30 <= 16'he814;
        src31 <= 16'h111c;
        src32 <= 16'h96fa;
        src33 <= 16'h5d7b;
        src34 <= 16'heb94;
        src35 <= 16'h9ab8;
        src36 <= 16'h9779;
        src37 <= 16'h9d20;
        src38 <= 16'hdbf4;
        src39 <= 16'hb5e;
        src40 <= 16'h64ee;
        src41 <= 16'hfc16;
        src42 <= 16'h1ba6;
        src43 <= 16'h5e0a;
        src44 <= 16'h5ee0;
        src45 <= 16'h6851;
        src46 <= 16'hb702;
        src47 <= 16'h6b7e;
        src48 <= 16'h2963;
        src49 <= 16'h854d;
        src50 <= 16'h8b3e;
        src51 <= 16'h1b44;
        src52 <= 16'h9bd1;
        src53 <= 16'h6534;
        exp <= 22'h1941ca;
        #1
        src0 <= 16'h9626;
        src1 <= 16'hf803;
        src2 <= 16'h47bd;
        src3 <= 16'h3f1;
        src4 <= 16'h4929;
        src5 <= 16'hbaa7;
        src6 <= 16'h18b4;
        src7 <= 16'h72a6;
        src8 <= 16'h6432;
        src9 <= 16'h5421;
        src10 <= 16'hc41c;
        src11 <= 16'h69d4;
        src12 <= 16'h8a4d;
        src13 <= 16'h245b;
        src14 <= 16'h728b;
        src15 <= 16'h3d78;
        src16 <= 16'h4b20;
        src17 <= 16'hf973;
        src18 <= 16'hc5f;
        src19 <= 16'hcc84;
        src20 <= 16'h7509;
        src21 <= 16'hb67a;
        src22 <= 16'h2e6e;
        src23 <= 16'hb90f;
        src24 <= 16'h24fc;
        src25 <= 16'h65d9;
        src26 <= 16'h2475;
        src27 <= 16'h2ec5;
        src28 <= 16'h1aa0;
        src29 <= 16'h3ec8;
        src30 <= 16'h5c2d;
        src31 <= 16'had9d;
        src32 <= 16'h526;
        src33 <= 16'h161e;
        src34 <= 16'hbaf0;
        src35 <= 16'h6db0;
        src36 <= 16'haa49;
        src37 <= 16'h62cb;
        src38 <= 16'h2bf9;
        src39 <= 16'h1f5;
        src40 <= 16'hb0c3;
        src41 <= 16'h194c;
        src42 <= 16'hc2c7;
        src43 <= 16'h7249;
        src44 <= 16'h460e;
        src45 <= 16'h3869;
        src46 <= 16'h245a;
        src47 <= 16'hcfeb;
        src48 <= 16'h9202;
        src49 <= 16'h356a;
        src50 <= 16'h410b;
        src51 <= 16'h4a59;
        src52 <= 16'h438b;
        src53 <= 16'h7ddf;
        exp <= 22'h1524a1;
        #1
        src0 <= 16'h67e9;
        src1 <= 16'h8204;
        src2 <= 16'h839f;
        src3 <= 16'hde86;
        src4 <= 16'hb385;
        src5 <= 16'hfbd9;
        src6 <= 16'he792;
        src7 <= 16'hb8ad;
        src8 <= 16'h67d0;
        src9 <= 16'ha710;
        src10 <= 16'h5a3;
        src11 <= 16'hc44c;
        src12 <= 16'h613c;
        src13 <= 16'h90b9;
        src14 <= 16'h68a7;
        src15 <= 16'hb0b1;
        src16 <= 16'h43f8;
        src17 <= 16'hdb3f;
        src18 <= 16'hd790;
        src19 <= 16'hbf67;
        src20 <= 16'hbdfb;
        src21 <= 16'h9476;
        src22 <= 16'h9af7;
        src23 <= 16'h6754;
        src24 <= 16'hf5f4;
        src25 <= 16'h2921;
        src26 <= 16'h3f44;
        src27 <= 16'h926a;
        src28 <= 16'hc9ae;
        src29 <= 16'h4469;
        src30 <= 16'h547c;
        src31 <= 16'h248a;
        src32 <= 16'h48d6;
        src33 <= 16'hf333;
        src34 <= 16'h13b;
        src35 <= 16'h2095;
        src36 <= 16'hdf0f;
        src37 <= 16'h233f;
        src38 <= 16'h8d5d;
        src39 <= 16'h4471;
        src40 <= 16'h7c3;
        src41 <= 16'h7a15;
        src42 <= 16'h9939;
        src43 <= 16'hae87;
        src44 <= 16'hf18b;
        src45 <= 16'ha6fa;
        src46 <= 16'h38fc;
        src47 <= 16'h400f;
        src48 <= 16'h2af0;
        src49 <= 16'h572f;
        src50 <= 16'h4044;
        src51 <= 16'h25a8;
        src52 <= 16'h6c6d;
        src53 <= 16'hfbac;
        exp <= 22'h1b5fd6;
        #1
        src0 <= 16'hb074;
        src1 <= 16'h7bfb;
        src2 <= 16'hd861;
        src3 <= 16'h1bd8;
        src4 <= 16'h6746;
        src5 <= 16'h7ee3;
        src6 <= 16'had6f;
        src7 <= 16'ha2b0;
        src8 <= 16'h189d;
        src9 <= 16'h7dbc;
        src10 <= 16'h8767;
        src11 <= 16'h713b;
        src12 <= 16'hc161;
        src13 <= 16'h81b8;
        src14 <= 16'h21b2;
        src15 <= 16'hec0a;
        src16 <= 16'h1999;
        src17 <= 16'h6064;
        src18 <= 16'h6e61;
        src19 <= 16'hdfe3;
        src20 <= 16'h5c7b;
        src21 <= 16'hef70;
        src22 <= 16'ha25e;
        src23 <= 16'h3b4e;
        src24 <= 16'h81d3;
        src25 <= 16'h25f2;
        src26 <= 16'h77ab;
        src27 <= 16'haa08;
        src28 <= 16'h6ea9;
        src29 <= 16'h20ad;
        src30 <= 16'haa17;
        src31 <= 16'hb276;
        src32 <= 16'hf93b;
        src33 <= 16'h25fa;
        src34 <= 16'h15b6;
        src35 <= 16'h9a15;
        src36 <= 16'h5255;
        src37 <= 16'hef24;
        src38 <= 16'h667b;
        src39 <= 16'haf0b;
        src40 <= 16'h1392;
        src41 <= 16'h4bfc;
        src42 <= 16'h5ff5;
        src43 <= 16'h87f5;
        src44 <= 16'h35b9;
        src45 <= 16'h23c8;
        src46 <= 16'h2340;
        src47 <= 16'hbfb8;
        src48 <= 16'h61d6;
        src49 <= 16'he951;
        src50 <= 16'he7ff;
        src51 <= 16'h4406;
        src52 <= 16'h735f;
        src53 <= 16'h204c;
        exp <= 22'h1992ba;
        #1
        src0 <= 16'hcdd6;
        src1 <= 16'h54a9;
        src2 <= 16'h25d4;
        src3 <= 16'ha5ab;
        src4 <= 16'h48fd;
        src5 <= 16'h81b;
        src6 <= 16'ha583;
        src7 <= 16'hee24;
        src8 <= 16'hb69d;
        src9 <= 16'h6500;
        src10 <= 16'he46;
        src11 <= 16'ha39f;
        src12 <= 16'h944;
        src13 <= 16'hf0d4;
        src14 <= 16'h2431;
        src15 <= 16'h54b1;
        src16 <= 16'h8cda;
        src17 <= 16'h34c1;
        src18 <= 16'hd872;
        src19 <= 16'hd3b4;
        src20 <= 16'h21e;
        src21 <= 16'h9c80;
        src22 <= 16'haed2;
        src23 <= 16'h2ae8;
        src24 <= 16'hbf0c;
        src25 <= 16'h4870;
        src26 <= 16'ha902;
        src27 <= 16'heb07;
        src28 <= 16'h12bd;
        src29 <= 16'hb6ed;
        src30 <= 16'hc92c;
        src31 <= 16'hfa2a;
        src32 <= 16'ha35;
        src33 <= 16'h9f74;
        src34 <= 16'h6683;
        src35 <= 16'hf89c;
        src36 <= 16'heb15;
        src37 <= 16'hd579;
        src38 <= 16'h64a1;
        src39 <= 16'hd6a5;
        src40 <= 16'h43bd;
        src41 <= 16'h2124;
        src42 <= 16'hb6fb;
        src43 <= 16'h343c;
        src44 <= 16'h72c4;
        src45 <= 16'h57;
        src46 <= 16'hab9f;
        src47 <= 16'ha4aa;
        src48 <= 16'h8656;
        src49 <= 16'h4c5d;
        src50 <= 16'hacec;
        src51 <= 16'hf833;
        src52 <= 16'h8f56;
        src53 <= 16'hc986;
        exp <= 22'h1c0a9d;
        #1
        src0 <= 16'h6efd;
        src1 <= 16'h27ce;
        src2 <= 16'h80ae;
        src3 <= 16'hcb74;
        src4 <= 16'h5738;
        src5 <= 16'h9075;
        src6 <= 16'hb9a0;
        src7 <= 16'h8b9d;
        src8 <= 16'h3725;
        src9 <= 16'h2e4e;
        src10 <= 16'h1828;
        src11 <= 16'h38a4;
        src12 <= 16'h36d2;
        src13 <= 16'h4d8b;
        src14 <= 16'h697e;
        src15 <= 16'he10d;
        src16 <= 16'hfbfa;
        src17 <= 16'h716b;
        src18 <= 16'hb062;
        src19 <= 16'h2605;
        src20 <= 16'h5657;
        src21 <= 16'h18d6;
        src22 <= 16'hb64c;
        src23 <= 16'h57ed;
        src24 <= 16'h442c;
        src25 <= 16'h3670;
        src26 <= 16'hb763;
        src27 <= 16'h23b0;
        src28 <= 16'hb9c7;
        src29 <= 16'h6989;
        src30 <= 16'h9206;
        src31 <= 16'habf8;
        src32 <= 16'hc345;
        src33 <= 16'h91f8;
        src34 <= 16'h157e;
        src35 <= 16'h41b3;
        src36 <= 16'h54f2;
        src37 <= 16'h8a64;
        src38 <= 16'hbd43;
        src39 <= 16'hb3e5;
        src40 <= 16'h55d5;
        src41 <= 16'h7193;
        src42 <= 16'hae92;
        src43 <= 16'hbed6;
        src44 <= 16'h5119;
        src45 <= 16'hf92;
        src46 <= 16'h93cd;
        src47 <= 16'h55e8;
        src48 <= 16'hab29;
        src49 <= 16'hbf5b;
        src50 <= 16'hbb06;
        src51 <= 16'h8151;
        src52 <= 16'h859;
        src53 <= 16'h399e;
        exp <= 22'h18721b;
        #1
        src0 <= 16'hdac8;
        src1 <= 16'hde95;
        src2 <= 16'h2693;
        src3 <= 16'h2bfb;
        src4 <= 16'haf06;
        src5 <= 16'h16e6;
        src6 <= 16'h2788;
        src7 <= 16'hd26e;
        src8 <= 16'h39f7;
        src9 <= 16'h705d;
        src10 <= 16'hdfa5;
        src11 <= 16'hcf1d;
        src12 <= 16'he52b;
        src13 <= 16'h175f;
        src14 <= 16'he5;
        src15 <= 16'h49ae;
        src16 <= 16'h957;
        src17 <= 16'h807;
        src18 <= 16'ha536;
        src19 <= 16'h524a;
        src20 <= 16'h60df;
        src21 <= 16'h64f5;
        src22 <= 16'h3780;
        src23 <= 16'h47cf;
        src24 <= 16'hc0b6;
        src25 <= 16'he251;
        src26 <= 16'h8730;
        src27 <= 16'hda4d;
        src28 <= 16'h62ef;
        src29 <= 16'ha0a0;
        src30 <= 16'h57f;
        src31 <= 16'h8a86;
        src32 <= 16'h310f;
        src33 <= 16'hf8ba;
        src34 <= 16'ha3c0;
        src35 <= 16'h9238;
        src36 <= 16'h89cf;
        src37 <= 16'h288c;
        src38 <= 16'h63ce;
        src39 <= 16'h415c;
        src40 <= 16'hfe31;
        src41 <= 16'h965b;
        src42 <= 16'h3753;
        src43 <= 16'h80b9;
        src44 <= 16'hd047;
        src45 <= 16'hbb56;
        src46 <= 16'h67ee;
        src47 <= 16'hf714;
        src48 <= 16'h21cd;
        src49 <= 16'h3437;
        src50 <= 16'hbdf4;
        src51 <= 16'h87af;
        src52 <= 16'he1e5;
        src53 <= 16'h69ff;
        exp <= 22'h1a2821;
        #1
        src0 <= 16'h23c3;
        src1 <= 16'h6b80;
        src2 <= 16'h93c;
        src3 <= 16'hdc94;
        src4 <= 16'hd8b4;
        src5 <= 16'hb5eb;
        src6 <= 16'hd7b7;
        src7 <= 16'h46de;
        src8 <= 16'h6875;
        src9 <= 16'hf93e;
        src10 <= 16'h703b;
        src11 <= 16'h16da;
        src12 <= 16'h66cd;
        src13 <= 16'hf48e;
        src14 <= 16'h23c4;
        src15 <= 16'h9b3;
        src16 <= 16'hed4a;
        src17 <= 16'ha454;
        src18 <= 16'ha9f4;
        src19 <= 16'hf952;
        src20 <= 16'hba8e;
        src21 <= 16'h4f95;
        src22 <= 16'he130;
        src23 <= 16'h962a;
        src24 <= 16'h9ee4;
        src25 <= 16'h2531;
        src26 <= 16'h23f0;
        src27 <= 16'hfb4c;
        src28 <= 16'hbd12;
        src29 <= 16'ha316;
        src30 <= 16'h9c7f;
        src31 <= 16'hf636;
        src32 <= 16'hf5d7;
        src33 <= 16'h337c;
        src34 <= 16'h649f;
        src35 <= 16'he1ce;
        src36 <= 16'h3dda;
        src37 <= 16'h2c48;
        src38 <= 16'hf7de;
        src39 <= 16'hfbbd;
        src40 <= 16'h7992;
        src41 <= 16'h39b8;
        src42 <= 16'h1edd;
        src43 <= 16'h77d3;
        src44 <= 16'hd9e4;
        src45 <= 16'h196b;
        src46 <= 16'hfb3e;
        src47 <= 16'ha2fe;
        src48 <= 16'h3e14;
        src49 <= 16'h14cd;
        src50 <= 16'he3a8;
        src51 <= 16'he119;
        src52 <= 16'h9743;
        src53 <= 16'hc724;
        exp <= 22'h1e3f7b;
        #1
        src0 <= 16'h4121;
        src1 <= 16'h87f5;
        src2 <= 16'h748d;
        src3 <= 16'h96be;
        src4 <= 16'h230d;
        src5 <= 16'h6bdf;
        src6 <= 16'h6adf;
        src7 <= 16'h87a4;
        src8 <= 16'h771a;
        src9 <= 16'he98e;
        src10 <= 16'hd59a;
        src11 <= 16'hb02a;
        src12 <= 16'h901e;
        src13 <= 16'h1ada;
        src14 <= 16'h660e;
        src15 <= 16'h276;
        src16 <= 16'hb6b6;
        src17 <= 16'hcff0;
        src18 <= 16'hba4a;
        src19 <= 16'h24b8;
        src20 <= 16'hbe5c;
        src21 <= 16'hf50;
        src22 <= 16'h5ae8;
        src23 <= 16'h7b38;
        src24 <= 16'h86c3;
        src25 <= 16'heb0;
        src26 <= 16'h8a10;
        src27 <= 16'h27eb;
        src28 <= 16'h625d;
        src29 <= 16'h157c;
        src30 <= 16'h41af;
        src31 <= 16'h349f;
        src32 <= 16'haf88;
        src33 <= 16'hf489;
        src34 <= 16'hbe42;
        src35 <= 16'h5205;
        src36 <= 16'hf096;
        src37 <= 16'hab41;
        src38 <= 16'hd6a4;
        src39 <= 16'he693;
        src40 <= 16'h707c;
        src41 <= 16'hbc95;
        src42 <= 16'h145d;
        src43 <= 16'hb03c;
        src44 <= 16'hc11d;
        src45 <= 16'h8299;
        src46 <= 16'h1199;
        src47 <= 16'h3c05;
        src48 <= 16'h2b7b;
        src49 <= 16'he6cb;
        src50 <= 16'he489;
        src51 <= 16'h3c7c;
        src52 <= 16'h61f4;
        src53 <= 16'h79eb;
        exp <= 22'h1a2e4f;
        #1
        src0 <= 16'h7d01;
        src1 <= 16'hdda5;
        src2 <= 16'hd06f;
        src3 <= 16'hff4d;
        src4 <= 16'h9016;
        src5 <= 16'h3068;
        src6 <= 16'h6ae8;
        src7 <= 16'hec4f;
        src8 <= 16'h9f0c;
        src9 <= 16'h98cd;
        src10 <= 16'hffaa;
        src11 <= 16'hcb02;
        src12 <= 16'h48d0;
        src13 <= 16'h487b;
        src14 <= 16'hb856;
        src15 <= 16'hacdc;
        src16 <= 16'h250f;
        src17 <= 16'h539e;
        src18 <= 16'haff4;
        src19 <= 16'hb5d5;
        src20 <= 16'hbf0c;
        src21 <= 16'h9e08;
        src22 <= 16'hc4fa;
        src23 <= 16'he1ec;
        src24 <= 16'h9996;
        src25 <= 16'hbb9f;
        src26 <= 16'ha9be;
        src27 <= 16'hb471;
        src28 <= 16'h558e;
        src29 <= 16'h445c;
        src30 <= 16'h1ee8;
        src31 <= 16'h3222;
        src32 <= 16'hf491;
        src33 <= 16'h7806;
        src34 <= 16'h1d87;
        src35 <= 16'h36fa;
        src36 <= 16'h2708;
        src37 <= 16'h26e6;
        src38 <= 16'h9512;
        src39 <= 16'he80f;
        src40 <= 16'h9d6d;
        src41 <= 16'ha14e;
        src42 <= 16'h76d3;
        src43 <= 16'he409;
        src44 <= 16'h1184;
        src45 <= 16'h6f08;
        src46 <= 16'he532;
        src47 <= 16'h5da;
        src48 <= 16'hc270;
        src49 <= 16'h1b76;
        src50 <= 16'hc51;
        src51 <= 16'hdb77;
        src52 <= 16'he338;
        src53 <= 16'h427e;
        exp <= 22'h1d389b;
        #1
        src0 <= 16'hff14;
        src1 <= 16'h37a2;
        src2 <= 16'hdbfc;
        src3 <= 16'h447c;
        src4 <= 16'h7968;
        src5 <= 16'hd9d6;
        src6 <= 16'h9bf4;
        src7 <= 16'h2e75;
        src8 <= 16'hfe4e;
        src9 <= 16'hf9ff;
        src10 <= 16'hdcea;
        src11 <= 16'h1a4e;
        src12 <= 16'ha847;
        src13 <= 16'hb9d1;
        src14 <= 16'hae2a;
        src15 <= 16'hd95c;
        src16 <= 16'h5393;
        src17 <= 16'h796e;
        src18 <= 16'h1048;
        src19 <= 16'h5715;
        src20 <= 16'ha46d;
        src21 <= 16'h49ae;
        src22 <= 16'hc447;
        src23 <= 16'h2fa8;
        src24 <= 16'hed52;
        src25 <= 16'h67ed;
        src26 <= 16'h471d;
        src27 <= 16'h905c;
        src28 <= 16'h3760;
        src29 <= 16'h5f38;
        src30 <= 16'h40a2;
        src31 <= 16'h3ccf;
        src32 <= 16'hd298;
        src33 <= 16'h220f;
        src34 <= 16'h9085;
        src35 <= 16'hd68a;
        src36 <= 16'h7194;
        src37 <= 16'he5aa;
        src38 <= 16'hc84;
        src39 <= 16'h6678;
        src40 <= 16'hb83c;
        src41 <= 16'ha906;
        src42 <= 16'h1bb8;
        src43 <= 16'h3080;
        src44 <= 16'hd983;
        src45 <= 16'hff4d;
        src46 <= 16'hf7f0;
        src47 <= 16'h3bfc;
        src48 <= 16'h89e8;
        src49 <= 16'he9db;
        src50 <= 16'ha44b;
        src51 <= 16'h8f4;
        src52 <= 16'he2a5;
        src53 <= 16'h2829;
        exp <= 22'h1cb117;
        #1
        src0 <= 16'h31f7;
        src1 <= 16'h6140;
        src2 <= 16'hf2d5;
        src3 <= 16'h593d;
        src4 <= 16'he553;
        src5 <= 16'h588;
        src6 <= 16'hac16;
        src7 <= 16'hf001;
        src8 <= 16'h7d85;
        src9 <= 16'h644d;
        src10 <= 16'hf506;
        src11 <= 16'h3039;
        src12 <= 16'h8797;
        src13 <= 16'h4ac2;
        src14 <= 16'h8ed3;
        src15 <= 16'h48b6;
        src16 <= 16'h38b5;
        src17 <= 16'h8abb;
        src18 <= 16'h34b8;
        src19 <= 16'hd337;
        src20 <= 16'h395e;
        src21 <= 16'h81bd;
        src22 <= 16'hc2c9;
        src23 <= 16'h8533;
        src24 <= 16'h2709;
        src25 <= 16'h7913;
        src26 <= 16'hca06;
        src27 <= 16'hb02a;
        src28 <= 16'hd3cd;
        src29 <= 16'h6a3;
        src30 <= 16'hed05;
        src31 <= 16'ha510;
        src32 <= 16'h96bb;
        src33 <= 16'hf581;
        src34 <= 16'hb733;
        src35 <= 16'hef89;
        src36 <= 16'hdf8b;
        src37 <= 16'h8968;
        src38 <= 16'h2f94;
        src39 <= 16'h857a;
        src40 <= 16'haf10;
        src41 <= 16'heff0;
        src42 <= 16'ha302;
        src43 <= 16'hc471;
        src44 <= 16'hb201;
        src45 <= 16'h640e;
        src46 <= 16'h1149;
        src47 <= 16'h4baf;
        src48 <= 16'h6b12;
        src49 <= 16'h4e64;
        src50 <= 16'h9e8d;
        src51 <= 16'h1c37;
        src52 <= 16'hbb18;
        src53 <= 16'hb3a4;
        exp <= 22'h1d19de;
        #1
        src0 <= 16'h1b92;
        src1 <= 16'h83b1;
        src2 <= 16'h4d98;
        src3 <= 16'h310b;
        src4 <= 16'h40b1;
        src5 <= 16'h886e;
        src6 <= 16'ha2f0;
        src7 <= 16'h464f;
        src8 <= 16'hd1f0;
        src9 <= 16'h6b4e;
        src10 <= 16'h1e67;
        src11 <= 16'hc7cd;
        src12 <= 16'h4ead;
        src13 <= 16'h9b9;
        src14 <= 16'h7f07;
        src15 <= 16'h57f6;
        src16 <= 16'h9383;
        src17 <= 16'h917f;
        src18 <= 16'h4395;
        src19 <= 16'h2ba0;
        src20 <= 16'h3e21;
        src21 <= 16'h254;
        src22 <= 16'he15f;
        src23 <= 16'h910b;
        src24 <= 16'ha1a4;
        src25 <= 16'hd9e0;
        src26 <= 16'hc958;
        src27 <= 16'h4fbd;
        src28 <= 16'h93ec;
        src29 <= 16'h50d4;
        src30 <= 16'h5a72;
        src31 <= 16'h77cc;
        src32 <= 16'h27d4;
        src33 <= 16'h30a4;
        src34 <= 16'h23c6;
        src35 <= 16'h6296;
        src36 <= 16'h4d88;
        src37 <= 16'h443f;
        src38 <= 16'hdd24;
        src39 <= 16'haa3;
        src40 <= 16'h2923;
        src41 <= 16'h5748;
        src42 <= 16'h3e8;
        src43 <= 16'h9a13;
        src44 <= 16'hd2;
        src45 <= 16'hf51a;
        src46 <= 16'hb95a;
        src47 <= 16'hf9f4;
        src48 <= 16'h7392;
        src49 <= 16'h57da;
        src50 <= 16'h8f04;
        src51 <= 16'hb34c;
        src52 <= 16'h44f;
        src53 <= 16'hfc4a;
        exp <= 22'h16e41d;
        #1
        src0 <= 16'h574c;
        src1 <= 16'h39ad;
        src2 <= 16'h72ad;
        src3 <= 16'h6bdb;
        src4 <= 16'hc9f4;
        src5 <= 16'ha995;
        src6 <= 16'hf695;
        src7 <= 16'h17c8;
        src8 <= 16'h41d2;
        src9 <= 16'hd4f7;
        src10 <= 16'hf239;
        src11 <= 16'hc82c;
        src12 <= 16'h6fc5;
        src13 <= 16'h21a2;
        src14 <= 16'h954c;
        src15 <= 16'hb87e;
        src16 <= 16'hbe3a;
        src17 <= 16'hca37;
        src18 <= 16'he026;
        src19 <= 16'hcadb;
        src20 <= 16'ha2cf;
        src21 <= 16'hf1c9;
        src22 <= 16'he5dd;
        src23 <= 16'hda8a;
        src24 <= 16'hc4b7;
        src25 <= 16'hfb94;
        src26 <= 16'hbf88;
        src27 <= 16'hfa2f;
        src28 <= 16'h6ab7;
        src29 <= 16'h60c1;
        src30 <= 16'hbff4;
        src31 <= 16'hd2ce;
        src32 <= 16'he75a;
        src33 <= 16'hdc01;
        src34 <= 16'h9377;
        src35 <= 16'h3f88;
        src36 <= 16'h3328;
        src37 <= 16'h9703;
        src38 <= 16'h4462;
        src39 <= 16'h6cd8;
        src40 <= 16'h7ae4;
        src41 <= 16'h29ac;
        src42 <= 16'hd875;
        src43 <= 16'hc41f;
        src44 <= 16'hdb22;
        src45 <= 16'hbeba;
        src46 <= 16'h4e;
        src47 <= 16'he942;
        src48 <= 16'hab75;
        src49 <= 16'h1f1c;
        src50 <= 16'h9ac6;
        src51 <= 16'he9d2;
        src52 <= 16'h7ed5;
        src53 <= 16'h6793;
        exp <= 22'h210e53;
        #1
        src0 <= 16'h29fd;
        src1 <= 16'hf2e3;
        src2 <= 16'h1aca;
        src3 <= 16'h2b6f;
        src4 <= 16'h8001;
        src5 <= 16'haa4a;
        src6 <= 16'h6d78;
        src7 <= 16'h8e80;
        src8 <= 16'hb9e;
        src9 <= 16'hf67b;
        src10 <= 16'hc823;
        src11 <= 16'h3fdc;
        src12 <= 16'hd8a7;
        src13 <= 16'h4ac8;
        src14 <= 16'h5f17;
        src15 <= 16'h226b;
        src16 <= 16'h1655;
        src17 <= 16'hc3b1;
        src18 <= 16'h5ee1;
        src19 <= 16'h1ae0;
        src20 <= 16'h3096;
        src21 <= 16'hd8f;
        src22 <= 16'hd5ad;
        src23 <= 16'hcbf1;
        src24 <= 16'he265;
        src25 <= 16'h387d;
        src26 <= 16'h86b;
        src27 <= 16'ha31;
        src28 <= 16'he9fb;
        src29 <= 16'hcfab;
        src30 <= 16'h32b2;
        src31 <= 16'h14f3;
        src32 <= 16'hb496;
        src33 <= 16'h2bc6;
        src34 <= 16'h99e;
        src35 <= 16'hf2f5;
        src36 <= 16'h1c1d;
        src37 <= 16'h4147;
        src38 <= 16'h570b;
        src39 <= 16'hbe4b;
        src40 <= 16'hfdb;
        src41 <= 16'h6137;
        src42 <= 16'h4d6d;
        src43 <= 16'hd1ba;
        src44 <= 16'h1e19;
        src45 <= 16'hd9cb;
        src46 <= 16'h41a0;
        src47 <= 16'h7635;
        src48 <= 16'h7e17;
        src49 <= 16'h1f25;
        src50 <= 16'hcd43;
        src51 <= 16'h1cc1;
        src52 <= 16'h433f;
        src53 <= 16'h7fee;
        exp <= 22'h1674c0;
        #1
        src0 <= 16'hf5eb;
        src1 <= 16'h9464;
        src2 <= 16'hc12a;
        src3 <= 16'h4cdc;
        src4 <= 16'h2cfe;
        src5 <= 16'h1541;
        src6 <= 16'h3127;
        src7 <= 16'h2caa;
        src8 <= 16'h15dd;
        src9 <= 16'h78b9;
        src10 <= 16'h2901;
        src11 <= 16'h6c38;
        src12 <= 16'h4e85;
        src13 <= 16'h9706;
        src14 <= 16'he92f;
        src15 <= 16'hf47c;
        src16 <= 16'h6509;
        src17 <= 16'h3fc0;
        src18 <= 16'hb744;
        src19 <= 16'h7961;
        src20 <= 16'he06e;
        src21 <= 16'hc3b9;
        src22 <= 16'hfa3e;
        src23 <= 16'hee6d;
        src24 <= 16'hd4c;
        src25 <= 16'hae1;
        src26 <= 16'h5e6b;
        src27 <= 16'h9503;
        src28 <= 16'h451;
        src29 <= 16'hcc9b;
        src30 <= 16'h2266;
        src31 <= 16'hb70f;
        src32 <= 16'h6487;
        src33 <= 16'h1893;
        src34 <= 16'hcc4b;
        src35 <= 16'hff33;
        src36 <= 16'hfbdc;
        src37 <= 16'h7340;
        src38 <= 16'h8b98;
        src39 <= 16'h1515;
        src40 <= 16'hd0e1;
        src41 <= 16'h670;
        src42 <= 16'h53c1;
        src43 <= 16'h7b8d;
        src44 <= 16'h4c1c;
        src45 <= 16'h45c0;
        src46 <= 16'h3cf2;
        src47 <= 16'h6cbc;
        src48 <= 16'h2be7;
        src49 <= 16'h84c2;
        src50 <= 16'h305c;
        src51 <= 16'h459c;
        src52 <= 16'hc718;
        src53 <= 16'haa30;
        exp <= 22'h190a19;
        #1
        src0 <= 16'hc528;
        src1 <= 16'hc6da;
        src2 <= 16'h5c22;
        src3 <= 16'h5395;
        src4 <= 16'h5d5c;
        src5 <= 16'h1274;
        src6 <= 16'hc7f6;
        src7 <= 16'hca15;
        src8 <= 16'hf744;
        src9 <= 16'hf199;
        src10 <= 16'hd03;
        src11 <= 16'haf0d;
        src12 <= 16'h9140;
        src13 <= 16'h1f75;
        src14 <= 16'hb89d;
        src15 <= 16'he3d3;
        src16 <= 16'hda80;
        src17 <= 16'hbae;
        src18 <= 16'hc914;
        src19 <= 16'h18ba;
        src20 <= 16'hb22;
        src21 <= 16'h6f7a;
        src22 <= 16'h3379;
        src23 <= 16'he04;
        src24 <= 16'hc588;
        src25 <= 16'h6765;
        src26 <= 16'h3b0e;
        src27 <= 16'hc74d;
        src28 <= 16'hfaf0;
        src29 <= 16'h34ca;
        src30 <= 16'h1e1;
        src31 <= 16'he394;
        src32 <= 16'h5a19;
        src33 <= 16'h1225;
        src34 <= 16'h3304;
        src35 <= 16'hd325;
        src36 <= 16'h9e3d;
        src37 <= 16'haf99;
        src38 <= 16'h97a8;
        src39 <= 16'he660;
        src40 <= 16'h1eac;
        src41 <= 16'h2f7b;
        src42 <= 16'ha37;
        src43 <= 16'hf3cc;
        src44 <= 16'h508d;
        src45 <= 16'h2207;
        src46 <= 16'h8081;
        src47 <= 16'h82d0;
        src48 <= 16'hddd2;
        src49 <= 16'hbfb4;
        src50 <= 16'h9c65;
        src51 <= 16'hfb56;
        src52 <= 16'h8216;
        src53 <= 16'h6789;
        exp <= 22'h1b1766;
        #1
        src0 <= 16'hc709;
        src1 <= 16'h509e;
        src2 <= 16'hf9fd;
        src3 <= 16'hd39d;
        src4 <= 16'h61e2;
        src5 <= 16'h1d7f;
        src6 <= 16'hc687;
        src7 <= 16'hbe1f;
        src8 <= 16'hbcf4;
        src9 <= 16'hcf6c;
        src10 <= 16'h9c01;
        src11 <= 16'hbee1;
        src12 <= 16'h3b31;
        src13 <= 16'hc5ae;
        src14 <= 16'hd002;
        src15 <= 16'h7919;
        src16 <= 16'hc750;
        src17 <= 16'he36f;
        src18 <= 16'h8974;
        src19 <= 16'hb3a4;
        src20 <= 16'h5b9a;
        src21 <= 16'hea87;
        src22 <= 16'hcef7;
        src23 <= 16'h7d6c;
        src24 <= 16'h34ac;
        src25 <= 16'hcdae;
        src26 <= 16'h8724;
        src27 <= 16'h3e58;
        src28 <= 16'h3cb2;
        src29 <= 16'h4f37;
        src30 <= 16'heb02;
        src31 <= 16'h65a1;
        src32 <= 16'hbce8;
        src33 <= 16'h1e36;
        src34 <= 16'hbc10;
        src35 <= 16'hda63;
        src36 <= 16'h6228;
        src37 <= 16'h7e31;
        src38 <= 16'hf519;
        src39 <= 16'h8480;
        src40 <= 16'h2832;
        src41 <= 16'h1cb8;
        src42 <= 16'hbca7;
        src43 <= 16'hcc1d;
        src44 <= 16'h2478;
        src45 <= 16'he04;
        src46 <= 16'h96a1;
        src47 <= 16'h6a3;
        src48 <= 16'h7345;
        src49 <= 16'h9c12;
        src50 <= 16'hc7e0;
        src51 <= 16'h98cb;
        src52 <= 16'h45d0;
        src53 <= 16'hd534;
        exp <= 22'h1e2d38;
        #1
        src0 <= 16'h7c83;
        src1 <= 16'h6e92;
        src2 <= 16'h6f1c;
        src3 <= 16'hd24b;
        src4 <= 16'h3914;
        src5 <= 16'h2a5b;
        src6 <= 16'h6f67;
        src7 <= 16'hae76;
        src8 <= 16'hf0db;
        src9 <= 16'h561d;
        src10 <= 16'hd0d2;
        src11 <= 16'h1417;
        src12 <= 16'hb1f5;
        src13 <= 16'h920c;
        src14 <= 16'hd4bc;
        src15 <= 16'h1bfd;
        src16 <= 16'h6ef8;
        src17 <= 16'hd3a4;
        src18 <= 16'hbb26;
        src19 <= 16'h43f9;
        src20 <= 16'hbe50;
        src21 <= 16'h4cc;
        src22 <= 16'he513;
        src23 <= 16'h3730;
        src24 <= 16'h3bc9;
        src25 <= 16'h7059;
        src26 <= 16'h1ce6;
        src27 <= 16'h8de;
        src28 <= 16'h2cb5;
        src29 <= 16'h42a7;
        src30 <= 16'hb213;
        src31 <= 16'hf110;
        src32 <= 16'hf928;
        src33 <= 16'he32e;
        src34 <= 16'h8710;
        src35 <= 16'h51ac;
        src36 <= 16'h4ca1;
        src37 <= 16'h311d;
        src38 <= 16'hc907;
        src39 <= 16'hdc19;
        src40 <= 16'hda8a;
        src41 <= 16'hbc64;
        src42 <= 16'h88bf;
        src43 <= 16'h1e90;
        src44 <= 16'h71c0;
        src45 <= 16'heb92;
        src46 <= 16'h2157;
        src47 <= 16'he865;
        src48 <= 16'h37c;
        src49 <= 16'hc61e;
        src50 <= 16'hbc72;
        src51 <= 16'h3075;
        src52 <= 16'h6bd9;
        src53 <= 16'h2992;
        exp <= 22'h1add09;
        #1
        src0 <= 16'hd043;
        src1 <= 16'h2bec;
        src2 <= 16'h47d0;
        src3 <= 16'h94af;
        src4 <= 16'he2c2;
        src5 <= 16'hf41f;
        src6 <= 16'hdaa4;
        src7 <= 16'hff20;
        src8 <= 16'h6f3;
        src9 <= 16'h6a40;
        src10 <= 16'h6d9b;
        src11 <= 16'h662b;
        src12 <= 16'h3e9e;
        src13 <= 16'h76b9;
        src14 <= 16'h5cbf;
        src15 <= 16'h6f00;
        src16 <= 16'h2b2;
        src17 <= 16'h8de;
        src18 <= 16'hd1db;
        src19 <= 16'hc9b7;
        src20 <= 16'hacf4;
        src21 <= 16'h7e9d;
        src22 <= 16'hda2a;
        src23 <= 16'h2fc1;
        src24 <= 16'hf271;
        src25 <= 16'h3bd2;
        src26 <= 16'h50ea;
        src27 <= 16'h3bdc;
        src28 <= 16'hcdc7;
        src29 <= 16'hff24;
        src30 <= 16'h6ab9;
        src31 <= 16'h1491;
        src32 <= 16'h7b04;
        src33 <= 16'ha22e;
        src34 <= 16'hc89d;
        src35 <= 16'h72ba;
        src36 <= 16'hcb00;
        src37 <= 16'h308f;
        src38 <= 16'hffa1;
        src39 <= 16'h6d2c;
        src40 <= 16'hd756;
        src41 <= 16'h3148;
        src42 <= 16'h66e7;
        src43 <= 16'hda9b;
        src44 <= 16'h706c;
        src45 <= 16'h8873;
        src46 <= 16'h8363;
        src47 <= 16'h3bf1;
        src48 <= 16'h117f;
        src49 <= 16'hc745;
        src50 <= 16'h6bc4;
        src51 <= 16'h429f;
        src52 <= 16'h39bc;
        src53 <= 16'hee3a;
        exp <= 22'h1ba593;
        #1
        src0 <= 16'heffc;
        src1 <= 16'h6bbb;
        src2 <= 16'hd646;
        src3 <= 16'h30a1;
        src4 <= 16'h1bb9;
        src5 <= 16'h2df9;
        src6 <= 16'h9f79;
        src7 <= 16'h90f4;
        src8 <= 16'h23ad;
        src9 <= 16'h71a6;
        src10 <= 16'hcbbd;
        src11 <= 16'h4715;
        src12 <= 16'hf57b;
        src13 <= 16'hf4ef;
        src14 <= 16'h7f1;
        src15 <= 16'he98a;
        src16 <= 16'h1224;
        src17 <= 16'heff1;
        src18 <= 16'hb820;
        src19 <= 16'h71eb;
        src20 <= 16'hb47a;
        src21 <= 16'hbd74;
        src22 <= 16'hc1f9;
        src23 <= 16'h4b83;
        src24 <= 16'hd228;
        src25 <= 16'h2bf9;
        src26 <= 16'ha3a9;
        src27 <= 16'hf1e1;
        src28 <= 16'h928a;
        src29 <= 16'hcafe;
        src30 <= 16'hb4f2;
        src31 <= 16'h6ff3;
        src32 <= 16'hfa3f;
        src33 <= 16'he640;
        src34 <= 16'h2c9f;
        src35 <= 16'h6884;
        src36 <= 16'hf3f6;
        src37 <= 16'h6ab9;
        src38 <= 16'h3ff5;
        src39 <= 16'h2f40;
        src40 <= 16'hd388;
        src41 <= 16'hc482;
        src42 <= 16'h43f8;
        src43 <= 16'h8b75;
        src44 <= 16'h912;
        src45 <= 16'h5df8;
        src46 <= 16'hfd46;
        src47 <= 16'hab96;
        src48 <= 16'h7a9b;
        src49 <= 16'hc99f;
        src50 <= 16'ha92d;
        src51 <= 16'h8fad;
        src52 <= 16'h14f0;
        src53 <= 16'hbcc2;
        exp <= 22'h1e2c12;
        #1
        src0 <= 16'hce4b;
        src1 <= 16'hd8e7;
        src2 <= 16'hcec;
        src3 <= 16'ha404;
        src4 <= 16'h94fa;
        src5 <= 16'he07e;
        src6 <= 16'haaac;
        src7 <= 16'h2d96;
        src8 <= 16'hfa3b;
        src9 <= 16'h42b7;
        src10 <= 16'hd897;
        src11 <= 16'hb8fc;
        src12 <= 16'hc41e;
        src13 <= 16'hbcb4;
        src14 <= 16'h8a6d;
        src15 <= 16'h227b;
        src16 <= 16'hff41;
        src17 <= 16'heb4d;
        src18 <= 16'h78fd;
        src19 <= 16'h7d82;
        src20 <= 16'h89cf;
        src21 <= 16'h6557;
        src22 <= 16'hb71e;
        src23 <= 16'h9afa;
        src24 <= 16'h408b;
        src25 <= 16'hcf24;
        src26 <= 16'h1032;
        src27 <= 16'hdaf9;
        src28 <= 16'h2a5;
        src29 <= 16'hdaa6;
        src30 <= 16'ha790;
        src31 <= 16'hdfa9;
        src32 <= 16'h9eb7;
        src33 <= 16'hc31a;
        src34 <= 16'h8572;
        src35 <= 16'h67e2;
        src36 <= 16'he90b;
        src37 <= 16'h5839;
        src38 <= 16'h5a34;
        src39 <= 16'h5c82;
        src40 <= 16'h66ff;
        src41 <= 16'hde50;
        src42 <= 16'h2237;
        src43 <= 16'h80ad;
        src44 <= 16'h7d26;
        src45 <= 16'h3d99;
        src46 <= 16'hc64b;
        src47 <= 16'hef49;
        src48 <= 16'he60f;
        src49 <= 16'h3790;
        src50 <= 16'h662a;
        src51 <= 16'h392e;
        src52 <= 16'h30ee;
        src53 <= 16'h1f5b;
        exp <= 22'h1dd0a9;
        #1
        src0 <= 16'h87e5;
        src1 <= 16'h40;
        src2 <= 16'hb31e;
        src3 <= 16'h8668;
        src4 <= 16'h61ba;
        src5 <= 16'ha9af;
        src6 <= 16'h5f6a;
        src7 <= 16'ha731;
        src8 <= 16'hb8b;
        src9 <= 16'hda1f;
        src10 <= 16'h31d1;
        src11 <= 16'h6c02;
        src12 <= 16'h80d2;
        src13 <= 16'h44a1;
        src14 <= 16'h5ccd;
        src15 <= 16'h641d;
        src16 <= 16'h53d3;
        src17 <= 16'h8be5;
        src18 <= 16'hcbb4;
        src19 <= 16'he308;
        src20 <= 16'h694;
        src21 <= 16'h4c60;
        src22 <= 16'h5d9f;
        src23 <= 16'he995;
        src24 <= 16'h47f0;
        src25 <= 16'h7280;
        src26 <= 16'ha01d;
        src27 <= 16'hef32;
        src28 <= 16'h998c;
        src29 <= 16'hdd6e;
        src30 <= 16'hc71d;
        src31 <= 16'h2e4c;
        src32 <= 16'h5a6c;
        src33 <= 16'hae46;
        src34 <= 16'h7046;
        src35 <= 16'h5fe3;
        src36 <= 16'hb2f3;
        src37 <= 16'h69e3;
        src38 <= 16'ha052;
        src39 <= 16'h61ed;
        src40 <= 16'h5083;
        src41 <= 16'hb385;
        src42 <= 16'h561c;
        src43 <= 16'he6b0;
        src44 <= 16'h385;
        src45 <= 16'hb9f9;
        src46 <= 16'hce81;
        src47 <= 16'hca03;
        src48 <= 16'h5e81;
        src49 <= 16'h62e1;
        src50 <= 16'h9c19;
        src51 <= 16'haa8b;
        src52 <= 16'hfd29;
        src53 <= 16'hd29f;
        exp <= 22'h1c22db;
        #1
        src0 <= 16'h580a;
        src1 <= 16'h898;
        src2 <= 16'h4138;
        src3 <= 16'h584a;
        src4 <= 16'hcc9a;
        src5 <= 16'h44be;
        src6 <= 16'haa61;
        src7 <= 16'hb44e;
        src8 <= 16'hcc91;
        src9 <= 16'h9bf7;
        src10 <= 16'hf208;
        src11 <= 16'h80c;
        src12 <= 16'hc443;
        src13 <= 16'hfa3f;
        src14 <= 16'hed60;
        src15 <= 16'hb1c2;
        src16 <= 16'h82cb;
        src17 <= 16'hae1e;
        src18 <= 16'hf9b9;
        src19 <= 16'h4a50;
        src20 <= 16'he717;
        src21 <= 16'h301b;
        src22 <= 16'hd998;
        src23 <= 16'h21a6;
        src24 <= 16'hada7;
        src25 <= 16'h8fad;
        src26 <= 16'hdb82;
        src27 <= 16'h80a9;
        src28 <= 16'h1695;
        src29 <= 16'h3402;
        src30 <= 16'h1048;
        src31 <= 16'hc63f;
        src32 <= 16'he3aa;
        src33 <= 16'hb0e4;
        src34 <= 16'hbab7;
        src35 <= 16'hbb1e;
        src36 <= 16'h9de4;
        src37 <= 16'hbc8d;
        src38 <= 16'h6dbc;
        src39 <= 16'h1b5d;
        src40 <= 16'hf066;
        src41 <= 16'hc235;
        src42 <= 16'hc8d3;
        src43 <= 16'he592;
        src44 <= 16'h2ecb;
        src45 <= 16'h8619;
        src46 <= 16'h1ac6;
        src47 <= 16'hb024;
        src48 <= 16'h742d;
        src49 <= 16'he8d3;
        src50 <= 16'h69c;
        src51 <= 16'hc1af;
        src52 <= 16'h5be9;
        src53 <= 16'h2f9e;
        exp <= 22'h1debf7;
        #1
        src0 <= 16'h7512;
        src1 <= 16'h971f;
        src2 <= 16'hac1;
        src3 <= 16'hb45;
        src4 <= 16'h3e5a;
        src5 <= 16'hb40a;
        src6 <= 16'hcc3b;
        src7 <= 16'h7be6;
        src8 <= 16'h3ad1;
        src9 <= 16'hf6a8;
        src10 <= 16'he619;
        src11 <= 16'hfb82;
        src12 <= 16'h219e;
        src13 <= 16'he841;
        src14 <= 16'h589f;
        src15 <= 16'h982f;
        src16 <= 16'hab45;
        src17 <= 16'h153;
        src18 <= 16'h8aac;
        src19 <= 16'hcea;
        src20 <= 16'h24e6;
        src21 <= 16'hd81f;
        src22 <= 16'h96de;
        src23 <= 16'h39be;
        src24 <= 16'h8c05;
        src25 <= 16'h88e6;
        src26 <= 16'h181d;
        src27 <= 16'hdbb7;
        src28 <= 16'h7d9d;
        src29 <= 16'h6c01;
        src30 <= 16'he4bf;
        src31 <= 16'hcbc4;
        src32 <= 16'h68ff;
        src33 <= 16'hb69e;
        src34 <= 16'hdbe1;
        src35 <= 16'hb0e;
        src36 <= 16'h9048;
        src37 <= 16'habd7;
        src38 <= 16'hdc2e;
        src39 <= 16'he69b;
        src40 <= 16'ha289;
        src41 <= 16'h6877;
        src42 <= 16'h7370;
        src43 <= 16'h9528;
        src44 <= 16'h3e7c;
        src45 <= 16'h479e;
        src46 <= 16'h5f41;
        src47 <= 16'h27a5;
        src48 <= 16'hcd73;
        src49 <= 16'hd382;
        src50 <= 16'hf72a;
        src51 <= 16'h550a;
        src52 <= 16'h25c7;
        src53 <= 16'h38ea;
        exp <= 22'h1b9112;
        #1
        src0 <= 16'hf808;
        src1 <= 16'h2e18;
        src2 <= 16'h2974;
        src3 <= 16'hab53;
        src4 <= 16'hbf39;
        src5 <= 16'ha9c0;
        src6 <= 16'h350c;
        src7 <= 16'hfa29;
        src8 <= 16'h4efc;
        src9 <= 16'h1fb3;
        src10 <= 16'h76f3;
        src11 <= 16'h87c4;
        src12 <= 16'h4d0f;
        src13 <= 16'hb09d;
        src14 <= 16'h2b37;
        src15 <= 16'hae85;
        src16 <= 16'hc6e4;
        src17 <= 16'hcbb5;
        src18 <= 16'hf0b3;
        src19 <= 16'h6e19;
        src20 <= 16'hdbee;
        src21 <= 16'h1e5e;
        src22 <= 16'hc20b;
        src23 <= 16'h6e26;
        src24 <= 16'h2950;
        src25 <= 16'hf60d;
        src26 <= 16'h6636;
        src27 <= 16'h9f6;
        src28 <= 16'h9317;
        src29 <= 16'hd06b;
        src30 <= 16'h2ee5;
        src31 <= 16'h725f;
        src32 <= 16'habe4;
        src33 <= 16'h7f5a;
        src34 <= 16'h9a99;
        src35 <= 16'h344;
        src36 <= 16'ha5a5;
        src37 <= 16'h6357;
        src38 <= 16'h1a8d;
        src39 <= 16'h5134;
        src40 <= 16'h410e;
        src41 <= 16'h7b01;
        src42 <= 16'h9d80;
        src43 <= 16'h3e27;
        src44 <= 16'h924d;
        src45 <= 16'h4e23;
        src46 <= 16'h6084;
        src47 <= 16'h34b4;
        src48 <= 16'hc9bf;
        src49 <= 16'h58dc;
        src50 <= 16'h1b46;
        src51 <= 16'h2b15;
        src52 <= 16'hea3c;
        src53 <= 16'h5b88;
        exp <= 22'h198204;
        #1
        src0 <= 16'h8fc7;
        src1 <= 16'hd827;
        src2 <= 16'hbab7;
        src3 <= 16'h6edd;
        src4 <= 16'h9e70;
        src5 <= 16'he3a1;
        src6 <= 16'hbf20;
        src7 <= 16'he995;
        src8 <= 16'h698;
        src9 <= 16'hae6b;
        src10 <= 16'h4088;
        src11 <= 16'h2541;
        src12 <= 16'hdcec;
        src13 <= 16'h1cbb;
        src14 <= 16'h6d32;
        src15 <= 16'hfdf1;
        src16 <= 16'hde03;
        src17 <= 16'hfcae;
        src18 <= 16'hc2c6;
        src19 <= 16'ha516;
        src20 <= 16'hfcce;
        src21 <= 16'h6cb;
        src22 <= 16'hd06;
        src23 <= 16'h2f7d;
        src24 <= 16'h52f1;
        src25 <= 16'hf176;
        src26 <= 16'he7fa;
        src27 <= 16'h9121;
        src28 <= 16'ha880;
        src29 <= 16'hb954;
        src30 <= 16'hef05;
        src31 <= 16'h4d6b;
        src32 <= 16'h9006;
        src33 <= 16'h1fbf;
        src34 <= 16'h7c39;
        src35 <= 16'hf253;
        src36 <= 16'hee36;
        src37 <= 16'h8012;
        src38 <= 16'hc8b9;
        src39 <= 16'heb0f;
        src40 <= 16'hc95a;
        src41 <= 16'he0a1;
        src42 <= 16'h122a;
        src43 <= 16'h590e;
        src44 <= 16'h7543;
        src45 <= 16'hb615;
        src46 <= 16'h5ff;
        src47 <= 16'hb1f4;
        src48 <= 16'hbcfe;
        src49 <= 16'hb9b4;
        src50 <= 16'h2e59;
        src51 <= 16'hb693;
        src52 <= 16'h496;
        src53 <= 16'h5f11;
        exp <= 22'h1f1271;
        #1
        src0 <= 16'h72c1;
        src1 <= 16'h1b9f;
        src2 <= 16'hca63;
        src3 <= 16'h4636;
        src4 <= 16'hf163;
        src5 <= 16'ha88a;
        src6 <= 16'he0a;
        src7 <= 16'hbbbd;
        src8 <= 16'hc556;
        src9 <= 16'h5f51;
        src10 <= 16'h369b;
        src11 <= 16'hf72f;
        src12 <= 16'h1755;
        src13 <= 16'h79b7;
        src14 <= 16'h5de;
        src15 <= 16'hea8d;
        src16 <= 16'h5585;
        src17 <= 16'h6b8;
        src18 <= 16'h6d8;
        src19 <= 16'hc648;
        src20 <= 16'h784d;
        src21 <= 16'he9cd;
        src22 <= 16'hd6c5;
        src23 <= 16'h3d31;
        src24 <= 16'hf58b;
        src25 <= 16'hd4d5;
        src26 <= 16'h5358;
        src27 <= 16'h9e0;
        src28 <= 16'h2046;
        src29 <= 16'h81bf;
        src30 <= 16'h7573;
        src31 <= 16'hf81c;
        src32 <= 16'h5304;
        src33 <= 16'h57b1;
        src34 <= 16'hb4be;
        src35 <= 16'hac84;
        src36 <= 16'h7a8f;
        src37 <= 16'h9ee4;
        src38 <= 16'hd603;
        src39 <= 16'h1134;
        src40 <= 16'h6b4e;
        src41 <= 16'h4bb;
        src42 <= 16'h9b9e;
        src43 <= 16'hec6a;
        src44 <= 16'heafe;
        src45 <= 16'hd987;
        src46 <= 16'h3051;
        src47 <= 16'h5d7b;
        src48 <= 16'h50c0;
        src49 <= 16'hb2b4;
        src50 <= 16'h87d8;
        src51 <= 16'h5c79;
        src52 <= 16'h2131;
        src53 <= 16'he08f;
        exp <= 22'h1aedb6;
        #1
        src0 <= 16'h1b77;
        src1 <= 16'h5f2;
        src2 <= 16'h27d;
        src3 <= 16'hb1f2;
        src4 <= 16'h28b;
        src5 <= 16'hf8e6;
        src6 <= 16'h7395;
        src7 <= 16'h4725;
        src8 <= 16'h2d79;
        src9 <= 16'hb370;
        src10 <= 16'ha065;
        src11 <= 16'h2092;
        src12 <= 16'hd447;
        src13 <= 16'h1d3b;
        src14 <= 16'h6ccc;
        src15 <= 16'h5638;
        src16 <= 16'h7b8f;
        src17 <= 16'h77a8;
        src18 <= 16'h1884;
        src19 <= 16'h5f24;
        src20 <= 16'h84d1;
        src21 <= 16'hdd16;
        src22 <= 16'h10cf;
        src23 <= 16'h9515;
        src24 <= 16'h66de;
        src25 <= 16'he1de;
        src26 <= 16'hd32a;
        src27 <= 16'hf4de;
        src28 <= 16'h7b84;
        src29 <= 16'hf26c;
        src30 <= 16'hbbe;
        src31 <= 16'h19b9;
        src32 <= 16'h58fa;
        src33 <= 16'hc569;
        src34 <= 16'h6cef;
        src35 <= 16'h549c;
        src36 <= 16'h6c60;
        src37 <= 16'hc76e;
        src38 <= 16'h9012;
        src39 <= 16'h1cb4;
        src40 <= 16'h2588;
        src41 <= 16'h4891;
        src42 <= 16'h5030;
        src43 <= 16'h1a01;
        src44 <= 16'h8b62;
        src45 <= 16'h684f;
        src46 <= 16'hd69e;
        src47 <= 16'h54dd;
        src48 <= 16'h4dba;
        src49 <= 16'h7664;
        src50 <= 16'ha890;
        src51 <= 16'h271;
        src52 <= 16'h3836;
        src53 <= 16'hef7b;
        exp <= 22'h174806;
        #1
        src0 <= 16'hecde;
        src1 <= 16'hd58c;
        src2 <= 16'hed76;
        src3 <= 16'h3cc7;
        src4 <= 16'h8a6e;
        src5 <= 16'hc407;
        src6 <= 16'h5fe2;
        src7 <= 16'hd3fe;
        src8 <= 16'hd338;
        src9 <= 16'h2f55;
        src10 <= 16'he7ad;
        src11 <= 16'h76f2;
        src12 <= 16'h2c92;
        src13 <= 16'h6ce2;
        src14 <= 16'h9b9a;
        src15 <= 16'h17f5;
        src16 <= 16'hcae3;
        src17 <= 16'h2a38;
        src18 <= 16'h1445;
        src19 <= 16'h6034;
        src20 <= 16'hf023;
        src21 <= 16'hedb0;
        src22 <= 16'h7826;
        src23 <= 16'hc714;
        src24 <= 16'h9565;
        src25 <= 16'hca89;
        src26 <= 16'hef98;
        src27 <= 16'ha2b4;
        src28 <= 16'h5bd8;
        src29 <= 16'h2a6f;
        src30 <= 16'h1c12;
        src31 <= 16'h1c76;
        src32 <= 16'hde4e;
        src33 <= 16'h998f;
        src34 <= 16'h1164;
        src35 <= 16'hf683;
        src36 <= 16'h7015;
        src37 <= 16'he5a3;
        src38 <= 16'h66a2;
        src39 <= 16'hfda0;
        src40 <= 16'h2d8f;
        src41 <= 16'h1cb7;
        src42 <= 16'he7e8;
        src43 <= 16'h2a63;
        src44 <= 16'h3850;
        src45 <= 16'hf744;
        src46 <= 16'h75ee;
        src47 <= 16'h9635;
        src48 <= 16'hd3f3;
        src49 <= 16'h8776;
        src50 <= 16'hdf9e;
        src51 <= 16'h7415;
        src52 <= 16'h638c;
        src53 <= 16'h2fb8;
        exp <= 22'h1d693b;
        #1
        src0 <= 16'hda52;
        src1 <= 16'h52d3;
        src2 <= 16'h88f7;
        src3 <= 16'hbac7;
        src4 <= 16'h7051;
        src5 <= 16'hf392;
        src6 <= 16'h9b75;
        src7 <= 16'h3371;
        src8 <= 16'h7ebf;
        src9 <= 16'hc587;
        src10 <= 16'hf477;
        src11 <= 16'h11c7;
        src12 <= 16'h4c72;
        src13 <= 16'hc00;
        src14 <= 16'h1c71;
        src15 <= 16'hc99e;
        src16 <= 16'h318f;
        src17 <= 16'hf21e;
        src18 <= 16'hf461;
        src19 <= 16'had3c;
        src20 <= 16'h3129;
        src21 <= 16'h2bdd;
        src22 <= 16'ha82a;
        src23 <= 16'hf559;
        src24 <= 16'h3c0c;
        src25 <= 16'hc804;
        src26 <= 16'h70bb;
        src27 <= 16'hf4e9;
        src28 <= 16'h6403;
        src29 <= 16'hff66;
        src30 <= 16'h1223;
        src31 <= 16'haf8a;
        src32 <= 16'h2066;
        src33 <= 16'hb9ab;
        src34 <= 16'h3073;
        src35 <= 16'h3c9d;
        src36 <= 16'he765;
        src37 <= 16'h604;
        src38 <= 16'h6daa;
        src39 <= 16'ha31f;
        src40 <= 16'h7ca4;
        src41 <= 16'h2c5e;
        src42 <= 16'hfc76;
        src43 <= 16'h7cb9;
        src44 <= 16'h64bf;
        src45 <= 16'h1e80;
        src46 <= 16'h875b;
        src47 <= 16'h982e;
        src48 <= 16'h6c26;
        src49 <= 16'hb57e;
        src50 <= 16'hc1b1;
        src51 <= 16'h1dcf;
        src52 <= 16'he79e;
        src53 <= 16'h3f92;
        exp <= 22'h1badee;
        #1
        src0 <= 16'hd17c;
        src1 <= 16'h2e60;
        src2 <= 16'hf0bf;
        src3 <= 16'h94a6;
        src4 <= 16'h160f;
        src5 <= 16'hbc59;
        src6 <= 16'hb47e;
        src7 <= 16'h91b6;
        src8 <= 16'h9472;
        src9 <= 16'hd0a2;
        src10 <= 16'h9531;
        src11 <= 16'h8e7f;
        src12 <= 16'hdf98;
        src13 <= 16'hf506;
        src14 <= 16'hce8c;
        src15 <= 16'h2a7;
        src16 <= 16'h3a6f;
        src17 <= 16'hc01f;
        src18 <= 16'h906c;
        src19 <= 16'hdc8;
        src20 <= 16'hf6cc;
        src21 <= 16'h1813;
        src22 <= 16'h38ba;
        src23 <= 16'h376f;
        src24 <= 16'h27c1;
        src25 <= 16'h62a;
        src26 <= 16'h3f77;
        src27 <= 16'h76d9;
        src28 <= 16'h63f4;
        src29 <= 16'he1f8;
        src30 <= 16'hb27a;
        src31 <= 16'hd257;
        src32 <= 16'h25f8;
        src33 <= 16'h3708;
        src34 <= 16'hd76f;
        src35 <= 16'h5d91;
        src36 <= 16'h4e82;
        src37 <= 16'h8281;
        src38 <= 16'h943f;
        src39 <= 16'h7ace;
        src40 <= 16'h54a4;
        src41 <= 16'h75e8;
        src42 <= 16'h6bcd;
        src43 <= 16'he9ae;
        src44 <= 16'h7b15;
        src45 <= 16'h419a;
        src46 <= 16'hddba;
        src47 <= 16'h8d50;
        src48 <= 16'had11;
        src49 <= 16'ha45a;
        src50 <= 16'h8d27;
        src51 <= 16'h78d5;
        src52 <= 16'h7a1f;
        src53 <= 16'habbf;
        exp <= 22'h1bca49;
        #1
        $finish;
    end
endmodule

