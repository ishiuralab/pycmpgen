module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37);
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    reg [53:0] src16;
    reg [53:0] src17;
    reg [53:0] src18;
    reg [53:0] src19;
    reg [53:0] src20;
    reg [53:0] src21;
    reg [53:0] src22;
    reg [53:0] src23;
    reg [53:0] src24;
    reg [53:0] src25;
    reg [53:0] src26;
    reg [53:0] src27;
    reg [53:0] src28;
    reg [53:0] src29;
    reg [53:0] src30;
    reg [53:0] src31;
    compressor_CLA54_32 compressor_CLA54_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37));
    initial begin
        src0 <= 54'h0;
        src1 <= 54'h0;
        src2 <= 54'h0;
        src3 <= 54'h0;
        src4 <= 54'h0;
        src5 <= 54'h0;
        src6 <= 54'h0;
        src7 <= 54'h0;
        src8 <= 54'h0;
        src9 <= 54'h0;
        src10 <= 54'h0;
        src11 <= 54'h0;
        src12 <= 54'h0;
        src13 <= 54'h0;
        src14 <= 54'h0;
        src15 <= 54'h0;
        src16 <= 54'h0;
        src17 <= 54'h0;
        src18 <= 54'h0;
        src19 <= 54'h0;
        src20 <= 54'h0;
        src21 <= 54'h0;
        src22 <= 54'h0;
        src23 <= 54'h0;
        src24 <= 54'h0;
        src25 <= 54'h0;
        src26 <= 54'h0;
        src27 <= 54'h0;
        src28 <= 54'h0;
        src29 <= 54'h0;
        src30 <= 54'h0;
        src31 <= 54'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA54_32(
    input [53:0]src0,
    input [53:0]src1,
    input [53:0]src2,
    input [53:0]src3,
    input [53:0]src4,
    input [53:0]src5,
    input [53:0]src6,
    input [53:0]src7,
    input [53:0]src8,
    input [53:0]src9,
    input [53:0]src10,
    input [53:0]src11,
    input [53:0]src12,
    input [53:0]src13,
    input [53:0]src14,
    input [53:0]src15,
    input [53:0]src16,
    input [53:0]src17,
    input [53:0]src18,
    input [53:0]src19,
    input [53:0]src20,
    input [53:0]src21,
    input [53:0]src22,
    input [53:0]src23,
    input [53:0]src24,
    input [53:0]src25,
    input [53:0]src26,
    input [53:0]src27,
    input [53:0]src28,
    input [53:0]src29,
    input [53:0]src30,
    input [53:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [0:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [0:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [0:0] comp_out37;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], 1'h0, comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], 1'h0, comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      input wire [53:0] src12,
      input wire [53:0] src13,
      input wire [53:0] src14,
      input wire [53:0] src15,
      input wire [53:0] src16,
      input wire [53:0] src17,
      input wire [53:0] src18,
      input wire [53:0] src19,
      input wire [53:0] src20,
      input wire [53:0] src21,
      input wire [53:0] src22,
      input wire [53:0] src23,
      input wire [53:0] src24,
      input wire [53:0] src25,
      input wire [53:0] src26,
      input wire [53:0] src27,
      input wire [53:0] src28,
      input wire [53:0] src29,
      input wire [53:0] src30,
      input wire [53:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [0:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [0:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [0:0] dst37);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [53:0] stage0_12;
   wire [53:0] stage0_13;
   wire [53:0] stage0_14;
   wire [53:0] stage0_15;
   wire [53:0] stage0_16;
   wire [53:0] stage0_17;
   wire [53:0] stage0_18;
   wire [53:0] stage0_19;
   wire [53:0] stage0_20;
   wire [53:0] stage0_21;
   wire [53:0] stage0_22;
   wire [53:0] stage0_23;
   wire [53:0] stage0_24;
   wire [53:0] stage0_25;
   wire [53:0] stage0_26;
   wire [53:0] stage0_27;
   wire [53:0] stage0_28;
   wire [53:0] stage0_29;
   wire [53:0] stage0_30;
   wire [53:0] stage0_31;
   wire [15:0] stage1_0;
   wire [16:0] stage1_1;
   wire [21:0] stage1_2;
   wire [21:0] stage1_3;
   wire [32:0] stage1_4;
   wire [26:0] stage1_5;
   wire [32:0] stage1_6;
   wire [20:0] stage1_7;
   wire [25:0] stage1_8;
   wire [35:0] stage1_9;
   wire [17:0] stage1_10;
   wire [28:0] stage1_11;
   wire [23:0] stage1_12;
   wire [31:0] stage1_13;
   wire [30:0] stage1_14;
   wire [27:0] stage1_15;
   wire [24:0] stage1_16;
   wire [19:0] stage1_17;
   wire [29:0] stage1_18;
   wire [31:0] stage1_19;
   wire [22:0] stage1_20;
   wire [29:0] stage1_21;
   wire [21:0] stage1_22;
   wire [28:0] stage1_23;
   wire [23:0] stage1_24;
   wire [22:0] stage1_25;
   wire [17:0] stage1_26;
   wire [24:0] stage1_27;
   wire [25:0] stage1_28;
   wire [24:0] stage1_29;
   wire [17:0] stage1_30;
   wire [23:0] stage1_31;
   wire [16:0] stage1_32;
   wire [7:0] stage1_33;
   wire [9:0] stage2_0;
   wire [11:0] stage2_1;
   wire [16:0] stage2_2;
   wire [10:0] stage2_3;
   wire [9:0] stage2_4;
   wire [11:0] stage2_5;
   wire [11:0] stage2_6;
   wire [15:0] stage2_7;
   wire [16:0] stage2_8;
   wire [9:0] stage2_9;
   wire [8:0] stage2_10;
   wire [9:0] stage2_11;
   wire [15:0] stage2_12;
   wire [18:0] stage2_13;
   wire [9:0] stage2_14;
   wire [11:0] stage2_15;
   wire [10:0] stage2_16;
   wire [11:0] stage2_17;
   wire [13:0] stage2_18;
   wire [9:0] stage2_19;
   wire [10:0] stage2_20;
   wire [11:0] stage2_21;
   wire [16:0] stage2_22;
   wire [16:0] stage2_23;
   wire [17:0] stage2_24;
   wire [11:0] stage2_25;
   wire [8:0] stage2_26;
   wire [6:0] stage2_27;
   wire [13:0] stage2_28;
   wire [17:0] stage2_29;
   wire [10:0] stage2_30;
   wire [9:0] stage2_31;
   wire [6:0] stage2_32;
   wire [6:0] stage2_33;
   wire [3:0] stage2_34;
   wire [1:0] stage2_35;
   wire [1:0] stage3_0;
   wire [11:0] stage3_1;
   wire [2:0] stage3_2;
   wire [12:0] stage3_3;
   wire [4:0] stage3_4;
   wire [2:0] stage3_5;
   wire [4:0] stage3_6;
   wire [8:0] stage3_7;
   wire [8:0] stage3_8;
   wire [7:0] stage3_9;
   wire [6:0] stage3_10;
   wire [3:0] stage3_11;
   wire [5:0] stage3_12;
   wire [6:0] stage3_13;
   wire [5:0] stage3_14;
   wire [5:0] stage3_15;
   wire [8:0] stage3_16;
   wire [2:0] stage3_17;
   wire [6:0] stage3_18;
   wire [6:0] stage3_19;
   wire [7:0] stage3_20;
   wire [6:0] stage3_21;
   wire [7:0] stage3_22;
   wire [6:0] stage3_23;
   wire [4:0] stage3_24;
   wire [5:0] stage3_25;
   wire [9:0] stage3_26;
   wire [2:0] stage3_27;
   wire [3:0] stage3_28;
   wire [18:0] stage3_29;
   wire [2:0] stage3_30;
   wire [6:0] stage3_31;
   wire [3:0] stage3_32;
   wire [1:0] stage3_33;
   wire [4:0] stage3_34;
   wire [3:0] stage3_35;
   wire [1:0] stage4_0;
   wire [3:0] stage4_1;
   wire [2:0] stage4_2;
   wire [2:0] stage4_3;
   wire [2:0] stage4_4;
   wire [2:0] stage4_5;
   wire [2:0] stage4_6;
   wire [2:0] stage4_7;
   wire [4:0] stage4_8;
   wire [3:0] stage4_9;
   wire [4:0] stage4_10;
   wire [2:0] stage4_11;
   wire [1:0] stage4_12;
   wire [2:0] stage4_13;
   wire [2:0] stage4_14;
   wire [3:0] stage4_15;
   wire [5:0] stage4_16;
   wire [1:0] stage4_17;
   wire [3:0] stage4_18;
   wire [1:0] stage4_19;
   wire [2:0] stage4_20;
   wire [2:0] stage4_21;
   wire [5:0] stage4_22;
   wire [2:0] stage4_23;
   wire [1:0] stage4_24;
   wire [5:0] stage4_25;
   wire [7:0] stage4_26;
   wire [0:0] stage4_27;
   wire [1:0] stage4_28;
   wire [5:0] stage4_29;
   wire [4:0] stage4_30;
   wire [5:0] stage4_31;
   wire [3:0] stage4_32;
   wire [0:0] stage4_33;
   wire [0:0] stage4_34;
   wire [1:0] stage4_35;
   wire [1:0] stage4_36;
   wire [0:0] stage4_37;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [0:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [1:0] stage5_19;
   wire [1:0] stage5_20;
   wire [0:0] stage5_21;
   wire [1:0] stage5_22;
   wire [1:0] stage5_23;
   wire [1:0] stage5_24;
   wire [1:0] stage5_25;
   wire [1:0] stage5_26;
   wire [1:0] stage5_27;
   wire [1:0] stage5_28;
   wire [1:0] stage5_29;
   wire [1:0] stage5_30;
   wire [1:0] stage5_31;
   wire [1:0] stage5_32;
   wire [1:0] stage5_33;
   wire [1:0] stage5_34;
   wire [1:0] stage5_35;
   wire [1:0] stage5_36;
   wire [0:0] stage5_37;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;
   assign dst22 = stage5_22;
   assign dst23 = stage5_23;
   assign dst24 = stage5_24;
   assign dst25 = stage5_25;
   assign dst26 = stage5_26;
   assign dst27 = stage5_27;
   assign dst28 = stage5_28;
   assign dst29 = stage5_29;
   assign dst30 = stage5_30;
   assign dst31 = stage5_31;
   assign dst32 = stage5_32;
   assign dst33 = stage5_33;
   assign dst34 = stage5_34;
   assign dst35 = stage5_35;
   assign dst36 = stage5_36;
   assign dst37 = stage5_37;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30]},
      {stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36]},
      {stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc615_5 gpc7 (
      {stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_1[15]},
      {stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc615_5 gpc8 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46]},
      {stage0_1[16]},
      {stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_1[17], stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21]},
      {stage0_2[29], stage0_2[30], stage0_2[31]},
      {stage0_3[10]},
      {stage0_4[0], stage0_4[1]},
      {stage1_5[0],stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27]},
      {stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16]},
      {stage1_5[1],stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33]},
      {stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22]},
      {stage1_5[2],stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39]},
      {stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28]},
      {stage1_5[3],stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45]},
      {stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34]},
      {stage1_5[4],stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51]},
      {stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40]},
      {stage1_5[5],stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14]}
   );
   gpc606_5 gpc15 (
      {stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37]},
      {stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5], stage0_4[6], stage0_4[7]},
      {stage1_6[0],stage1_5[6],stage1_4[15],stage1_3[15],stage1_2[15]}
   );
   gpc606_5 gpc16 (
      {stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43]},
      {stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13]},
      {stage1_6[1],stage1_5[7],stage1_4[16],stage1_3[16],stage1_2[16]}
   );
   gpc606_5 gpc17 (
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49]},
      {stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage1_6[2],stage1_5[8],stage1_4[17],stage1_3[17],stage1_2[17]}
   );
   gpc606_5 gpc18 (
      {stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[3],stage1_5[9],stage1_4[18],stage1_3[18]}
   );
   gpc615_5 gpc19 (
      {stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage0_4[20]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[4],stage1_5[10],stage1_4[19],stage1_3[19]}
   );
   gpc606_5 gpc20 (
      {stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[2],stage1_6[5],stage1_5[11],stage1_4[20]}
   );
   gpc606_5 gpc21 (
      {stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[3],stage1_6[6],stage1_5[12],stage1_4[21]}
   );
   gpc606_5 gpc22 (
      {stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[4],stage1_6[7],stage1_5[13],stage1_4[22]}
   );
   gpc606_5 gpc23 (
      {stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[5],stage1_6[8],stage1_5[14],stage1_4[23]}
   );
   gpc606_5 gpc24 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[4],stage1_7[6],stage1_6[9],stage1_5[15]}
   );
   gpc606_5 gpc25 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[5],stage1_7[7],stage1_6[10],stage1_5[16]}
   );
   gpc606_5 gpc26 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[6],stage1_7[8],stage1_6[11],stage1_5[17]}
   );
   gpc606_5 gpc27 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[7],stage1_7[9],stage1_6[12],stage1_5[18]}
   );
   gpc606_5 gpc28 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[8],stage1_7[10],stage1_6[13],stage1_5[19]}
   );
   gpc606_5 gpc29 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[9],stage1_7[11],stage1_6[14],stage1_5[20]}
   );
   gpc615_5 gpc30 (
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28]},
      {stage0_7[36]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[6],stage1_8[10],stage1_7[12],stage1_6[15]}
   );
   gpc615_5 gpc31 (
      {stage0_6[29], stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33]},
      {stage0_7[37]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[7],stage1_8[11],stage1_7[13],stage1_6[16]}
   );
   gpc615_5 gpc32 (
      {stage0_6[34], stage0_6[35], stage0_6[36], stage0_6[37], stage0_6[38]},
      {stage0_7[38]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[8],stage1_8[12],stage1_7[14],stage1_6[17]}
   );
   gpc606_5 gpc33 (
      {stage0_7[39], stage0_7[40], stage0_7[41], stage0_7[42], stage0_7[43], stage0_7[44]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[9],stage1_8[13],stage1_7[15]}
   );
   gpc615_5 gpc34 (
      {stage0_7[45], stage0_7[46], stage0_7[47], stage0_7[48], stage0_7[49]},
      {stage0_8[18]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[4],stage1_9[10],stage1_8[14],stage1_7[16]}
   );
   gpc1163_5 gpc35 (
      {stage0_8[19], stage0_8[20], stage0_8[21]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage0_10[0]},
      {stage0_11[0]},
      {stage1_12[0],stage1_11[2],stage1_10[5],stage1_9[11],stage1_8[15]}
   );
   gpc606_5 gpc36 (
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6]},
      {stage1_12[1],stage1_11[3],stage1_10[6],stage1_9[12],stage1_8[16]}
   );
   gpc606_5 gpc37 (
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11], stage0_10[12]},
      {stage1_12[2],stage1_11[4],stage1_10[7],stage1_9[13],stage1_8[17]}
   );
   gpc615_5 gpc38 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38]},
      {stage0_9[18]},
      {stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17], stage0_10[18]},
      {stage1_12[3],stage1_11[5],stage1_10[8],stage1_9[14],stage1_8[18]}
   );
   gpc615_5 gpc39 (
      {stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_9[19]},
      {stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23], stage0_10[24]},
      {stage1_12[4],stage1_11[6],stage1_10[9],stage1_9[15],stage1_8[19]}
   );
   gpc615_5 gpc40 (
      {stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_9[20]},
      {stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29], stage0_10[30]},
      {stage1_12[5],stage1_11[7],stage1_10[10],stage1_9[16],stage1_8[20]}
   );
   gpc606_5 gpc41 (
      {stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6]},
      {stage1_13[0],stage1_12[6],stage1_11[8],stage1_10[11],stage1_9[17]}
   );
   gpc606_5 gpc42 (
      {stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32]},
      {stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12]},
      {stage1_13[1],stage1_12[7],stage1_11[9],stage1_10[12],stage1_9[18]}
   );
   gpc615_5 gpc43 (
      {stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_10[31]},
      {stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17], stage0_11[18]},
      {stage1_13[2],stage1_12[8],stage1_11[10],stage1_10[13],stage1_9[19]}
   );
   gpc606_5 gpc44 (
      {stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35], stage0_10[36], stage0_10[37]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[3],stage1_12[9],stage1_11[11],stage1_10[14]}
   );
   gpc606_5 gpc45 (
      {stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[4],stage1_12[10],stage1_11[12],stage1_10[15]}
   );
   gpc615_5 gpc46 (
      {stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47], stage0_10[48]},
      {stage0_11[19]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[5],stage1_12[11],stage1_11[13],stage1_10[16]}
   );
   gpc615_5 gpc47 (
      {stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage0_11[20]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[6],stage1_12[12],stage1_11[14],stage1_10[17]}
   );
   gpc606_5 gpc48 (
      {stage0_11[21], stage0_11[22], stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[4],stage1_13[7],stage1_12[13],stage1_11[15]}
   );
   gpc606_5 gpc49 (
      {stage0_11[27], stage0_11[28], stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[5],stage1_13[8],stage1_12[14],stage1_11[16]}
   );
   gpc606_5 gpc50 (
      {stage0_11[33], stage0_11[34], stage0_11[35], stage0_11[36], stage0_11[37], stage0_11[38]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[6],stage1_13[9],stage1_12[15],stage1_11[17]}
   );
   gpc615_5 gpc51 (
      {stage0_11[39], stage0_11[40], stage0_11[41], stage0_11[42], stage0_11[43]},
      {stage0_12[24]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[7],stage1_13[10],stage1_12[16],stage1_11[18]}
   );
   gpc1423_5 gpc52 (
      {stage0_12[25], stage0_12[26], stage0_12[27]},
      {stage0_13[24], stage0_13[25]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3]},
      {stage0_15[0]},
      {stage1_16[0],stage1_15[4],stage1_14[8],stage1_13[11],stage1_12[17]}
   );
   gpc606_5 gpc53 (
      {stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33]},
      {stage0_14[4], stage0_14[5], stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9]},
      {stage1_16[1],stage1_15[5],stage1_14[9],stage1_13[12],stage1_12[18]}
   );
   gpc606_5 gpc54 (
      {stage0_12[34], stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39]},
      {stage0_14[10], stage0_14[11], stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15]},
      {stage1_16[2],stage1_15[6],stage1_14[10],stage1_13[13],stage1_12[19]}
   );
   gpc606_5 gpc55 (
      {stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45]},
      {stage0_14[16], stage0_14[17], stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21]},
      {stage1_16[3],stage1_15[7],stage1_14[11],stage1_13[14],stage1_12[20]}
   );
   gpc606_5 gpc56 (
      {stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51]},
      {stage0_14[22], stage0_14[23], stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27]},
      {stage1_16[4],stage1_15[8],stage1_14[12],stage1_13[15],stage1_12[21]}
   );
   gpc615_5 gpc57 (
      {stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29], stage0_13[30]},
      {stage0_14[28]},
      {stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5], stage0_15[6]},
      {stage1_17[0],stage1_16[5],stage1_15[9],stage1_14[13],stage1_13[16]}
   );
   gpc615_5 gpc58 (
      {stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_14[29]},
      {stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11], stage0_15[12]},
      {stage1_17[1],stage1_16[6],stage1_15[10],stage1_14[14],stage1_13[17]}
   );
   gpc615_5 gpc59 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40]},
      {stage0_14[30]},
      {stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17], stage0_15[18]},
      {stage1_17[2],stage1_16[7],stage1_15[11],stage1_14[15],stage1_13[18]}
   );
   gpc615_5 gpc60 (
      {stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage0_15[19]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[3],stage1_16[8],stage1_15[12],stage1_14[16]}
   );
   gpc615_5 gpc61 (
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40]},
      {stage0_15[20]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[4],stage1_16[9],stage1_15[13],stage1_14[17]}
   );
   gpc606_5 gpc62 (
      {stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24], stage0_15[25], stage0_15[26]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[2],stage1_17[5],stage1_16[10],stage1_15[14]}
   );
   gpc606_5 gpc63 (
      {stage0_15[27], stage0_15[28], stage0_15[29], stage0_15[30], stage0_15[31], stage0_15[32]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[3],stage1_17[6],stage1_16[11],stage1_15[15]}
   );
   gpc606_5 gpc64 (
      {stage0_15[33], stage0_15[34], stage0_15[35], stage0_15[36], stage0_15[37], stage0_15[38]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[4],stage1_17[7],stage1_16[12],stage1_15[16]}
   );
   gpc615_5 gpc65 (
      {stage0_15[39], stage0_15[40], stage0_15[41], stage0_15[42], stage0_15[43]},
      {stage0_16[12]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[5],stage1_17[8],stage1_16[13],stage1_15[17]}
   );
   gpc606_5 gpc66 (
      {stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17], stage0_16[18]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[4],stage1_18[6],stage1_17[9],stage1_16[14]}
   );
   gpc606_5 gpc67 (
      {stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23], stage0_16[24]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[5],stage1_18[7],stage1_17[10],stage1_16[15]}
   );
   gpc606_5 gpc68 (
      {stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[6],stage1_18[8],stage1_17[11],stage1_16[16]}
   );
   gpc606_5 gpc69 (
      {stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35], stage0_16[36]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[7],stage1_18[9],stage1_17[12],stage1_16[17]}
   );
   gpc606_5 gpc70 (
      {stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[8],stage1_18[10],stage1_17[13],stage1_16[18]}
   );
   gpc606_5 gpc71 (
      {stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47], stage0_16[48]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[9],stage1_18[11],stage1_17[14],stage1_16[19]}
   );
   gpc606_5 gpc72 (
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[6],stage1_19[10],stage1_18[12],stage1_17[15]}
   );
   gpc606_5 gpc73 (
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[7],stage1_19[11],stage1_18[13],stage1_17[16]}
   );
   gpc606_5 gpc74 (
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[8],stage1_19[12],stage1_18[14],stage1_17[17]}
   );
   gpc606_5 gpc75 (
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[9],stage1_19[13],stage1_18[15],stage1_17[18]}
   );
   gpc606_5 gpc76 (
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[10],stage1_19[14],stage1_18[16],stage1_17[19]}
   );
   gpc606_5 gpc77 (
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[5],stage1_20[11],stage1_19[15],stage1_18[17]}
   );
   gpc615_5 gpc78 (
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34]},
      {stage0_20[6]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[1],stage1_21[6],stage1_20[12],stage1_19[16]}
   );
   gpc615_5 gpc79 (
      {stage0_19[35], stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39]},
      {stage0_20[7]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[2],stage1_21[7],stage1_20[13],stage1_19[17]}
   );
   gpc606_5 gpc80 (
      {stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11], stage0_20[12], stage0_20[13]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[2],stage1_22[3],stage1_21[8],stage1_20[14]}
   );
   gpc606_5 gpc81 (
      {stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17], stage0_20[18], stage0_20[19]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[3],stage1_22[4],stage1_21[9],stage1_20[15]}
   );
   gpc606_5 gpc82 (
      {stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23], stage0_20[24], stage0_20[25]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[4],stage1_22[5],stage1_21[10],stage1_20[16]}
   );
   gpc606_5 gpc83 (
      {stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[5],stage1_22[6],stage1_21[11],stage1_20[17]}
   );
   gpc606_5 gpc84 (
      {stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[6],stage1_22[7],stage1_21[12],stage1_20[18]}
   );
   gpc615_5 gpc85 (
      {stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42]},
      {stage0_21[12]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[7],stage1_22[8],stage1_21[13],stage1_20[19]}
   );
   gpc615_5 gpc86 (
      {stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage0_21[13]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[8],stage1_22[9],stage1_21[14],stage1_20[20]}
   );
   gpc615_5 gpc87 (
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[14]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[9],stage1_22[10],stage1_21[15],stage1_20[21]}
   );
   gpc606_5 gpc88 (
      {stage0_21[15], stage0_21[16], stage0_21[17], stage0_21[18], stage0_21[19], stage0_21[20]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[8],stage1_23[10],stage1_22[11],stage1_21[16]}
   );
   gpc606_5 gpc89 (
      {stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25], stage0_21[26]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[9],stage1_23[11],stage1_22[12],stage1_21[17]}
   );
   gpc606_5 gpc90 (
      {stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30], stage0_21[31], stage0_21[32]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[10],stage1_23[12],stage1_22[13],stage1_21[18]}
   );
   gpc606_5 gpc91 (
      {stage0_21[33], stage0_21[34], stage0_21[35], stage0_21[36], stage0_21[37], stage0_21[38]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[11],stage1_23[13],stage1_22[14],stage1_21[19]}
   );
   gpc606_5 gpc92 (
      {stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42], stage0_21[43], stage0_21[44]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[12],stage1_23[14],stage1_22[15],stage1_21[20]}
   );
   gpc606_5 gpc93 (
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[0],stage1_25[5],stage1_24[13],stage1_23[15]}
   );
   gpc606_5 gpc94 (
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[1],stage1_25[6],stage1_24[14],stage1_23[16]}
   );
   gpc606_5 gpc95 (
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[2],stage1_26[2],stage1_25[7],stage1_24[15]}
   );
   gpc606_5 gpc96 (
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[3],stage1_26[3],stage1_25[8],stage1_24[16]}
   );
   gpc606_5 gpc97 (
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[4],stage1_26[4],stage1_25[9],stage1_24[17]}
   );
   gpc606_5 gpc98 (
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[5],stage1_26[5],stage1_25[10],stage1_24[18]}
   );
   gpc606_5 gpc99 (
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[6],stage1_26[6],stage1_25[11],stage1_24[19]}
   );
   gpc606_5 gpc100 (
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[7],stage1_26[7],stage1_25[12],stage1_24[20]}
   );
   gpc606_5 gpc101 (
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[8],stage1_26[8],stage1_25[13],stage1_24[21]}
   );
   gpc606_5 gpc102 (
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[9],stage1_26[9],stage1_25[14],stage1_24[22]}
   );
   gpc606_5 gpc103 (
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[10],stage1_26[10],stage1_25[15],stage1_24[23]}
   );
   gpc606_5 gpc104 (
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[9],stage1_27[11],stage1_26[11],stage1_25[16]}
   );
   gpc606_5 gpc105 (
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[10],stage1_27[12],stage1_26[12],stage1_25[17]}
   );
   gpc606_5 gpc106 (
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[11],stage1_27[13],stage1_26[13],stage1_25[18]}
   );
   gpc606_5 gpc107 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[12],stage1_27[14],stage1_26[14],stage1_25[19]}
   );
   gpc606_5 gpc108 (
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[13],stage1_27[15],stage1_26[15],stage1_25[20]}
   );
   gpc606_5 gpc109 (
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[14],stage1_27[16],stage1_26[16],stage1_25[21]}
   );
   gpc606_5 gpc110 (
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[15],stage1_27[17],stage1_26[17],stage1_25[22]}
   );
   gpc606_5 gpc111 (
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[0],stage1_29[7],stage1_28[16],stage1_27[18]}
   );
   gpc606_5 gpc112 (
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[1],stage1_30[1],stage1_29[8],stage1_28[17]}
   );
   gpc606_5 gpc113 (
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[2],stage1_30[2],stage1_29[9],stage1_28[18]}
   );
   gpc606_5 gpc114 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[3],stage1_30[3],stage1_29[10],stage1_28[19]}
   );
   gpc606_5 gpc115 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[4],stage1_30[4],stage1_29[11],stage1_28[20]}
   );
   gpc606_5 gpc116 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[5],stage1_30[5],stage1_29[12],stage1_28[21]}
   );
   gpc606_5 gpc117 (
      {stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[6],stage1_30[6],stage1_29[13],stage1_28[22]}
   );
   gpc606_5 gpc118 (
      {stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[7],stage1_30[7],stage1_29[14],stage1_28[23]}
   );
   gpc606_5 gpc119 (
      {stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[8],stage1_30[8],stage1_29[15],stage1_28[24]}
   );
   gpc606_5 gpc120 (
      {stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[9],stage1_30[9],stage1_29[16],stage1_28[25]}
   );
   gpc606_5 gpc121 (
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[9],stage1_31[10],stage1_30[10],stage1_29[17]}
   );
   gpc606_5 gpc122 (
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[10],stage1_31[11],stage1_30[11],stage1_29[18]}
   );
   gpc606_5 gpc123 (
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[11],stage1_31[12],stage1_30[12],stage1_29[19]}
   );
   gpc606_5 gpc124 (
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[12],stage1_31[13],stage1_30[13],stage1_29[20]}
   );
   gpc606_5 gpc125 (
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[13],stage1_31[14],stage1_30[14],stage1_29[21]}
   );
   gpc606_5 gpc126 (
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[14],stage1_31[15],stage1_30[15],stage1_29[22]}
   );
   gpc606_5 gpc127 (
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[15],stage1_31[16],stage1_30[16],stage1_29[23]}
   );
   gpc606_5 gpc128 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[16],stage1_31[17],stage1_30[17],stage1_29[24]}
   );
   gpc1_1 gpc129 (
      {stage0_0[47]},
      {stage1_0[9]}
   );
   gpc1_1 gpc130 (
      {stage0_0[48]},
      {stage1_0[10]}
   );
   gpc1_1 gpc131 (
      {stage0_0[49]},
      {stage1_0[11]}
   );
   gpc1_1 gpc132 (
      {stage0_0[50]},
      {stage1_0[12]}
   );
   gpc1_1 gpc133 (
      {stage0_0[51]},
      {stage1_0[13]}
   );
   gpc1_1 gpc134 (
      {stage0_0[52]},
      {stage1_0[14]}
   );
   gpc1_1 gpc135 (
      {stage0_0[53]},
      {stage1_0[15]}
   );
   gpc1_1 gpc136 (
      {stage0_1[52]},
      {stage1_1[15]}
   );
   gpc1_1 gpc137 (
      {stage0_1[53]},
      {stage1_1[16]}
   );
   gpc1_1 gpc138 (
      {stage0_2[50]},
      {stage1_2[18]}
   );
   gpc1_1 gpc139 (
      {stage0_2[51]},
      {stage1_2[19]}
   );
   gpc1_1 gpc140 (
      {stage0_2[52]},
      {stage1_2[20]}
   );
   gpc1_1 gpc141 (
      {stage0_2[53]},
      {stage1_2[21]}
   );
   gpc1_1 gpc142 (
      {stage0_3[52]},
      {stage1_3[20]}
   );
   gpc1_1 gpc143 (
      {stage0_3[53]},
      {stage1_3[21]}
   );
   gpc1_1 gpc144 (
      {stage0_4[45]},
      {stage1_4[24]}
   );
   gpc1_1 gpc145 (
      {stage0_4[46]},
      {stage1_4[25]}
   );
   gpc1_1 gpc146 (
      {stage0_4[47]},
      {stage1_4[26]}
   );
   gpc1_1 gpc147 (
      {stage0_4[48]},
      {stage1_4[27]}
   );
   gpc1_1 gpc148 (
      {stage0_4[49]},
      {stage1_4[28]}
   );
   gpc1_1 gpc149 (
      {stage0_4[50]},
      {stage1_4[29]}
   );
   gpc1_1 gpc150 (
      {stage0_4[51]},
      {stage1_4[30]}
   );
   gpc1_1 gpc151 (
      {stage0_4[52]},
      {stage1_4[31]}
   );
   gpc1_1 gpc152 (
      {stage0_4[53]},
      {stage1_4[32]}
   );
   gpc1_1 gpc153 (
      {stage0_5[48]},
      {stage1_5[21]}
   );
   gpc1_1 gpc154 (
      {stage0_5[49]},
      {stage1_5[22]}
   );
   gpc1_1 gpc155 (
      {stage0_5[50]},
      {stage1_5[23]}
   );
   gpc1_1 gpc156 (
      {stage0_5[51]},
      {stage1_5[24]}
   );
   gpc1_1 gpc157 (
      {stage0_5[52]},
      {stage1_5[25]}
   );
   gpc1_1 gpc158 (
      {stage0_5[53]},
      {stage1_5[26]}
   );
   gpc1_1 gpc159 (
      {stage0_6[39]},
      {stage1_6[18]}
   );
   gpc1_1 gpc160 (
      {stage0_6[40]},
      {stage1_6[19]}
   );
   gpc1_1 gpc161 (
      {stage0_6[41]},
      {stage1_6[20]}
   );
   gpc1_1 gpc162 (
      {stage0_6[42]},
      {stage1_6[21]}
   );
   gpc1_1 gpc163 (
      {stage0_6[43]},
      {stage1_6[22]}
   );
   gpc1_1 gpc164 (
      {stage0_6[44]},
      {stage1_6[23]}
   );
   gpc1_1 gpc165 (
      {stage0_6[45]},
      {stage1_6[24]}
   );
   gpc1_1 gpc166 (
      {stage0_6[46]},
      {stage1_6[25]}
   );
   gpc1_1 gpc167 (
      {stage0_6[47]},
      {stage1_6[26]}
   );
   gpc1_1 gpc168 (
      {stage0_6[48]},
      {stage1_6[27]}
   );
   gpc1_1 gpc169 (
      {stage0_6[49]},
      {stage1_6[28]}
   );
   gpc1_1 gpc170 (
      {stage0_6[50]},
      {stage1_6[29]}
   );
   gpc1_1 gpc171 (
      {stage0_6[51]},
      {stage1_6[30]}
   );
   gpc1_1 gpc172 (
      {stage0_6[52]},
      {stage1_6[31]}
   );
   gpc1_1 gpc173 (
      {stage0_6[53]},
      {stage1_6[32]}
   );
   gpc1_1 gpc174 (
      {stage0_7[50]},
      {stage1_7[17]}
   );
   gpc1_1 gpc175 (
      {stage0_7[51]},
      {stage1_7[18]}
   );
   gpc1_1 gpc176 (
      {stage0_7[52]},
      {stage1_7[19]}
   );
   gpc1_1 gpc177 (
      {stage0_7[53]},
      {stage1_7[20]}
   );
   gpc1_1 gpc178 (
      {stage0_8[49]},
      {stage1_8[21]}
   );
   gpc1_1 gpc179 (
      {stage0_8[50]},
      {stage1_8[22]}
   );
   gpc1_1 gpc180 (
      {stage0_8[51]},
      {stage1_8[23]}
   );
   gpc1_1 gpc181 (
      {stage0_8[52]},
      {stage1_8[24]}
   );
   gpc1_1 gpc182 (
      {stage0_8[53]},
      {stage1_8[25]}
   );
   gpc1_1 gpc183 (
      {stage0_9[38]},
      {stage1_9[20]}
   );
   gpc1_1 gpc184 (
      {stage0_9[39]},
      {stage1_9[21]}
   );
   gpc1_1 gpc185 (
      {stage0_9[40]},
      {stage1_9[22]}
   );
   gpc1_1 gpc186 (
      {stage0_9[41]},
      {stage1_9[23]}
   );
   gpc1_1 gpc187 (
      {stage0_9[42]},
      {stage1_9[24]}
   );
   gpc1_1 gpc188 (
      {stage0_9[43]},
      {stage1_9[25]}
   );
   gpc1_1 gpc189 (
      {stage0_9[44]},
      {stage1_9[26]}
   );
   gpc1_1 gpc190 (
      {stage0_9[45]},
      {stage1_9[27]}
   );
   gpc1_1 gpc191 (
      {stage0_9[46]},
      {stage1_9[28]}
   );
   gpc1_1 gpc192 (
      {stage0_9[47]},
      {stage1_9[29]}
   );
   gpc1_1 gpc193 (
      {stage0_9[48]},
      {stage1_9[30]}
   );
   gpc1_1 gpc194 (
      {stage0_9[49]},
      {stage1_9[31]}
   );
   gpc1_1 gpc195 (
      {stage0_9[50]},
      {stage1_9[32]}
   );
   gpc1_1 gpc196 (
      {stage0_9[51]},
      {stage1_9[33]}
   );
   gpc1_1 gpc197 (
      {stage0_9[52]},
      {stage1_9[34]}
   );
   gpc1_1 gpc198 (
      {stage0_9[53]},
      {stage1_9[35]}
   );
   gpc1_1 gpc199 (
      {stage0_11[44]},
      {stage1_11[19]}
   );
   gpc1_1 gpc200 (
      {stage0_11[45]},
      {stage1_11[20]}
   );
   gpc1_1 gpc201 (
      {stage0_11[46]},
      {stage1_11[21]}
   );
   gpc1_1 gpc202 (
      {stage0_11[47]},
      {stage1_11[22]}
   );
   gpc1_1 gpc203 (
      {stage0_11[48]},
      {stage1_11[23]}
   );
   gpc1_1 gpc204 (
      {stage0_11[49]},
      {stage1_11[24]}
   );
   gpc1_1 gpc205 (
      {stage0_11[50]},
      {stage1_11[25]}
   );
   gpc1_1 gpc206 (
      {stage0_11[51]},
      {stage1_11[26]}
   );
   gpc1_1 gpc207 (
      {stage0_11[52]},
      {stage1_11[27]}
   );
   gpc1_1 gpc208 (
      {stage0_11[53]},
      {stage1_11[28]}
   );
   gpc1_1 gpc209 (
      {stage0_12[52]},
      {stage1_12[22]}
   );
   gpc1_1 gpc210 (
      {stage0_12[53]},
      {stage1_12[23]}
   );
   gpc1_1 gpc211 (
      {stage0_13[41]},
      {stage1_13[19]}
   );
   gpc1_1 gpc212 (
      {stage0_13[42]},
      {stage1_13[20]}
   );
   gpc1_1 gpc213 (
      {stage0_13[43]},
      {stage1_13[21]}
   );
   gpc1_1 gpc214 (
      {stage0_13[44]},
      {stage1_13[22]}
   );
   gpc1_1 gpc215 (
      {stage0_13[45]},
      {stage1_13[23]}
   );
   gpc1_1 gpc216 (
      {stage0_13[46]},
      {stage1_13[24]}
   );
   gpc1_1 gpc217 (
      {stage0_13[47]},
      {stage1_13[25]}
   );
   gpc1_1 gpc218 (
      {stage0_13[48]},
      {stage1_13[26]}
   );
   gpc1_1 gpc219 (
      {stage0_13[49]},
      {stage1_13[27]}
   );
   gpc1_1 gpc220 (
      {stage0_13[50]},
      {stage1_13[28]}
   );
   gpc1_1 gpc221 (
      {stage0_13[51]},
      {stage1_13[29]}
   );
   gpc1_1 gpc222 (
      {stage0_13[52]},
      {stage1_13[30]}
   );
   gpc1_1 gpc223 (
      {stage0_13[53]},
      {stage1_13[31]}
   );
   gpc1_1 gpc224 (
      {stage0_14[41]},
      {stage1_14[18]}
   );
   gpc1_1 gpc225 (
      {stage0_14[42]},
      {stage1_14[19]}
   );
   gpc1_1 gpc226 (
      {stage0_14[43]},
      {stage1_14[20]}
   );
   gpc1_1 gpc227 (
      {stage0_14[44]},
      {stage1_14[21]}
   );
   gpc1_1 gpc228 (
      {stage0_14[45]},
      {stage1_14[22]}
   );
   gpc1_1 gpc229 (
      {stage0_14[46]},
      {stage1_14[23]}
   );
   gpc1_1 gpc230 (
      {stage0_14[47]},
      {stage1_14[24]}
   );
   gpc1_1 gpc231 (
      {stage0_14[48]},
      {stage1_14[25]}
   );
   gpc1_1 gpc232 (
      {stage0_14[49]},
      {stage1_14[26]}
   );
   gpc1_1 gpc233 (
      {stage0_14[50]},
      {stage1_14[27]}
   );
   gpc1_1 gpc234 (
      {stage0_14[51]},
      {stage1_14[28]}
   );
   gpc1_1 gpc235 (
      {stage0_14[52]},
      {stage1_14[29]}
   );
   gpc1_1 gpc236 (
      {stage0_14[53]},
      {stage1_14[30]}
   );
   gpc1_1 gpc237 (
      {stage0_15[44]},
      {stage1_15[18]}
   );
   gpc1_1 gpc238 (
      {stage0_15[45]},
      {stage1_15[19]}
   );
   gpc1_1 gpc239 (
      {stage0_15[46]},
      {stage1_15[20]}
   );
   gpc1_1 gpc240 (
      {stage0_15[47]},
      {stage1_15[21]}
   );
   gpc1_1 gpc241 (
      {stage0_15[48]},
      {stage1_15[22]}
   );
   gpc1_1 gpc242 (
      {stage0_15[49]},
      {stage1_15[23]}
   );
   gpc1_1 gpc243 (
      {stage0_15[50]},
      {stage1_15[24]}
   );
   gpc1_1 gpc244 (
      {stage0_15[51]},
      {stage1_15[25]}
   );
   gpc1_1 gpc245 (
      {stage0_15[52]},
      {stage1_15[26]}
   );
   gpc1_1 gpc246 (
      {stage0_15[53]},
      {stage1_15[27]}
   );
   gpc1_1 gpc247 (
      {stage0_16[49]},
      {stage1_16[20]}
   );
   gpc1_1 gpc248 (
      {stage0_16[50]},
      {stage1_16[21]}
   );
   gpc1_1 gpc249 (
      {stage0_16[51]},
      {stage1_16[22]}
   );
   gpc1_1 gpc250 (
      {stage0_16[52]},
      {stage1_16[23]}
   );
   gpc1_1 gpc251 (
      {stage0_16[53]},
      {stage1_16[24]}
   );
   gpc1_1 gpc252 (
      {stage0_18[42]},
      {stage1_18[18]}
   );
   gpc1_1 gpc253 (
      {stage0_18[43]},
      {stage1_18[19]}
   );
   gpc1_1 gpc254 (
      {stage0_18[44]},
      {stage1_18[20]}
   );
   gpc1_1 gpc255 (
      {stage0_18[45]},
      {stage1_18[21]}
   );
   gpc1_1 gpc256 (
      {stage0_18[46]},
      {stage1_18[22]}
   );
   gpc1_1 gpc257 (
      {stage0_18[47]},
      {stage1_18[23]}
   );
   gpc1_1 gpc258 (
      {stage0_18[48]},
      {stage1_18[24]}
   );
   gpc1_1 gpc259 (
      {stage0_18[49]},
      {stage1_18[25]}
   );
   gpc1_1 gpc260 (
      {stage0_18[50]},
      {stage1_18[26]}
   );
   gpc1_1 gpc261 (
      {stage0_18[51]},
      {stage1_18[27]}
   );
   gpc1_1 gpc262 (
      {stage0_18[52]},
      {stage1_18[28]}
   );
   gpc1_1 gpc263 (
      {stage0_18[53]},
      {stage1_18[29]}
   );
   gpc1_1 gpc264 (
      {stage0_19[40]},
      {stage1_19[18]}
   );
   gpc1_1 gpc265 (
      {stage0_19[41]},
      {stage1_19[19]}
   );
   gpc1_1 gpc266 (
      {stage0_19[42]},
      {stage1_19[20]}
   );
   gpc1_1 gpc267 (
      {stage0_19[43]},
      {stage1_19[21]}
   );
   gpc1_1 gpc268 (
      {stage0_19[44]},
      {stage1_19[22]}
   );
   gpc1_1 gpc269 (
      {stage0_19[45]},
      {stage1_19[23]}
   );
   gpc1_1 gpc270 (
      {stage0_19[46]},
      {stage1_19[24]}
   );
   gpc1_1 gpc271 (
      {stage0_19[47]},
      {stage1_19[25]}
   );
   gpc1_1 gpc272 (
      {stage0_19[48]},
      {stage1_19[26]}
   );
   gpc1_1 gpc273 (
      {stage0_19[49]},
      {stage1_19[27]}
   );
   gpc1_1 gpc274 (
      {stage0_19[50]},
      {stage1_19[28]}
   );
   gpc1_1 gpc275 (
      {stage0_19[51]},
      {stage1_19[29]}
   );
   gpc1_1 gpc276 (
      {stage0_19[52]},
      {stage1_19[30]}
   );
   gpc1_1 gpc277 (
      {stage0_19[53]},
      {stage1_19[31]}
   );
   gpc1_1 gpc278 (
      {stage0_20[53]},
      {stage1_20[22]}
   );
   gpc1_1 gpc279 (
      {stage0_21[45]},
      {stage1_21[21]}
   );
   gpc1_1 gpc280 (
      {stage0_21[46]},
      {stage1_21[22]}
   );
   gpc1_1 gpc281 (
      {stage0_21[47]},
      {stage1_21[23]}
   );
   gpc1_1 gpc282 (
      {stage0_21[48]},
      {stage1_21[24]}
   );
   gpc1_1 gpc283 (
      {stage0_21[49]},
      {stage1_21[25]}
   );
   gpc1_1 gpc284 (
      {stage0_21[50]},
      {stage1_21[26]}
   );
   gpc1_1 gpc285 (
      {stage0_21[51]},
      {stage1_21[27]}
   );
   gpc1_1 gpc286 (
      {stage0_21[52]},
      {stage1_21[28]}
   );
   gpc1_1 gpc287 (
      {stage0_21[53]},
      {stage1_21[29]}
   );
   gpc1_1 gpc288 (
      {stage0_22[48]},
      {stage1_22[16]}
   );
   gpc1_1 gpc289 (
      {stage0_22[49]},
      {stage1_22[17]}
   );
   gpc1_1 gpc290 (
      {stage0_22[50]},
      {stage1_22[18]}
   );
   gpc1_1 gpc291 (
      {stage0_22[51]},
      {stage1_22[19]}
   );
   gpc1_1 gpc292 (
      {stage0_22[52]},
      {stage1_22[20]}
   );
   gpc1_1 gpc293 (
      {stage0_22[53]},
      {stage1_22[21]}
   );
   gpc1_1 gpc294 (
      {stage0_23[42]},
      {stage1_23[17]}
   );
   gpc1_1 gpc295 (
      {stage0_23[43]},
      {stage1_23[18]}
   );
   gpc1_1 gpc296 (
      {stage0_23[44]},
      {stage1_23[19]}
   );
   gpc1_1 gpc297 (
      {stage0_23[45]},
      {stage1_23[20]}
   );
   gpc1_1 gpc298 (
      {stage0_23[46]},
      {stage1_23[21]}
   );
   gpc1_1 gpc299 (
      {stage0_23[47]},
      {stage1_23[22]}
   );
   gpc1_1 gpc300 (
      {stage0_23[48]},
      {stage1_23[23]}
   );
   gpc1_1 gpc301 (
      {stage0_23[49]},
      {stage1_23[24]}
   );
   gpc1_1 gpc302 (
      {stage0_23[50]},
      {stage1_23[25]}
   );
   gpc1_1 gpc303 (
      {stage0_23[51]},
      {stage1_23[26]}
   );
   gpc1_1 gpc304 (
      {stage0_23[52]},
      {stage1_23[27]}
   );
   gpc1_1 gpc305 (
      {stage0_23[53]},
      {stage1_23[28]}
   );
   gpc1_1 gpc306 (
      {stage0_27[48]},
      {stage1_27[19]}
   );
   gpc1_1 gpc307 (
      {stage0_27[49]},
      {stage1_27[20]}
   );
   gpc1_1 gpc308 (
      {stage0_27[50]},
      {stage1_27[21]}
   );
   gpc1_1 gpc309 (
      {stage0_27[51]},
      {stage1_27[22]}
   );
   gpc1_1 gpc310 (
      {stage0_27[52]},
      {stage1_27[23]}
   );
   gpc1_1 gpc311 (
      {stage0_27[53]},
      {stage1_27[24]}
   );
   gpc1_1 gpc312 (
      {stage0_31[48]},
      {stage1_31[18]}
   );
   gpc1_1 gpc313 (
      {stage0_31[49]},
      {stage1_31[19]}
   );
   gpc1_1 gpc314 (
      {stage0_31[50]},
      {stage1_31[20]}
   );
   gpc1_1 gpc315 (
      {stage0_31[51]},
      {stage1_31[21]}
   );
   gpc1_1 gpc316 (
      {stage0_31[52]},
      {stage1_31[22]}
   );
   gpc1_1 gpc317 (
      {stage0_31[53]},
      {stage1_31[23]}
   );
   gpc1163_5 gpc318 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc615_5 gpc319 (
      {stage1_0[3], stage1_0[4], stage1_0[5], stage1_0[6], stage1_0[7]},
      {stage1_1[6]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc320 (
      {stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage1_4[0]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[2],stage2_3[2]}
   );
   gpc615_5 gpc321 (
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10]},
      {stage1_4[1]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[3],stage2_3[3]}
   );
   gpc615_5 gpc322 (
      {stage1_3[11], stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15]},
      {stage1_4[2]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[2],stage2_5[2],stage2_4[4],stage2_3[4]}
   );
   gpc606_5 gpc323 (
      {stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[3],stage2_6[3],stage2_5[3],stage2_4[5]}
   );
   gpc606_5 gpc324 (
      {stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[4],stage2_6[4],stage2_5[4],stage2_4[6]}
   );
   gpc606_5 gpc325 (
      {stage1_4[15], stage1_4[16], stage1_4[17], stage1_4[18], stage1_4[19], stage1_4[20]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[5],stage2_6[5],stage2_5[5],stage2_4[7]}
   );
   gpc606_5 gpc326 (
      {stage1_4[21], stage1_4[22], stage1_4[23], stage1_4[24], stage1_4[25], stage1_4[26]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[6],stage2_6[6],stage2_5[6],stage2_4[8]}
   );
   gpc606_5 gpc327 (
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[7],stage2_6[7],stage2_5[7],stage2_4[9]}
   );
   gpc606_5 gpc328 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[5],stage2_7[8],stage2_6[8],stage2_5[8]}
   );
   gpc615_5 gpc329 (
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[1],stage2_8[6],stage2_7[9]}
   );
   gpc615_5 gpc330 (
      {stage1_7[11], stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15]},
      {stage1_8[1]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[1],stage2_9[2],stage2_8[7],stage2_7[10]}
   );
   gpc606_5 gpc331 (
      {stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5], stage1_8[6], stage1_8[7]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[2],stage2_10[2],stage2_9[3],stage2_8[8]}
   );
   gpc606_5 gpc332 (
      {stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11], stage1_8[12], stage1_8[13]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[3],stage2_10[3],stage2_9[4],stage2_8[9]}
   );
   gpc606_5 gpc333 (
      {stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[4],stage2_10[4],stage2_9[5],stage2_8[10]}
   );
   gpc606_5 gpc334 (
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[3],stage2_11[5],stage2_10[5],stage2_9[6]}
   );
   gpc606_5 gpc335 (
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[4],stage2_11[6],stage2_10[6],stage2_9[7]}
   );
   gpc606_5 gpc336 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[5],stage2_11[7],stage2_10[7],stage2_9[8]}
   );
   gpc606_5 gpc337 (
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[6],stage2_11[8],stage2_10[8],stage2_9[9]}
   );
   gpc615_5 gpc338 (
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28]},
      {stage1_12[0]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[0],stage2_13[4],stage2_12[7],stage2_11[9]}
   );
   gpc606_5 gpc339 (
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[1],stage2_14[1],stage2_13[5],stage2_12[8]}
   );
   gpc606_5 gpc340 (
      {stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[2],stage2_14[2],stage2_13[6],stage2_12[9]}
   );
   gpc606_5 gpc341 (
      {stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[3],stage2_14[3],stage2_13[7],stage2_12[10]}
   );
   gpc606_5 gpc342 (
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[3],stage2_15[4],stage2_14[4],stage2_13[8]}
   );
   gpc606_5 gpc343 (
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[4],stage2_15[5],stage2_14[5],stage2_13[9]}
   );
   gpc606_5 gpc344 (
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[5],stage2_15[6],stage2_14[6],stage2_13[10]}
   );
   gpc1163_5 gpc345 (
      {stage1_14[18], stage1_14[19], stage1_14[20]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage1_16[0]},
      {stage1_17[0]},
      {stage2_18[0],stage2_17[3],stage2_16[6],stage2_15[7],stage2_14[7]}
   );
   gpc615_5 gpc346 (
      {stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25]},
      {stage1_15[24]},
      {stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage2_18[1],stage2_17[4],stage2_16[7],stage2_15[8],stage2_14[8]}
   );
   gpc615_5 gpc347 (
      {stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30]},
      {stage1_15[25]},
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12]},
      {stage2_18[2],stage2_17[5],stage2_16[8],stage2_15[9],stage2_14[9]}
   );
   gpc606_5 gpc348 (
      {stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17], stage1_16[18]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[0],stage2_18[3],stage2_17[6],stage2_16[9]}
   );
   gpc606_5 gpc349 (
      {stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23], stage1_16[24]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[1],stage2_18[4],stage2_17[7],stage2_16[10]}
   );
   gpc606_5 gpc350 (
      {stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5], stage1_17[6]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[5],stage2_17[8]}
   );
   gpc606_5 gpc351 (
      {stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11], stage1_17[12]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[3],stage2_19[3],stage2_18[6],stage2_17[9]}
   );
   gpc606_5 gpc352 (
      {stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17], stage1_17[18]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[4],stage2_19[4],stage2_18[7],stage2_17[10]}
   );
   gpc615_5 gpc353 (
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16]},
      {stage1_19[18]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[3],stage2_20[5],stage2_19[5],stage2_18[8]}
   );
   gpc615_5 gpc354 (
      {stage1_18[17], stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21]},
      {stage1_19[19]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[4],stage2_20[6],stage2_19[6],stage2_18[9]}
   );
   gpc615_5 gpc355 (
      {stage1_18[22], stage1_18[23], stage1_18[24], stage1_18[25], stage1_18[26]},
      {stage1_19[20]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[5],stage2_20[7],stage2_19[7],stage2_18[10]}
   );
   gpc606_5 gpc356 (
      {stage1_19[21], stage1_19[22], stage1_19[23], stage1_19[24], stage1_19[25], stage1_19[26]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[3],stage2_21[6],stage2_20[8],stage2_19[8]}
   );
   gpc606_5 gpc357 (
      {stage1_19[27], stage1_19[28], stage1_19[29], stage1_19[30], stage1_19[31], 1'b0},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[4],stage2_21[7],stage2_20[9],stage2_19[9]}
   );
   gpc606_5 gpc358 (
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], 1'b0},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[2],stage2_22[5],stage2_21[8],stage2_20[10]}
   );
   gpc606_5 gpc359 (
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[1],stage2_23[3],stage2_22[6],stage2_21[9]}
   );
   gpc606_5 gpc360 (
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[2],stage2_23[4],stage2_22[7],stage2_21[10]}
   );
   gpc606_5 gpc361 (
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[3],stage2_23[5],stage2_22[8],stage2_21[11]}
   );
   gpc615_5 gpc362 (
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10]},
      {stage1_23[18]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[3],stage2_24[4],stage2_23[6],stage2_22[9]}
   );
   gpc615_5 gpc363 (
      {stage1_22[11], stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15]},
      {stage1_23[19]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[4],stage2_24[5],stage2_23[7],stage2_22[10]}
   );
   gpc1415_5 gpc364 (
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4]},
      {stage1_26[0]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3]},
      {stage1_28[0]},
      {stage2_29[0],stage2_28[0],stage2_27[0],stage2_26[2],stage2_25[5]}
   );
   gpc615_5 gpc365 (
      {stage1_25[5], stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9]},
      {stage1_26[1]},
      {stage1_27[4], stage1_27[5], stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9]},
      {stage2_29[1],stage2_28[1],stage2_27[1],stage2_26[3],stage2_25[6]}
   );
   gpc615_5 gpc366 (
      {stage1_25[10], stage1_25[11], stage1_25[12], stage1_25[13], stage1_25[14]},
      {stage1_26[2]},
      {stage1_27[10], stage1_27[11], stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15]},
      {stage2_29[2],stage2_28[2],stage2_27[2],stage2_26[4],stage2_25[7]}
   );
   gpc615_5 gpc367 (
      {stage1_25[15], stage1_25[16], stage1_25[17], stage1_25[18], stage1_25[19]},
      {stage1_26[3]},
      {stage1_27[16], stage1_27[17], stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21]},
      {stage2_29[3],stage2_28[3],stage2_27[3],stage2_26[5],stage2_25[8]}
   );
   gpc615_5 gpc368 (
      {stage1_26[4], stage1_26[5], stage1_26[6], stage1_26[7], stage1_26[8]},
      {stage1_27[22]},
      {stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5], stage1_28[6]},
      {stage2_30[0],stage2_29[4],stage2_28[4],stage2_27[4],stage2_26[6]}
   );
   gpc615_5 gpc369 (
      {stage1_26[9], stage1_26[10], stage1_26[11], stage1_26[12], stage1_26[13]},
      {stage1_27[23]},
      {stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12]},
      {stage2_30[1],stage2_29[5],stage2_28[5],stage2_27[5],stage2_26[7]}
   );
   gpc615_5 gpc370 (
      {stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17], 1'b0},
      {stage1_27[24]},
      {stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17], stage1_28[18]},
      {stage2_30[2],stage2_29[6],stage2_28[6],stage2_27[6],stage2_26[8]}
   );
   gpc2135_5 gpc371 (
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4]},
      {stage1_30[0], stage1_30[1], stage1_30[2]},
      {stage1_31[0]},
      {stage1_32[0], stage1_32[1]},
      {stage2_33[0],stage2_32[0],stage2_31[0],stage2_30[3],stage2_29[7]}
   );
   gpc1406_5 gpc372 (
      {stage1_29[5], stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10]},
      {stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4]},
      {stage1_32[2]},
      {stage2_33[1],stage2_32[1],stage2_31[1],stage2_30[4],stage2_29[8]}
   );
   gpc606_5 gpc373 (
      {stage1_29[11], stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16]},
      {stage1_31[5], stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10]},
      {stage2_33[2],stage2_32[2],stage2_31[2],stage2_30[5],stage2_29[9]}
   );
   gpc606_5 gpc374 (
      {stage1_30[3], stage1_30[4], stage1_30[5], stage1_30[6], stage1_30[7], stage1_30[8]},
      {stage1_32[3], stage1_32[4], stage1_32[5], stage1_32[6], stage1_32[7], stage1_32[8]},
      {stage2_34[0],stage2_33[3],stage2_32[3],stage2_31[3],stage2_30[6]}
   );
   gpc606_5 gpc375 (
      {stage1_30[9], stage1_30[10], stage1_30[11], stage1_30[12], stage1_30[13], stage1_30[14]},
      {stage1_32[9], stage1_32[10], stage1_32[11], stage1_32[12], stage1_32[13], stage1_32[14]},
      {stage2_34[1],stage2_33[4],stage2_32[4],stage2_31[4],stage2_30[7]}
   );
   gpc615_5 gpc376 (
      {stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15]},
      {stage1_32[15]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[2],stage2_33[5],stage2_32[5],stage2_31[5]}
   );
   gpc615_5 gpc377 (
      {stage1_31[16], stage1_31[17], stage1_31[18], stage1_31[19], stage1_31[20]},
      {stage1_32[16]},
      {stage1_33[6], stage1_33[7], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage2_35[1],stage2_34[3],stage2_33[6],stage2_32[6],stage2_31[6]}
   );
   gpc1_1 gpc378 (
      {stage1_0[8]},
      {stage2_0[2]}
   );
   gpc1_1 gpc379 (
      {stage1_0[9]},
      {stage2_0[3]}
   );
   gpc1_1 gpc380 (
      {stage1_0[10]},
      {stage2_0[4]}
   );
   gpc1_1 gpc381 (
      {stage1_0[11]},
      {stage2_0[5]}
   );
   gpc1_1 gpc382 (
      {stage1_0[12]},
      {stage2_0[6]}
   );
   gpc1_1 gpc383 (
      {stage1_0[13]},
      {stage2_0[7]}
   );
   gpc1_1 gpc384 (
      {stage1_0[14]},
      {stage2_0[8]}
   );
   gpc1_1 gpc385 (
      {stage1_0[15]},
      {stage2_0[9]}
   );
   gpc1_1 gpc386 (
      {stage1_1[7]},
      {stage2_1[2]}
   );
   gpc1_1 gpc387 (
      {stage1_1[8]},
      {stage2_1[3]}
   );
   gpc1_1 gpc388 (
      {stage1_1[9]},
      {stage2_1[4]}
   );
   gpc1_1 gpc389 (
      {stage1_1[10]},
      {stage2_1[5]}
   );
   gpc1_1 gpc390 (
      {stage1_1[11]},
      {stage2_1[6]}
   );
   gpc1_1 gpc391 (
      {stage1_1[12]},
      {stage2_1[7]}
   );
   gpc1_1 gpc392 (
      {stage1_1[13]},
      {stage2_1[8]}
   );
   gpc1_1 gpc393 (
      {stage1_1[14]},
      {stage2_1[9]}
   );
   gpc1_1 gpc394 (
      {stage1_1[15]},
      {stage2_1[10]}
   );
   gpc1_1 gpc395 (
      {stage1_1[16]},
      {stage2_1[11]}
   );
   gpc1_1 gpc396 (
      {stage1_2[7]},
      {stage2_2[2]}
   );
   gpc1_1 gpc397 (
      {stage1_2[8]},
      {stage2_2[3]}
   );
   gpc1_1 gpc398 (
      {stage1_2[9]},
      {stage2_2[4]}
   );
   gpc1_1 gpc399 (
      {stage1_2[10]},
      {stage2_2[5]}
   );
   gpc1_1 gpc400 (
      {stage1_2[11]},
      {stage2_2[6]}
   );
   gpc1_1 gpc401 (
      {stage1_2[12]},
      {stage2_2[7]}
   );
   gpc1_1 gpc402 (
      {stage1_2[13]},
      {stage2_2[8]}
   );
   gpc1_1 gpc403 (
      {stage1_2[14]},
      {stage2_2[9]}
   );
   gpc1_1 gpc404 (
      {stage1_2[15]},
      {stage2_2[10]}
   );
   gpc1_1 gpc405 (
      {stage1_2[16]},
      {stage2_2[11]}
   );
   gpc1_1 gpc406 (
      {stage1_2[17]},
      {stage2_2[12]}
   );
   gpc1_1 gpc407 (
      {stage1_2[18]},
      {stage2_2[13]}
   );
   gpc1_1 gpc408 (
      {stage1_2[19]},
      {stage2_2[14]}
   );
   gpc1_1 gpc409 (
      {stage1_2[20]},
      {stage2_2[15]}
   );
   gpc1_1 gpc410 (
      {stage1_2[21]},
      {stage2_2[16]}
   );
   gpc1_1 gpc411 (
      {stage1_3[16]},
      {stage2_3[5]}
   );
   gpc1_1 gpc412 (
      {stage1_3[17]},
      {stage2_3[6]}
   );
   gpc1_1 gpc413 (
      {stage1_3[18]},
      {stage2_3[7]}
   );
   gpc1_1 gpc414 (
      {stage1_3[19]},
      {stage2_3[8]}
   );
   gpc1_1 gpc415 (
      {stage1_3[20]},
      {stage2_3[9]}
   );
   gpc1_1 gpc416 (
      {stage1_3[21]},
      {stage2_3[10]}
   );
   gpc1_1 gpc417 (
      {stage1_5[24]},
      {stage2_5[9]}
   );
   gpc1_1 gpc418 (
      {stage1_5[25]},
      {stage2_5[10]}
   );
   gpc1_1 gpc419 (
      {stage1_5[26]},
      {stage2_5[11]}
   );
   gpc1_1 gpc420 (
      {stage1_6[30]},
      {stage2_6[9]}
   );
   gpc1_1 gpc421 (
      {stage1_6[31]},
      {stage2_6[10]}
   );
   gpc1_1 gpc422 (
      {stage1_6[32]},
      {stage2_6[11]}
   );
   gpc1_1 gpc423 (
      {stage1_7[16]},
      {stage2_7[11]}
   );
   gpc1_1 gpc424 (
      {stage1_7[17]},
      {stage2_7[12]}
   );
   gpc1_1 gpc425 (
      {stage1_7[18]},
      {stage2_7[13]}
   );
   gpc1_1 gpc426 (
      {stage1_7[19]},
      {stage2_7[14]}
   );
   gpc1_1 gpc427 (
      {stage1_7[20]},
      {stage2_7[15]}
   );
   gpc1_1 gpc428 (
      {stage1_8[20]},
      {stage2_8[11]}
   );
   gpc1_1 gpc429 (
      {stage1_8[21]},
      {stage2_8[12]}
   );
   gpc1_1 gpc430 (
      {stage1_8[22]},
      {stage2_8[13]}
   );
   gpc1_1 gpc431 (
      {stage1_8[23]},
      {stage2_8[14]}
   );
   gpc1_1 gpc432 (
      {stage1_8[24]},
      {stage2_8[15]}
   );
   gpc1_1 gpc433 (
      {stage1_8[25]},
      {stage2_8[16]}
   );
   gpc1_1 gpc434 (
      {stage1_12[19]},
      {stage2_12[11]}
   );
   gpc1_1 gpc435 (
      {stage1_12[20]},
      {stage2_12[12]}
   );
   gpc1_1 gpc436 (
      {stage1_12[21]},
      {stage2_12[13]}
   );
   gpc1_1 gpc437 (
      {stage1_12[22]},
      {stage2_12[14]}
   );
   gpc1_1 gpc438 (
      {stage1_12[23]},
      {stage2_12[15]}
   );
   gpc1_1 gpc439 (
      {stage1_13[24]},
      {stage2_13[11]}
   );
   gpc1_1 gpc440 (
      {stage1_13[25]},
      {stage2_13[12]}
   );
   gpc1_1 gpc441 (
      {stage1_13[26]},
      {stage2_13[13]}
   );
   gpc1_1 gpc442 (
      {stage1_13[27]},
      {stage2_13[14]}
   );
   gpc1_1 gpc443 (
      {stage1_13[28]},
      {stage2_13[15]}
   );
   gpc1_1 gpc444 (
      {stage1_13[29]},
      {stage2_13[16]}
   );
   gpc1_1 gpc445 (
      {stage1_13[30]},
      {stage2_13[17]}
   );
   gpc1_1 gpc446 (
      {stage1_13[31]},
      {stage2_13[18]}
   );
   gpc1_1 gpc447 (
      {stage1_15[26]},
      {stage2_15[10]}
   );
   gpc1_1 gpc448 (
      {stage1_15[27]},
      {stage2_15[11]}
   );
   gpc1_1 gpc449 (
      {stage1_17[19]},
      {stage2_17[11]}
   );
   gpc1_1 gpc450 (
      {stage1_18[27]},
      {stage2_18[11]}
   );
   gpc1_1 gpc451 (
      {stage1_18[28]},
      {stage2_18[12]}
   );
   gpc1_1 gpc452 (
      {stage1_18[29]},
      {stage2_18[13]}
   );
   gpc1_1 gpc453 (
      {stage1_22[16]},
      {stage2_22[11]}
   );
   gpc1_1 gpc454 (
      {stage1_22[17]},
      {stage2_22[12]}
   );
   gpc1_1 gpc455 (
      {stage1_22[18]},
      {stage2_22[13]}
   );
   gpc1_1 gpc456 (
      {stage1_22[19]},
      {stage2_22[14]}
   );
   gpc1_1 gpc457 (
      {stage1_22[20]},
      {stage2_22[15]}
   );
   gpc1_1 gpc458 (
      {stage1_22[21]},
      {stage2_22[16]}
   );
   gpc1_1 gpc459 (
      {stage1_23[20]},
      {stage2_23[8]}
   );
   gpc1_1 gpc460 (
      {stage1_23[21]},
      {stage2_23[9]}
   );
   gpc1_1 gpc461 (
      {stage1_23[22]},
      {stage2_23[10]}
   );
   gpc1_1 gpc462 (
      {stage1_23[23]},
      {stage2_23[11]}
   );
   gpc1_1 gpc463 (
      {stage1_23[24]},
      {stage2_23[12]}
   );
   gpc1_1 gpc464 (
      {stage1_23[25]},
      {stage2_23[13]}
   );
   gpc1_1 gpc465 (
      {stage1_23[26]},
      {stage2_23[14]}
   );
   gpc1_1 gpc466 (
      {stage1_23[27]},
      {stage2_23[15]}
   );
   gpc1_1 gpc467 (
      {stage1_23[28]},
      {stage2_23[16]}
   );
   gpc1_1 gpc468 (
      {stage1_24[12]},
      {stage2_24[6]}
   );
   gpc1_1 gpc469 (
      {stage1_24[13]},
      {stage2_24[7]}
   );
   gpc1_1 gpc470 (
      {stage1_24[14]},
      {stage2_24[8]}
   );
   gpc1_1 gpc471 (
      {stage1_24[15]},
      {stage2_24[9]}
   );
   gpc1_1 gpc472 (
      {stage1_24[16]},
      {stage2_24[10]}
   );
   gpc1_1 gpc473 (
      {stage1_24[17]},
      {stage2_24[11]}
   );
   gpc1_1 gpc474 (
      {stage1_24[18]},
      {stage2_24[12]}
   );
   gpc1_1 gpc475 (
      {stage1_24[19]},
      {stage2_24[13]}
   );
   gpc1_1 gpc476 (
      {stage1_24[20]},
      {stage2_24[14]}
   );
   gpc1_1 gpc477 (
      {stage1_24[21]},
      {stage2_24[15]}
   );
   gpc1_1 gpc478 (
      {stage1_24[22]},
      {stage2_24[16]}
   );
   gpc1_1 gpc479 (
      {stage1_24[23]},
      {stage2_24[17]}
   );
   gpc1_1 gpc480 (
      {stage1_25[20]},
      {stage2_25[9]}
   );
   gpc1_1 gpc481 (
      {stage1_25[21]},
      {stage2_25[10]}
   );
   gpc1_1 gpc482 (
      {stage1_25[22]},
      {stage2_25[11]}
   );
   gpc1_1 gpc483 (
      {stage1_28[19]},
      {stage2_28[7]}
   );
   gpc1_1 gpc484 (
      {stage1_28[20]},
      {stage2_28[8]}
   );
   gpc1_1 gpc485 (
      {stage1_28[21]},
      {stage2_28[9]}
   );
   gpc1_1 gpc486 (
      {stage1_28[22]},
      {stage2_28[10]}
   );
   gpc1_1 gpc487 (
      {stage1_28[23]},
      {stage2_28[11]}
   );
   gpc1_1 gpc488 (
      {stage1_28[24]},
      {stage2_28[12]}
   );
   gpc1_1 gpc489 (
      {stage1_28[25]},
      {stage2_28[13]}
   );
   gpc1_1 gpc490 (
      {stage1_29[17]},
      {stage2_29[10]}
   );
   gpc1_1 gpc491 (
      {stage1_29[18]},
      {stage2_29[11]}
   );
   gpc1_1 gpc492 (
      {stage1_29[19]},
      {stage2_29[12]}
   );
   gpc1_1 gpc493 (
      {stage1_29[20]},
      {stage2_29[13]}
   );
   gpc1_1 gpc494 (
      {stage1_29[21]},
      {stage2_29[14]}
   );
   gpc1_1 gpc495 (
      {stage1_29[22]},
      {stage2_29[15]}
   );
   gpc1_1 gpc496 (
      {stage1_29[23]},
      {stage2_29[16]}
   );
   gpc1_1 gpc497 (
      {stage1_29[24]},
      {stage2_29[17]}
   );
   gpc1_1 gpc498 (
      {stage1_30[15]},
      {stage2_30[8]}
   );
   gpc1_1 gpc499 (
      {stage1_30[16]},
      {stage2_30[9]}
   );
   gpc1_1 gpc500 (
      {stage1_30[17]},
      {stage2_30[10]}
   );
   gpc1_1 gpc501 (
      {stage1_31[21]},
      {stage2_31[7]}
   );
   gpc1_1 gpc502 (
      {stage1_31[22]},
      {stage2_31[8]}
   );
   gpc1_1 gpc503 (
      {stage1_31[23]},
      {stage2_31[9]}
   );
   gpc615_5 gpc504 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc505 (
      {stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9]},
      {stage2_1[1]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc506 (
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16]},
      {stage2_3[0]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc1163_5 gpc507 (
      {stage2_4[6], stage2_4[7], stage2_4[8]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage2_6[0]},
      {stage2_7[0]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[1],stage3_4[3]}
   );
   gpc606_5 gpc508 (
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6]},
      {stage3_9[0],stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[2]}
   );
   gpc606_5 gpc509 (
      {stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[1],stage3_8[2],stage3_7[2],stage3_6[3]}
   );
   gpc606_5 gpc510 (
      {stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11], 1'b0},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[2],stage3_8[3],stage3_7[3],stage3_6[4]}
   );
   gpc615_5 gpc511 (
      {stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage2_8[12]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[3],stage3_8[4],stage3_7[4]}
   );
   gpc606_5 gpc512 (
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[0],stage3_11[1],stage3_10[3]}
   );
   gpc615_5 gpc513 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[1],stage3_12[1],stage3_11[2]}
   );
   gpc615_5 gpc514 (
      {stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9]},
      {stage2_12[7]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[2],stage3_13[2],stage3_12[2],stage3_11[3]}
   );
   gpc606_5 gpc515 (
      {stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[2],stage3_14[3],stage3_13[3],stage3_12[3]}
   );
   gpc135_4 gpc516 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16]},
      {stage2_14[6], stage2_14[7], stage2_14[8]},
      {stage2_15[0]},
      {stage3_16[1],stage3_15[3],stage3_14[4],stage3_13[4]}
   );
   gpc606_5 gpc517 (
      {stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[0],stage3_17[0],stage3_16[2],stage3_15[4]}
   );
   gpc615_5 gpc518 (
      {stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage2_16[0]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[1],stage3_17[1],stage3_16[3],stage3_15[5]}
   );
   gpc606_5 gpc519 (
      {stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[2],stage3_18[2],stage3_17[2],stage3_16[4]}
   );
   gpc1343_5 gpc520 (
      {stage2_18[6], stage2_18[7], stage2_18[8]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3]},
      {stage2_20[0], stage2_20[1], stage2_20[2]},
      {stage2_21[0]},
      {stage3_22[0],stage3_21[0],stage3_20[1],stage3_19[3],stage3_18[3]}
   );
   gpc1343_5 gpc521 (
      {stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage2_19[4], stage2_19[5], stage2_19[6], stage2_19[7]},
      {stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage2_21[1]},
      {stage3_22[1],stage3_21[1],stage3_20[2],stage3_19[4],stage3_18[4]}
   );
   gpc606_5 gpc522 (
      {stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5], stage2_21[6], stage2_21[7]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[2],stage3_21[2]}
   );
   gpc615_5 gpc523 (
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4]},
      {stage2_23[6]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[3]}
   );
   gpc615_5 gpc524 (
      {stage2_22[5], stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9]},
      {stage2_23[7]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[4]}
   );
   gpc615_5 gpc525 (
      {stage2_22[10], stage2_22[11], stage2_22[12], stage2_22[13], stage2_22[14]},
      {stage2_23[8]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[5]}
   );
   gpc606_5 gpc526 (
      {stage2_23[9], stage2_23[10], stage2_23[11], stage2_23[12], stage2_23[13], stage2_23[14]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[3],stage3_25[4],stage3_24[4],stage3_23[4]}
   );
   gpc606_5 gpc527 (
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[0],stage3_27[1],stage3_26[4],stage3_25[5]}
   );
   gpc1415_5 gpc528 (
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4]},
      {stage2_27[6]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3]},
      {stage2_29[0]},
      {stage3_30[0],stage3_29[1],stage3_28[1],stage3_27[2],stage3_26[5]}
   );
   gpc615_5 gpc529 (
      {stage2_28[4], stage2_28[5], stage2_28[6], stage2_28[7], stage2_28[8]},
      {stage2_29[1]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[0],stage3_30[1],stage3_29[2],stage3_28[2]}
   );
   gpc615_5 gpc530 (
      {stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13]},
      {stage2_29[2]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], 1'b0},
      {stage3_32[1],stage3_31[1],stage3_30[2],stage3_29[3],stage3_28[3]}
   );
   gpc606_5 gpc531 (
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[0],stage3_33[0],stage3_32[2],stage3_31[2]}
   );
   gpc117_4 gpc532 (
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5], stage2_32[6]},
      {stage2_33[6]},
      {stage2_34[0]},
      {stage3_35[1],stage3_34[1],stage3_33[1],stage3_32[3]}
   );
   gpc1_1 gpc533 (
      {stage2_1[2]},
      {stage3_1[2]}
   );
   gpc1_1 gpc534 (
      {stage2_1[3]},
      {stage3_1[3]}
   );
   gpc1_1 gpc535 (
      {stage2_1[4]},
      {stage3_1[4]}
   );
   gpc1_1 gpc536 (
      {stage2_1[5]},
      {stage3_1[5]}
   );
   gpc1_1 gpc537 (
      {stage2_1[6]},
      {stage3_1[6]}
   );
   gpc1_1 gpc538 (
      {stage2_1[7]},
      {stage3_1[7]}
   );
   gpc1_1 gpc539 (
      {stage2_1[8]},
      {stage3_1[8]}
   );
   gpc1_1 gpc540 (
      {stage2_1[9]},
      {stage3_1[9]}
   );
   gpc1_1 gpc541 (
      {stage2_1[10]},
      {stage3_1[10]}
   );
   gpc1_1 gpc542 (
      {stage2_1[11]},
      {stage3_1[11]}
   );
   gpc1_1 gpc543 (
      {stage2_3[1]},
      {stage3_3[3]}
   );
   gpc1_1 gpc544 (
      {stage2_3[2]},
      {stage3_3[4]}
   );
   gpc1_1 gpc545 (
      {stage2_3[3]},
      {stage3_3[5]}
   );
   gpc1_1 gpc546 (
      {stage2_3[4]},
      {stage3_3[6]}
   );
   gpc1_1 gpc547 (
      {stage2_3[5]},
      {stage3_3[7]}
   );
   gpc1_1 gpc548 (
      {stage2_3[6]},
      {stage3_3[8]}
   );
   gpc1_1 gpc549 (
      {stage2_3[7]},
      {stage3_3[9]}
   );
   gpc1_1 gpc550 (
      {stage2_3[8]},
      {stage3_3[10]}
   );
   gpc1_1 gpc551 (
      {stage2_3[9]},
      {stage3_3[11]}
   );
   gpc1_1 gpc552 (
      {stage2_3[10]},
      {stage3_3[12]}
   );
   gpc1_1 gpc553 (
      {stage2_4[9]},
      {stage3_4[4]}
   );
   gpc1_1 gpc554 (
      {stage2_7[12]},
      {stage3_7[5]}
   );
   gpc1_1 gpc555 (
      {stage2_7[13]},
      {stage3_7[6]}
   );
   gpc1_1 gpc556 (
      {stage2_7[14]},
      {stage3_7[7]}
   );
   gpc1_1 gpc557 (
      {stage2_7[15]},
      {stage3_7[8]}
   );
   gpc1_1 gpc558 (
      {stage2_8[13]},
      {stage3_8[5]}
   );
   gpc1_1 gpc559 (
      {stage2_8[14]},
      {stage3_8[6]}
   );
   gpc1_1 gpc560 (
      {stage2_8[15]},
      {stage3_8[7]}
   );
   gpc1_1 gpc561 (
      {stage2_8[16]},
      {stage3_8[8]}
   );
   gpc1_1 gpc562 (
      {stage2_9[6]},
      {stage3_9[4]}
   );
   gpc1_1 gpc563 (
      {stage2_9[7]},
      {stage3_9[5]}
   );
   gpc1_1 gpc564 (
      {stage2_9[8]},
      {stage3_9[6]}
   );
   gpc1_1 gpc565 (
      {stage2_9[9]},
      {stage3_9[7]}
   );
   gpc1_1 gpc566 (
      {stage2_10[6]},
      {stage3_10[4]}
   );
   gpc1_1 gpc567 (
      {stage2_10[7]},
      {stage3_10[5]}
   );
   gpc1_1 gpc568 (
      {stage2_10[8]},
      {stage3_10[6]}
   );
   gpc1_1 gpc569 (
      {stage2_12[14]},
      {stage3_12[4]}
   );
   gpc1_1 gpc570 (
      {stage2_12[15]},
      {stage3_12[5]}
   );
   gpc1_1 gpc571 (
      {stage2_13[17]},
      {stage3_13[5]}
   );
   gpc1_1 gpc572 (
      {stage2_13[18]},
      {stage3_13[6]}
   );
   gpc1_1 gpc573 (
      {stage2_14[9]},
      {stage3_14[5]}
   );
   gpc1_1 gpc574 (
      {stage2_16[7]},
      {stage3_16[5]}
   );
   gpc1_1 gpc575 (
      {stage2_16[8]},
      {stage3_16[6]}
   );
   gpc1_1 gpc576 (
      {stage2_16[9]},
      {stage3_16[7]}
   );
   gpc1_1 gpc577 (
      {stage2_16[10]},
      {stage3_16[8]}
   );
   gpc1_1 gpc578 (
      {stage2_18[12]},
      {stage3_18[5]}
   );
   gpc1_1 gpc579 (
      {stage2_18[13]},
      {stage3_18[6]}
   );
   gpc1_1 gpc580 (
      {stage2_19[8]},
      {stage3_19[5]}
   );
   gpc1_1 gpc581 (
      {stage2_19[9]},
      {stage3_19[6]}
   );
   gpc1_1 gpc582 (
      {stage2_20[6]},
      {stage3_20[3]}
   );
   gpc1_1 gpc583 (
      {stage2_20[7]},
      {stage3_20[4]}
   );
   gpc1_1 gpc584 (
      {stage2_20[8]},
      {stage3_20[5]}
   );
   gpc1_1 gpc585 (
      {stage2_20[9]},
      {stage3_20[6]}
   );
   gpc1_1 gpc586 (
      {stage2_20[10]},
      {stage3_20[7]}
   );
   gpc1_1 gpc587 (
      {stage2_21[8]},
      {stage3_21[3]}
   );
   gpc1_1 gpc588 (
      {stage2_21[9]},
      {stage3_21[4]}
   );
   gpc1_1 gpc589 (
      {stage2_21[10]},
      {stage3_21[5]}
   );
   gpc1_1 gpc590 (
      {stage2_21[11]},
      {stage3_21[6]}
   );
   gpc1_1 gpc591 (
      {stage2_22[15]},
      {stage3_22[6]}
   );
   gpc1_1 gpc592 (
      {stage2_22[16]},
      {stage3_22[7]}
   );
   gpc1_1 gpc593 (
      {stage2_23[15]},
      {stage3_23[5]}
   );
   gpc1_1 gpc594 (
      {stage2_23[16]},
      {stage3_23[6]}
   );
   gpc1_1 gpc595 (
      {stage2_26[5]},
      {stage3_26[6]}
   );
   gpc1_1 gpc596 (
      {stage2_26[6]},
      {stage3_26[7]}
   );
   gpc1_1 gpc597 (
      {stage2_26[7]},
      {stage3_26[8]}
   );
   gpc1_1 gpc598 (
      {stage2_26[8]},
      {stage3_26[9]}
   );
   gpc1_1 gpc599 (
      {stage2_29[3]},
      {stage3_29[4]}
   );
   gpc1_1 gpc600 (
      {stage2_29[4]},
      {stage3_29[5]}
   );
   gpc1_1 gpc601 (
      {stage2_29[5]},
      {stage3_29[6]}
   );
   gpc1_1 gpc602 (
      {stage2_29[6]},
      {stage3_29[7]}
   );
   gpc1_1 gpc603 (
      {stage2_29[7]},
      {stage3_29[8]}
   );
   gpc1_1 gpc604 (
      {stage2_29[8]},
      {stage3_29[9]}
   );
   gpc1_1 gpc605 (
      {stage2_29[9]},
      {stage3_29[10]}
   );
   gpc1_1 gpc606 (
      {stage2_29[10]},
      {stage3_29[11]}
   );
   gpc1_1 gpc607 (
      {stage2_29[11]},
      {stage3_29[12]}
   );
   gpc1_1 gpc608 (
      {stage2_29[12]},
      {stage3_29[13]}
   );
   gpc1_1 gpc609 (
      {stage2_29[13]},
      {stage3_29[14]}
   );
   gpc1_1 gpc610 (
      {stage2_29[14]},
      {stage3_29[15]}
   );
   gpc1_1 gpc611 (
      {stage2_29[15]},
      {stage3_29[16]}
   );
   gpc1_1 gpc612 (
      {stage2_29[16]},
      {stage3_29[17]}
   );
   gpc1_1 gpc613 (
      {stage2_29[17]},
      {stage3_29[18]}
   );
   gpc1_1 gpc614 (
      {stage2_31[6]},
      {stage3_31[3]}
   );
   gpc1_1 gpc615 (
      {stage2_31[7]},
      {stage3_31[4]}
   );
   gpc1_1 gpc616 (
      {stage2_31[8]},
      {stage3_31[5]}
   );
   gpc1_1 gpc617 (
      {stage2_31[9]},
      {stage3_31[6]}
   );
   gpc1_1 gpc618 (
      {stage2_34[1]},
      {stage3_34[2]}
   );
   gpc1_1 gpc619 (
      {stage2_34[2]},
      {stage3_34[3]}
   );
   gpc1_1 gpc620 (
      {stage2_34[3]},
      {stage3_34[4]}
   );
   gpc1_1 gpc621 (
      {stage2_35[0]},
      {stage3_35[2]}
   );
   gpc1_1 gpc622 (
      {stage2_35[1]},
      {stage3_35[3]}
   );
   gpc615_5 gpc623 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4]},
      {stage3_2[0]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc615_5 gpc624 (
      {stage3_1[5], stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9]},
      {stage3_2[1]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc2135_5 gpc625 (
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4]},
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[0]},
      {stage3_7[0], stage3_7[1]},
      {stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[2],stage4_4[2]}
   );
   gpc623_5 gpc626 (
      {stage3_6[1], stage3_6[2], stage3_6[3]},
      {stage3_7[2], stage3_7[3]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[1]}
   );
   gpc615_5 gpc627 (
      {stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7], stage3_7[8]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[2]}
   );
   gpc615_5 gpc628 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4]},
      {stage3_11[0]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[2]}
   );
   gpc623_5 gpc629 (
      {stage3_11[1], stage3_11[2], stage3_11[3]},
      {1'b0, 1'b0},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1],stage4_11[2]}
   );
   gpc1406_5 gpc630 (
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3]},
      {stage3_17[0]},
      {stage4_18[0],stage4_17[0],stage4_16[0],stage4_15[1],stage4_14[2]}
   );
   gpc215_4 gpc631 (
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4]},
      {stage3_16[4]},
      {stage3_17[1], stage3_17[2]},
      {stage4_18[1],stage4_17[1],stage4_16[1],stage4_15[2]}
   );
   gpc606_5 gpc632 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage4_22[0],stage4_21[0],stage4_20[0],stage4_19[0],stage4_18[2]}
   );
   gpc117_4 gpc633 (
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6]},
      {stage3_20[6]},
      {stage3_21[0]},
      {stage4_22[1],stage4_21[1],stage4_20[1],stage4_19[1]}
   );
   gpc606_5 gpc634 (
      {stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5], stage3_21[6]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[0],stage4_23[0],stage4_22[2],stage4_21[2]}
   );
   gpc606_5 gpc635 (
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], 1'b0},
      {stage4_26[0],stage4_25[1],stage4_24[1],stage4_23[1],stage4_22[3]}
   );
   gpc1343_5 gpc636 (
      {stage3_25[0], stage3_25[1], stage3_25[2]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3]},
      {stage3_27[0], stage3_27[1], stage3_27[2]},
      {stage3_28[0]},
      {stage4_29[0],stage4_28[0],stage4_27[0],stage4_26[1],stage4_25[2]}
   );
   gpc135_4 gpc637 (
      {stage3_28[1], stage3_28[2], stage3_28[3], 1'b0, 1'b0},
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[0]},
      {stage4_31[0],stage4_30[0],stage4_29[1],stage4_28[1]}
   );
   gpc207_4 gpc638 (
      {stage3_29[3], stage3_29[4], stage3_29[5], stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9]},
      {stage3_31[0], stage3_31[1]},
      {stage4_32[0],stage4_31[1],stage4_30[1],stage4_29[2]}
   );
   gpc207_4 gpc639 (
      {stage3_29[10], stage3_29[11], stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16]},
      {stage3_31[2], stage3_31[3]},
      {stage4_32[1],stage4_31[2],stage4_30[2],stage4_29[3]}
   );
   gpc623_5 gpc640 (
      {stage3_32[0], stage3_32[1], stage3_32[2]},
      {stage3_33[0], stage3_33[1]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], 1'b0},
      {stage4_36[0],stage4_35[0],stage4_34[0],stage4_33[0],stage4_32[2]}
   );
   gpc215_4 gpc641 (
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], 1'b0},
      {1'b0},
      {1'b0, 1'b0},
      {stage4_37[0],stage4_36[1],stage4_35[1]}
   );
   gpc1_1 gpc642 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc643 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc644 (
      {stage3_1[10]},
      {stage4_1[2]}
   );
   gpc1_1 gpc645 (
      {stage3_1[11]},
      {stage4_1[3]}
   );
   gpc1_1 gpc646 (
      {stage3_2[2]},
      {stage4_2[2]}
   );
   gpc1_1 gpc647 (
      {stage3_3[12]},
      {stage4_3[2]}
   );
   gpc1_1 gpc648 (
      {stage3_6[4]},
      {stage4_6[2]}
   );
   gpc1_1 gpc649 (
      {stage3_8[7]},
      {stage4_8[3]}
   );
   gpc1_1 gpc650 (
      {stage3_8[8]},
      {stage4_8[4]}
   );
   gpc1_1 gpc651 (
      {stage3_9[6]},
      {stage4_9[2]}
   );
   gpc1_1 gpc652 (
      {stage3_9[7]},
      {stage4_9[3]}
   );
   gpc1_1 gpc653 (
      {stage3_10[5]},
      {stage4_10[3]}
   );
   gpc1_1 gpc654 (
      {stage3_10[6]},
      {stage4_10[4]}
   );
   gpc1_1 gpc655 (
      {stage3_13[6]},
      {stage4_13[2]}
   );
   gpc1_1 gpc656 (
      {stage3_15[5]},
      {stage4_15[3]}
   );
   gpc1_1 gpc657 (
      {stage3_16[5]},
      {stage4_16[2]}
   );
   gpc1_1 gpc658 (
      {stage3_16[6]},
      {stage4_16[3]}
   );
   gpc1_1 gpc659 (
      {stage3_16[7]},
      {stage4_16[4]}
   );
   gpc1_1 gpc660 (
      {stage3_16[8]},
      {stage4_16[5]}
   );
   gpc1_1 gpc661 (
      {stage3_18[6]},
      {stage4_18[3]}
   );
   gpc1_1 gpc662 (
      {stage3_20[7]},
      {stage4_20[2]}
   );
   gpc1_1 gpc663 (
      {stage3_22[6]},
      {stage4_22[4]}
   );
   gpc1_1 gpc664 (
      {stage3_22[7]},
      {stage4_22[5]}
   );
   gpc1_1 gpc665 (
      {stage3_23[6]},
      {stage4_23[2]}
   );
   gpc1_1 gpc666 (
      {stage3_25[3]},
      {stage4_25[3]}
   );
   gpc1_1 gpc667 (
      {stage3_25[4]},
      {stage4_25[4]}
   );
   gpc1_1 gpc668 (
      {stage3_25[5]},
      {stage4_25[5]}
   );
   gpc1_1 gpc669 (
      {stage3_26[4]},
      {stage4_26[2]}
   );
   gpc1_1 gpc670 (
      {stage3_26[5]},
      {stage4_26[3]}
   );
   gpc1_1 gpc671 (
      {stage3_26[6]},
      {stage4_26[4]}
   );
   gpc1_1 gpc672 (
      {stage3_26[7]},
      {stage4_26[5]}
   );
   gpc1_1 gpc673 (
      {stage3_26[8]},
      {stage4_26[6]}
   );
   gpc1_1 gpc674 (
      {stage3_26[9]},
      {stage4_26[7]}
   );
   gpc1_1 gpc675 (
      {stage3_29[17]},
      {stage4_29[4]}
   );
   gpc1_1 gpc676 (
      {stage3_29[18]},
      {stage4_29[5]}
   );
   gpc1_1 gpc677 (
      {stage3_30[1]},
      {stage4_30[3]}
   );
   gpc1_1 gpc678 (
      {stage3_30[2]},
      {stage4_30[4]}
   );
   gpc1_1 gpc679 (
      {stage3_31[4]},
      {stage4_31[3]}
   );
   gpc1_1 gpc680 (
      {stage3_31[5]},
      {stage4_31[4]}
   );
   gpc1_1 gpc681 (
      {stage3_31[6]},
      {stage4_31[5]}
   );
   gpc1_1 gpc682 (
      {stage3_32[3]},
      {stage4_32[3]}
   );
   gpc23_3 gpc683 (
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0], stage4_2[1]},
      {stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc2223_5 gpc684 (
      {stage4_3[0], stage4_3[1], stage4_3[2]},
      {stage4_4[0], stage4_4[1]},
      {stage4_5[0], stage4_5[1]},
      {stage4_6[0], stage4_6[1]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[1]}
   );
   gpc1343_5 gpc685 (
      {stage4_7[0], stage4_7[1], stage4_7[2]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3]},
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[1]}
   );
   gpc135_4 gpc686 (
      {stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], 1'b0},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[1],stage5_10[1]}
   );
   gpc1423_5 gpc687 (
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0], stage4_14[1]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3]},
      {stage4_16[0]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[1]}
   );
   gpc1325_5 gpc688 (
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage4_17[0], stage4_17[1]},
      {stage4_18[0], stage4_18[1], stage4_18[2]},
      {stage4_19[0]},
      {stage5_20[0],stage5_19[0],stage5_18[0],stage5_17[1],stage5_16[1]}
   );
   gpc1343_5 gpc689 (
      {stage4_20[0], stage4_20[1], stage4_20[2]},
      {stage4_21[0], stage4_21[1], stage4_21[2], 1'b0},
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[0]},
      {stage5_24[0],stage5_23[0],stage5_22[0],stage5_21[0],stage5_20[1]}
   );
   gpc223_4 gpc690 (
      {stage4_22[3], stage4_22[4], stage4_22[5]},
      {stage4_23[1], stage4_23[2]},
      {stage4_24[0], stage4_24[1]},
      {stage5_25[0],stage5_24[1],stage5_23[1],stage5_22[1]}
   );
   gpc2116_5 gpc691 (
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage4_26[0]},
      {stage4_27[0]},
      {stage4_28[0], stage4_28[1]},
      {stage5_29[0],stage5_28[0],stage5_27[0],stage5_26[0],stage5_25[1]}
   );
   gpc7_3 gpc692 (
      {stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5], stage4_26[6], stage4_26[7]},
      {stage5_28[1],stage5_27[1],stage5_26[1]}
   );
   gpc606_5 gpc693 (
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[0],stage5_29[1]}
   );
   gpc1415_5 gpc694 (
      {stage4_30[0], stage4_30[1], stage4_30[2], stage4_30[3], stage4_30[4]},
      {1'b0},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3]},
      {stage4_33[0]},
      {stage5_34[0],stage5_33[1],stage5_32[1],stage5_31[1],stage5_30[1]}
   );
   gpc1_1 gpc695 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc696 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc697 (
      {stage4_1[3]},
      {stage5_1[1]}
   );
   gpc1_1 gpc698 (
      {stage4_2[2]},
      {stage5_2[1]}
   );
   gpc1_1 gpc699 (
      {stage4_4[2]},
      {stage5_4[1]}
   );
   gpc1_1 gpc700 (
      {stage4_5[2]},
      {stage5_5[1]}
   );
   gpc1_1 gpc701 (
      {stage4_6[2]},
      {stage5_6[1]}
   );
   gpc1_1 gpc702 (
      {stage4_8[4]},
      {stage5_8[1]}
   );
   gpc1_1 gpc703 (
      {stage4_9[3]},
      {stage5_9[1]}
   );
   gpc1_1 gpc704 (
      {stage4_12[1]},
      {stage5_12[1]}
   );
   gpc1_1 gpc705 (
      {stage4_14[2]},
      {stage5_14[1]}
   );
   gpc1_1 gpc706 (
      {stage4_18[3]},
      {stage5_18[1]}
   );
   gpc1_1 gpc707 (
      {stage4_19[1]},
      {stage5_19[1]}
   );
   gpc1_1 gpc708 (
      {stage4_34[0]},
      {stage5_34[1]}
   );
   gpc1_1 gpc709 (
      {stage4_35[0]},
      {stage5_35[0]}
   );
   gpc1_1 gpc710 (
      {stage4_35[1]},
      {stage5_35[1]}
   );
   gpc1_1 gpc711 (
      {stage4_36[0]},
      {stage5_36[0]}
   );
   gpc1_1 gpc712 (
      {stage4_36[1]},
      {stage5_36[1]}
   );
   gpc1_1 gpc713 (
      {stage4_37[0]},
      {stage5_37[0]}
   );
endmodule

module testbench();
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    reg [53:0] src16;
    reg [53:0] src17;
    reg [53:0] src18;
    reg [53:0] src19;
    reg [53:0] src20;
    reg [53:0] src21;
    reg [53:0] src22;
    reg [53:0] src23;
    reg [53:0] src24;
    reg [53:0] src25;
    reg [53:0] src26;
    reg [53:0] src27;
    reg [53:0] src28;
    reg [53:0] src29;
    reg [53:0] src30;
    reg [53:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [37:0] srcsum;
    wire [37:0] dstsum;
    wire test;
    compressor_CLA54_32 compressor_CLA54_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h9122c691b3a4db9e93e9f3480090d3ec609364c782910caf8b8cf4b378cc89329979254146cdd023e8c3d93d96f0c65a2b5358018b0b25babebe1bd5e660b9e8fb86ae25d11ccb843e3c36e8a9f6f6bccb7a9368d5416676c809dfc435d54b074f3ed99db2b34fc26a70de33274006baad286d5b0369b437fef88501c58543fbbfbe92dc14e239ee61ebef0c46bd728b4e1571c32520f5fd7e838c7ff21540766385deb9ae39db23eb7d5c9b02f932d7fbb3fce3b42a72a18ab94cd13970ec013ea1a38748eea7fe40e4d895be1f9d3c14a805f9565f7a4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'haca671c2e64ced66c289435c7f6397e8c994639191797e89f11bc9673edc7f2940d8bc7d8dcf3cdd67ab0c28f1e32edda2737a851f2db34fa9ea361e1f7572fdba4d408a6e19caf2090cf5ab7d6dae890d23a4c0479ddd581217225147e79ddbe7ffa3dca3d7dbfc86b4df86624b38f5d3d9e3bbf63bf602e36dcf331237a15e508653dc722a7f2bb632753ea32b9f6a0aba74d19d65d2cfc0d42b2da3f1244821eaea0c2a57bb007d1ae385c992bc6b5f368709165265b34982798de04782edfc2c8c588fceed15b3cadce970a436927269f52e22247ab4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'he67d39a069b9025889557ee0286836d1aa66722b44d01cbcb2edd35af69a868486a3837fd9873c23048036d4bb682e255dc59e52b7b4750227b0eb110a9785a8bce7b75b94857ee796832dc287064ee5e4b9507d0dbbc710462f96abc557cd9fc7454990b44b29ecb3fbdfefefe3c7a0aff96da5e04bf2f93d07449a28200cf7b6936adf514cab993458c70711d8bb3d1fa039228743a63e2479cb14b15f8b72e0027d2cd59bcc38d22c4617a6d3a6c348d69aad6092a0647248b7a8d1c8585ea56da8dd2296318bebae9ec3afec36e33a669d6f4dfa64c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd38a0b11ef073b7695222f11fd3069fda50a748b09480e64f8eef8613eea5de6278c9e687b2a9509f28030b7a2734dbc0b05d73b42036f69019e669d612d333d52012d5d51d2b2b2bc2ad96b09ea5d3224909e97f309607484aa94e6d846f4cb2373ab13a30cd51b3c599a5906b55d9375ee16c9e96aa4e9b6910daf1f2643efa3059f349fb94e03c9e3f44aa94562456d4549d196d8291291ddfa9db0340dfaa3acf482b32b2af05d183ba9d82c599e47b02aff054adec6bb19eb4c385114e35dc3daf4b56c6b10665eb9da9dd83c3de4dda36b029cddb8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h714fa3084defe5bdc70badb9f55bc38c8662f5f56733075438d3f0a856a7006fec883d55220515dbd99dc5b67cde211bf237034635719ba69347d23a298d724a47c03975e4bfa671e7ee74f437e9d533ec32be0dd773087724509f05d188714201f7250c636793361a2f07072ca16aeeb572e798aa033e1c66da3b1ec92d558d462be9b38c3a994bfe359466423caa5a823faa5a7a19f6cc21deeebfe8fec31e3acb1313077f0697380e4f82773f2e09de8c2864dc8f10cd9b12decb78e476a4882fd4ec2052c6af32dafa133b0a6b96c2f667ac0154eac0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hde585faca937dde3a6189919a889aed7ec478e6b86bb744de7bf50a61c0bd7ab8fa959c6661a70bd980ae454f702bfe74b2030d467bb78b39afbaa55940858b67e511a3021a140deb5b10b7d7db8bcb4c4f78a1a8b131b23c6b7057e2fac822aa2b77a97518fb7e4930a24872e99c471a1e94b13ac7320efc3e4b235100e90b8e2d217b4e8c86c5035edcd07f5028258938a4153795cbb740e88ecdecc15cabee891447611d82049e330f52594763bc5a5722c597aac01ab7f6c388c4230ebb73e8936d85d921d2ee06a0ab9c01951f0d5c657d2f1033649;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hbbee86c9e96971b772248bcd7c1b2c27a44504b6d78aa51590940a4f24889f3bc5b64f9f00b1f609952b4e5c3bd166d9c0db0be6b66736c60bd7d89dff17bcb3ed8b46e678767a75449bc8bbaf905e35fd317e5377488a3a5cecf7fd075f2a2e14b1b737febe8b7b0cc2c8c4b7f044464d63e2e4b61e4932b4fe95b3d861e03fd4a6ae45758d27c6fa2e3f06a565f3c4a5be458ed796468dd4588d9c02c37b597d7cf3e8b86da91800cbb6bf75e7fe9f1e5f30e1d9f46ea282199dd1f7acbfdb13c73736e432141eaea2d4e5bef2f2dd5e5f05a6fce4fe18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h7134094ca68a64ef7a4f90743d50cc02e9afa50aa9c78fa1c791a429d9250e5820464e8b976e24ff5bd32aec34bbd6821df22e750f2d6152d075a28222a58541e104f339185e5a230be562f22aa33d30ce5a107d1cadbe9fa9f27c6524decc304af90aaf09c247ef62a5fddbf27f1ce452930fcc2e27c549149af6bdb43ccd52bf71e5a21769ee23d70ff319165672708f87f392abfa2062e8a0484d7533dd7c634e980b2df43e570c2c8a3f30e188dc96c0211f3532a444884f7c21137cba115e1870c61d533f4e36e14d0324e557c7e9dad6236feb15de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8473bf0643e71688af64d07850b504ed74e336a8b0b6bafb31e7fd16c1c7cf842296382c672de3c80e374688a498d7f2fe361307a1febd6779692f862d09c6b9550c78ca5e6e837f968437e1e14023a5a35769b4e0670c6d59cfc5cee9f90285c2325f4be6536947869890678401665fe0d863da7ad946f38e776a3714929a5fdd43c31d23d0bf7baaca5d66ea39a7777fb5a91b584481f4c5a8eca4d4d8f656118cd60cded9e31f54f687f9ea6209e7ba7997d6cb98f35ead6c47153234a752f0c729e2080b2aa5cf78cf0eddd9c34c3ec4f577614f525f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hadbf6ae70a992fce0a6af16dbde4d9b8966c4dd9790dfddb5e093ba5cd15d5fc69c56fae90f20a50d8aaefebf442f75c27b3529a1f22ffefba3fe805c47112f290309cebc0153de19c7cc3d891cd3e2f81ca84abea8bb42a9973030a34faf807d7422872db47e2493ad7d8c59ed8d3f6b8ea6157ac8630e920b429eccc44b570289bf934182e4e5b7e94621b8d83dff82d7752fef9972b42ac2988c296245f2215894c2195f66e6071d8799d0dbc47c50c7e77ad8d9cfb57e3fd1caf83f6c2be38eca7b2b7c74fbf9e8ea0231d44ec154c3695d1e6c5cd9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hf63781544b8600d485b6e5451dad54a96fb9ceb059b40ccbdce8b1954ec6975215246050430f4998faad9fbc5efbf800e3112d805fefb74d1d0b90252cb747738c76c8ab6363471996d0d86841f2db82990884acda872c4e5c37e91f207149f27e1c7155c9ed025618a1b4a0853ff015361ee96d5fe045a7470d41e849f6b846f164793c3052ef62ada0f31e9f813b5d4b7bc068e145d1ab177af876abc4984dba78004bd193c6644d73286b542c77066d2dc4002bdfb8c5851901f97e2ab21db8093baac3fc6f1c0aeb8559b9acc3ff836e5ea64a9b6983;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h75ad50a009e886ccb7ed36df8960724df16fb3a5900637658a6f2615c8967fcb004ac035ce9ed29175e6967581ef332374078561cf02c31458af41741881df7bc442987b472fa79a94576da2dd1337df870c006ece742b86332478124fb8e6112c3898514780950bc4a307520fc90740fbd0ac19203b6fb712314d94bd77b595e77f2831f4c499b5d3103109a72a014b076c1ab608d3bf928927467aa98b40c6f5b06d4a92e9a47dc636f7f274c4aaad5b1c2956babe537c706b4f3941ee6b631ce792d9ddd997a9440a6b69705c417b09ed03983c32376c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h638a28123da9cd710f62be8677459d949c6877ef0ec1d36934611eb1b541eb1bf250d6cbcd9b3dbb1cc0f63fd55124b73d574566f319669f599fbdef2ad81679d489a279be637e78c58cc7fa2121fb016edadf3066cf6cd5f0eecf87c80a851afeb8d609d1d29aaeadfdbe214517d7a8b4864889fcc497f9bb454ebf41207cfc8107565742ca949555a14c30f4f268aff57424aea44e194a49b615171dc7c6ac4b91435a98808ae586d2165d030d9bb06c0cf34539efa256275fa27a4b05cb007ca59ba51043ae5a09888baa67e778f902d2725067d223d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hbe4a7401479fa26b7b5fb63f3e501aa355688f5dd082b77f04a99224d7658f615d9b36f162587e7812d185e9c5009e021eaefead960f6b6835a219942600a5331da04789c292836466ca83fac9075ef32450da7f244e5fc17ef57f6209fed2fd09e144d13283248663a18e127c911a0a81157a145a1b6c11bd68027c013fbb23e465c099f0dffc437fbc2adb97390ce11bb7b1815ec5b31bd413f254f41e544324d1fd9230b0962e20e63809638a0a467814666ef3ca69c88406bfee0145d084884a7b4d404bc928acf23a6b6d3099dfc4601704a2764572;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h11dbe687de602b620ccfccce83d46930a8dce09cb10bdefa475540f3e53d9761291a541a3c1d2dcf07b42d6fbe08cf04cad7c8a2109b7358cd3cffcb6e9d3945eaefdcc6dc7f2c1ee6b44314190741e7bf17a9dc0c9b799ac5f3c5e3a43341ec0c7cd879296dd927c0d79c912082190a4434c454fb6d872d85e3933ee9434194c565670464b6bcd99b16da8a365cb4839f951d1421a8596a06fb9e0169821db37b58fa3bb92ad16cc33f707806470480abb0cc6bea9a2edff2952d546e5a62040a44d3bc0b230b459ff15096918e52418e7dcb3fe0f71163;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h2cb5ea83f547c3c6ea97aba49f1fbcfdd490f0b5c4ed40e22312691b10f3949b498c9d288f6b2797209aeaac2fbe65c8b7c231eda90d9c61b67e4ab8c0ad052a5d3f9f5f0352aa85d573164e799bc6d7719e33f30ebb1f6b3730213102790f9e7e07e6237ecac81f6c8bd6c4b3180e5c209c2fdd6d72092580de12361816046c076bcf38d8dc2d7668167cbc06c9c217eac44f255adfcf3630322eb1930cd157c6c346a6cb04b297434fa1a0b71d1c1557c272fca9520fb2d2d278da83b8ae6cf04e7c59a351b4fd1f9bd5afc28fb4a9f20de04b7ca61589;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hfb68b3412256ae76fb15538740896fb57119a4f940228cc9f84329db766ab263894641007610ce217797af918dc0bdba3d8fbd9d5a31951c2b5d785050fcf3f8219362b0d83395cd52a59307c85bd54ea6b8be881c6d2b65bd3b4ce42349a7fc660114c6427c66b41643918b6099824b624cf93c988865738f797079f1cdd444a3060365179cd5e809db219b83e53328f7d612988e598f7660f2aea0a660d639fc9d37395552a63a74d647c5bec9cd8f5d532ecdea6d38b2fa71ff0d788d49d873d0e2804dabb8eacd89c05c96eb701061df0d39848da38b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd7baa543a2838e89e970b405a502a80e389b765073f610021bbc27173662c63bba097a1bda6ff4ab4ef8101ee3f9f583e874ca12c85895825c1b8c728223cb8cb8062fcec41e8199b3be5fec8c265d1d12336da26913ef1ef3d7894fcd69c747bfd299d7beb0133a54eef0fd21e18ca79c7e1c19bf2f4de63b2eb211b5bbed9cfb2bd33103796c6d5d6e034ac3d1b15b27dc7e9b499b770c365185fe536097c6899ff51ea6cfed03407ae71b696f98472a07e5d4404e0cf485a691aef294947f148a24683857167c2e98b8b6efa3a1f0e1ea59c20d14a16f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hfc76337451be019fcf464cacc6597371133e6fef98e126b6163162429581f1212c62550b7b2dbcc8a531a92df247ede6dc5947f3edd32f0e074864a0606bdd2837c308b24b3bc281d6032d401aaa143248c2220d314f640279261ecfc1c4a42d87f319ae319a7eb50db17b97edc9ddfc3632870103b7cd343ff1ea6fb522ef8ce23deb3057160be1b1c4ac04a262b74badfb2e738e53dede58e88b939f2e8d5409b7d9158539ff0f46ac01fa703638e817c139d11b5e2abc5584c16ac72f529a0eb922dfb4ca74cf8ce52b1005ffbc70ad95f12286c1f21f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h12a96e44c3f84825d09ff1e83c1208f9484a55c48791357d2fa57ac1ed3a451ae46b9aeb8a027f7b8193a5575bfa23fb7c8220a3f78a3430eda7f13a1d031fa5f4885d5e74f2e6ee893c173ab2d768657c0addd7bcead08ac704cd1037e12e1250f81248a5f90b115e11267f2cad983072b5e5bf3c029709675131761955376bf457fc06e20ace20e512de6eb9738de3fce461101ceb657f86db7c63ebda08e30920b5f56f4263b067d9be2461bac8c9115372200464d46b3bce2cfed6752791dcbf933743d317868965ebba6855be2ca5e8d283b74cad5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h6caa6b12e37c684bac56cdf2515c9aa25fbfcba274befcad236a8687d86460f239d3eed79623ec12e220058f2b273f99ae35c87bbb9e6e6fae73ca273686279d37f625fa69a8691fa4760318108c55c6fded3544ef42966d2f9963d7976195574358235f9a4adc484cff091b3df592ae85453ae52377b22a014f72940deb2826f4c42605ad98c62f361570381b63c3372fb063e8ec4c512a5aa0577df12b781705d23538e438ef5a66aab6e7c93cfa0f745d7f4a5193cb8afce0fe574f684bc5305190aee4f48acecb313cf3ee16524a72beca288d948bd2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h9f550057ea3eab3be976120fd00aaf61bdd3830587458ee8a7877566b6013eedc92edd25a386aebded7f32d832d9c25a09abd1ca86ee774fddcf1d0c90ba2a8f1e96ac2b44a66289ac2083a4f9df9c6dee71b7017ca82c3d591a07e4682f64dc902ae27808437df4da8cd0c7b9c4843b8f967bc1a918666a2123773582b60225617bc5990ef80a388db78c22d3513a2b9f6f8343598fe71799ab4ede81e4a7c8b24e3a33f28f42b5d09b1016423f7d73f2e166e8f755bd20495c140457b643ebf5963792160fcb6e0b77ecaf60c00aa750d2fbe23b7966b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h638aa9c154d16313cf6704eef9081ed9d4984d8a5047ed8e486e165bc8c0a501d89253822a08e97d1f2e51bf08112e7de79e89657f1ee6d098385cab03236b010942c3a39d8e449591c4a9b2b6279b5d388aa10ff06c2d8d4b8a8c192e82f7ca37a355507dadd289d082024995e057c47bd98ce175bd0c6f364c1da0ade74468a5d640e8b633a0ded669eeb536d255945b830bceaa94b7aa03784232a25931b7f442f47537da4873be36a5dae95e940e8c7effd4a42ad8b1c7f29ccca9ed18924de62df619270f1aa46ff936a869e11c1982bbe6105cb4b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hfc9ea22fc371b89bb764e88d7f853b5b7e282343863c112c6f852bc84df0f3cc15146ad3de3696fd97a44f619a304e9db25c3eb7487765e26904c3561cf236dfef02bba7f3295d9e462f4a69b3818fe48bef5d19f249876f06c0af6ff9370fb9d8d7a3c5cf5b107eac11131dcf0e7f9bb9934a3f18e6c3311d8f5c31093a0ed94829473462482d9c14b3cc3a6745129e1d73aac20d2d3464d4a417e388642294b3b6b0c380ea6681f00292c2d3640944cfe7d44223c04014bbe94511aeff3842e825288a4b973161e59129ee07db90a58963f788e36a1dfc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd5b28278b173b0f056639748ee5c97b3f10b6511ddb4e85f9477107be7898ff9f241559340400638b10df1b97b3d275848a8296f550c58d001303f71d721fa80ae4c85b4e45994ba16556685a6a139d28263e0edb2c7a276dfd27af61d0fe238d445d37cd25a10da9ecae2e854c1951ad18c04de928694ecbc96dc589aec0892d805cf130abf2c8a16c559f0108187daa4b55904e5ad523e36bc7692c3d6a9a2f558b240710e8afb060bf8355f5167b9bf1eb93a9854ff4c48fc26fcc9e87f01e40abd00d28d95f648c5a0fbff839bd8f01c0704f8716a67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h5ffbddf952429089988a8f3085f0c1ef0a46d64b70434381d8cdb3484b1e81efb05d43f986dd219bfaba08fc55a25106291fb111fb79e6b5049ed0966353d026c0fdef21d7773d5044323604695609e442f33d22a7d9401a81fe51d9bf967b263d9df57fd4e4f8d37784a91129437f5244ea806f512c51fef921527dda7fe3fc3f0937ef4d374ebeed179a7d690392d093c4951ac185eb4b6aeae8d47050a76daa622d1f3fef626483bc0028cd51ffd505b0c7832d2bf1b3f32414d53f2720a332ad6d0ee190763d7d8a796d5fb3221e8977d56cf64484dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'heba1cff900992a59b08a5f459af3201a6ccc7d710ccffdb07d8c4108e2fb928c34503db7784cbafbbc7db3c0604cf5b90642f8ffcdb399c667c26dcfbd3fcd77df1ef46d8f4c5e836dcbe09ff51b7b1bd942edf4a2c9b05bc1313298eb9fc23db6f5833875b6d83f11bd34793cd234c51c729798a15e89e6ee3078209164e25b23d4745d5467dae9a7b61827442af7eab82bfa86f19f3855c6a409ffdc0d3eed784c75e0b11dddbbaf80c4c498f614ef2dc52332e2ee7c2c895f938f2749eca3d3f2ab25f533c5cebe3ff7cd6cbef6b1037f13f157c754a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h7181581e18281ca97ec27f07ee9a0a9763fb7d8f7390a7890d8a925d7fd9ee3efdf3bb19340c3f4ea78f5b12fdfac0bdddc901f6d4dce953f3791620b69f73b525408fb28eb7532d99fc8b8ba8b576c51f910324ef897e717bcb938a8667d41671cacb4cbccaa3b0a577215917d846f9dbd0c97245a55f37f673b6484f3baf474f100222bf74da04492cb5cf0ad5b3ee9ada13c0266563cdbe147ec1168d40328abdf9b86ce4853f9dfe90ba61d511dd3f08a29ba25df27866611bc9960a7604b188d18b1fe6f30beec3b809c75a51b7d8fb31e89356e5ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hafb6aee4444445dc322b327025f152655236d61714330da6a20670b692026b40b41513ca5520de08b8eeca7d1fece873a32c1fa3c4111a1bca852ac38b9e1421485e17ca276ed7d36371c76885b5bada31d66101184ba6defa39b3802ae2d0464f93b66ce48fb72b52da37e016d69090f35caedf3f8dea752895cf8888a7202e24c6731e192da5cfc8f560e1ba0c8a1fef2e70e79e9894f8726e4cdb6d1632bb627663ab570b81e899705a593dc651db05af45a19ab8b0f03d08bb3f33760908297dcec67d94c80650ca05a3435290819b1db082c260a3af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hef0e448005b9a14f71ceaaa3e1562434a56b865ff3f3f520ce4c2fc129df879ca72173bc9b90022b7ad63041bb9722c5bb9544d8b6a720cfb7805216f7cbb16868ae96b302938f0f6f47b88587e536f1f86ff14666f65d7607f932914726a8b1f8bf9fcce3491ff475d7b8d157e2ec09e9ac31befd66ea22d6edb808a44134cd032274aa055dd6cdcd285c5e5c6b76645c97f64b8867ef4280c7f675d13173cf02a1f154339d8668e4cf78be7b1701eebae2e4fe7b4083e4659e740d28ed750bdfed5780c6c218215deaa723fc483eda95fac14972a9aa4b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h5af445372dfe29cf3a92885c92cf1adb56abf5b98ed9537c7c96540984434cbea5b88883e4464a4daa187c6fd5410dac44e6d6373448dbb8b4fb88d2bd0cc002379b0c8b6e6363cf780a3a49830d755afc0e582bc97e6ca9a7e866a867cbcea7dcdf558e449ce7020204816f86fcb6aefe211600bef78426cb36963cc29c20679959b4b02262f6ca9a446e90e637c5caa4b478b786e6c7d5cb1e486d264f542284cad477f67e15d44dfeb432aca6ee095ebbd2d29b65ecbb2e02136fb0c3517b79bffb367020e22e9cdb67275a1e196a3cc2fc0a4b2840f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h5fc4575ce590a034d165c68dfba7659f6e28a06792e50ed2e939b105584cb1e1d16dd5598c3b8b393f0f0c0a093287c1bd9727b8e44a84adf7ea68699ecc6271b5f0f443dcf77228de902d01254a41386a97f445fd3dab80bb997713d299798e71bbe5d7b605fcf54025dfcb0423101e7c2b2cd0680cccebf5249221aa1758e6cb13fe4f105f6bc90d95cbfa39a28c8c55671ca534ee96a44da9baf0082fcc12b81e2f1b9dca0b61c5e438a8501b9898cd54255f583dd933ba41236bd17d372733f8875b0f212293abb0383e19d5936d1dc86f06da4a6a3f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8ca34c296801b072dcbc2115a94e18b6d1d7bdfc21d8642aec12da6d0abecca29790f0468bc93af3d385fff71214671e53c45ef1df2db0a2b2a0e124f7f50ea1911db590c410fcb81042cf05940bc6be3087c9da94d75b1f704efb8eba11593cd8ea506f0e67f8c05a27e33317669aa0e18d43179b0be2daea75cb42c08a10c10b2cc2d0901b812c475ff8bc6a0cf07bb429972ef29675a279c1aa3b2a9bc624a47c13cb2bcfee19c74fa65f5d6d31bd97d52ae99889b7d463c7bb40d30a6bd08ec6f8349f5b6d9f5abd4a864ab9790b0576311ebc27133e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hf9e73041106603784fd1d10dbd43105ad38bf9fc0800d2f016b835f2f0473216b1e25a10e96ad4bf3fff77e4c68ec4ea156dd63a4084139d0536fb4e89f06874cd2cdb4605250ad3450c1446e910b38547304b59a6692b87398affdfb348a86ca5494994e381e455028a573a2a0dc7a983c0676263e627d0fd96311bc9def075df35de0467d291424f096f01732ff93014935f4f8bcaa965e6104e5aec4ab9dcd8da9056d832a91bf8e43bfa18957156010c8001b984a1e6698f0f3d603a07644b29bce87e0f91a3fa4f0f82b76bc00f3101ba193d306f00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h17d5f183fcf54eee3d228179a65f32e1722cc85569ac28171f2d9631dc4da9bc0c85f5d23116fa32c43749f2d133417300ddd307e8484683eca21ab1096b7cdf4cb6c29992a43d58e5383d46af0a945c0838a6e688a2e547a34b6970d72469aef8a04de87ca935a119de131e6501e5aaf1a07acb53a9076a0489632fe36f822d17bc0c78dfac05c7f2d5877e7762eca64ab34045df3212a1d0a4e7a6b42eb75f52119704077310f8e2e31a290db6afc2082d7bc5261f0f0f0b68a6fcb58b42d1956fdcdd7d516ff1df6c9b1b70e8e5a75fb6cda0568943c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hc9169803fb038eda43dd873fdda4747b6553fbe784078ad78e45d89311f2b6114d1e01b97dc2f55c368e702c393bfd652c14fa3ff0eba40fa3b98c5c61b93a024d7515f62591fa2a9a116241bd7ebcf9ac0f1fc144d7b420596b7231c7f3729972db40f34fb011d3eb6667e1aca9d904feabc6b0fba40f9228ee98502edbac84c1ba3af3602d963dd731ef7ff9905c956f9e129e44628ca45428d018d834f5987adf78a17f8cf47db58445865be8e449b8d7063b4f2efe783cd96fbb6238a02999b61096cf6301bff5754323f5c067fe9c850c555fb9a775;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h88e0a1e1e330dc01dc77cb347be91dfff90dfe3b90527de62ab8b4fff10fc188ec190a7580771f2aef541478e8308db8d79ffcb7c103101afe56fedc3728b053560c2e51b3b2f4bbd81fec3e53a60eec6a6aa04b2de40e03f93f88fef60624a2cd6d5a29227d6b6150edeb82846d6da64fb3db78b513699e30c9b9d5e2956a4aa00f72e7ab5383408feade49873c3e025210d2a4157266fec8bf7af24441f939019e6190fd0b52358f3e19d84687b259ad5e3b4e602012f882629a4cad6384000f6655524071b44e3093953871b987f6c803da69180bc5fc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd6ac243209b9a5185f1706c626063230416a10f183511a6814a579b06cdfc92d65ffcbcf104fb6dd9e40bcd3a89aea4c420af7d8100909894a94153858bd84d6bc073dce102895f3d00bbce2071dcfa4370f336fcccb64e0155caa7f060728476d377d3953f684bd7213f0afae93c015b12b379f6b2c3e512541d163d2cf7b2c7c73a44e02cd6eb65de28f9aa76dc04f57c35c65d12879a4cbc9141178ad5a3effd41e3d30019ba15820d2b0d6c0effe7bbeb01068da8d57626d8a7f5dee020ce1d34cc18440799724134a86e1c3951dc07581ded6bdc1de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3c7bffadb66e212421254380f8a1bf4da575d638c8c4e674e23aa262730e15ead1c910fc73755c71581832deecb59c86487ea90a85dbe74b4872c0298421e3731d17674d0473bbff410fd4b42e22603e9a6ce0de9075c0f1418b8dfbfc21b489edff94a4f7d3a8db979f3e34356b702861978df1c30b6666219d80e77d6ec23e3fd0119a664bff1afb8366dcf3b06585cb8751cb1e2e22de79182828883b3e983bbd4242e4237d2ccd0bb89c583db50a5b17e9419d435b6dddbbad346313b2b0b383fad5f0530db52fd612f73e330efe661ca1dca53bff99;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hb138326f909d57448377b0e7306537b92b20eb04d7ed4195482531aed5455c7b0f7effeb8e99414ef84b4acc56cfd47a98224df104339fc77f9a53513a666b20745fb8c38d96be185a249c941934f5bae675cfa15b747f9feaa1163f56b0db886cd2b497fa5817d474a3504b0d0505f5ce506cfe1673f36a32154ca5b7cd7c4f3af61d10b29d1226b765e3bca80f6e5ef447f11cca0bc93a1fb645bef20e94048d05379841109df8400e316cdb84ccdcfaf5f33633ce7eeee3ae2edc84d4d59ca2604f482e3414cfb572c1e800a07c5bfa793a3e1b29c2ac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h626fd62b63cb176197b75f229a820a446857fa3b1e60948e5606687d2b6300005b840b9159d3fa40930ae4df86eac1df771250b331aaf5dd964de3827d0da6d71aee44f3d58bb5ba029621ef047c6705be436e403d225aaee334f3c640838e2c64cd9d0c9862d3e8735ce367fcc4da8c3a5b42e6fd4abad1755824745b62866a592f587b5be96e250c89eda5b5f1094d38364ae05938b8a2452af325df7010de1f27d937950ebb4c653b769e8ac5748f69a10649a7e3bf3e5e8cf23e9e8fae34cc13996c4f41cce5ec904ea8ef0c175cdb45b2ccb5772875;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'he5ebb6e1aba7b2b726638e65405b78e7ff2473fe36e3d1345a24ac0cb8cfde279b959b7bbcbd896e48f6ee5832d72338b4ffa506e95a72307ba00a2cc9048a39eafe5745909f20c3b662313f3f5df3a1b7c91aeddd39859030dc91c45acac0996725d96fdc2d560d75fbfc06300d5d66b4fe4752229cffc5a684fb2a085ba2c1c1762b6a685d487d1e9bff94eaff05727d52d5d0ca9dbbe9d1518a7b97e33ecc6f1b6b7079eea208ad56dc05d7b4b174f183db73bf62f0ea195dcf4dca7c5fa349106184463d7a2fc4f65ce48b17f7250106821607591a2f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3fb24a638d7f14a81a8162bb156b4b43060b63402194937f818a7d93f0b55dd9eb535214ebd28850b2158509c6412dc8ca0a4d749b6c62c5a24073605159aeeef99f02b550ef104d97612ccc2759df01707351349134f40adba5be010d8c587579db037e6e4ae641d235dbc9cd4d19919c2869e7554288ebae3cbb2de1e58b29123c79f670577aa411ca36e35dd8cf8ad79a629b74d859c56958450499155d108bcdcf2cd942d425476ce7b15b3b286e40491f595564541480d7c016ef8bd563868e4981184efe7c79854fc367d0e5aed2dcc0a4ed729bdf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd580f3284794371fc892f3514772611c15b004f07076c9b0e54e5c9b76cb4762ee76d146ebe1a8449321b4b6117e766d004dde7af59fec652ee2f4c012edeb3077e764cf20bb8a7407390907504a34eaf162458273a31a0bd4eb8d54a8443ba1bd03d36e46d5e8bbcdae2aa504edfd1d4d8fa89ae709663de56dc88040a92aedb9d39db53de1efec40bd01969bbfe0f69a5f73b64683eec4fe3afec8053ea13c191bd9a2faa84164b6dfc4bd69c33162cdda5bbe9c9891503223c2359670a185c6b9f7458c7a8c4503aeb8f44aad44453bb498ce8fb9196;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h9a98271c449c5ddcac4abae17ff5d250d2e16e2288f6e690c6c76abe282e15da14ca61fb54bf52ee5b9565a68e9dec48ed4b45955bb89e18967960062456cbb42282588d4bce4ddc6b5df50bdfb6497567c5f3938173ee7b8fec206cbaa395d41bac098520d125133c7fcfabc6a81f75d74d1ebdb377dcfd13cc07e8ae9ffe9de0b4cd6b1cd3e812e4467134928129792c5cf3923837209609b448bf47e0d136837da2e50a803939370daeced60b10567bc58e7ff5497a8686e1086da8fc763b05bcd4de37e1a6c182e097ef1eeded8eb56eb29daf3a66cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd6efec331a1282ed4b3bc70d45d59e48e5e7c31fcc71c1b5cb4a081d6853271bfa1926effb96a3a164b82733e2816f6474eaf72484734a58e7a47fd682c51e98b90c5c92d93cb3d532cf5015805583ffddad61177dbf5698ae244489512a91905739458ae63d4565a21c84ded9232db0eae8e95568b2a33c7a5c211c71f3f7fb27ad4d6395e76e41d03d5cbd9dc9d63fd61baa55f353b5086c50bc4baaea0785d3f80826966579580ff7cbf6cb4115424152292f18bb2856d000c395c59e57a2d4da15549b47add3fccd51c493c6943a1913cf53fe2e037b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h1324541ff281495ccba166374ea0dc05e4b7e97b8c21c13731afb4e5bae5522fdfa8371184d08c71c58dea5b622e88e29a687e6fb1ba3ae0f89d2717c836f8107ccfe97f343abdabe007b7d4a07d29dfb7df0d0463011909af7e010f3bb71e76ca8996075f58092dea3ced0b33d020158eb33b5b94d9eb2764d8229ba9e6a45ffa77c4f2b0cc3212f573d4db57caadd61903140c801f839739a3d7e824fd0d66a3b2a2f5d6324b0fb9cbbe132daef843b53956dcc20eef351c4919899759cd72454f1aa219918c31d316c5fb0b6acfe565a068281416a4ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hc2528d88e8c611289e73644de8e16daad0ee5826906ec1acbdd5f77f786e2d02ef808216a28cae47cc8268faa868a7d2daac82f308967a371b1945f3747e5d9e4361c802c2fd102db38fb1afb0b31058e8226dc0763ecd922468642448dc65e072bf247508504f2b942d190633c8b493d84956e71fc337f56115520dccf87a00c7c020b1d024d4bdb4300d46b92d3be27b2a877b33457911391dde2ce7937bbb0585d27bc665ad5186e1c1a767e2fb9ed274b3b11a60df8bffbf4742a484e5b589caa626ba67afb7eb3c3e8057ec88f39d7644c49bb36bb5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h229e5d7a7271d90fa1a9eb3bc56467b7f21dda29613d965689bf60c7e69a955b5f70a6307af540395343ff070413be17f2de79eac3e7c8275f65e3fa326a4c25a02cdda4fdf50f9fa559ed7cb028ef576657a9a3440cad5dfae206dcad4aa39e41a7816a2e47a6eb7603fb0c7dfc2537b7638c95ff2090d7ab548f522c99f30b8dd114fee71301fb1ab6b0f7e1c40af5d39a22cddb0c6958b184b5065a6e6244abe7dc0b9bcd71e287da1ff1d78b3a59016047c7a33b8b6f6e744925573ede8d6802d0fab6631a1fbcdd892e5a395d927a9aeae5a6186150;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h425874280dfda1c5531c7f92f54f7d13346411939fc5c65e529ce7cbceb55a827dc492aa4ecd1c8f9818caa3191bbe534d094a7b0f91f231751de67981f2f35186e38e74bb4611eec66501a4294770983d74a6d5e2f809ac7286347026e4cf3443d03c4526e72a5bef973296b6b1db0cdd7ae35d2b4fbc60d48f667b6044a4ef169e6993fa4be09bca964547d831655bfae8b455a219d6a4ad8e97876acd0ac995d02534a17a9a7d518136784c4809cafc7c3e4a21d4b238f2087dd34403ca2e77c5f4bc81921ba22e71bd789b29140bce309824e177e655;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hc79e1f33696e530f862d49f4a6a0e75ceb0ac20ca29e8bb751f01361541c94f5d183dba8c9bec2aa5b3a385e50bfc5282355c88c9812b18932eb8b21b12534e2c0c41cce222aa8dcdbd0b2987a1a500a6210982cfe8dd672d8c7aba3167cfd4dbe7a2ff50d1069012add5a5b38b8eaccd6b2fafccded602f2ace94d67bd9e76afe9ac081003c74558004f41f51860b40861b4aba321953b25a79643c4463573a3c765b5db3c38c8ffadbe89c7068e4cd448084f3cf82eb551c7fe01538ff3a3f203d45674a7c27aeb3adbce65946c30c6865556d695a7228;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h862d714567cfd33980f6e72ef79bdd0aed89781651fa3289c09cdbc1e050bb1366234c415e5a8e0ad3d232be576e6a85d405d2d22f475f7ced8b9aa5db10fbe67e586ba5a38671a60d4d0d9f57536930fbf04b3bb79145f00ba908d51f9da2cb0feb2b0af1f0c3f190719a2cf8ddb84b94dc33800a9a4bb752a6652b23e3521235199ac9cf03dbca0875f7e9a38ea2ea7040cc64d55f99b83aacb3223f3f90ed3fb80b458e802c815f3d6cca4b114077c32304abda14499bad532f5766e8709b16fe5e02041a4a8f583828c8a54eb24a2bffdb41b3ea8b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h1b901e6ab30fa15afc32bdc54094c75f8dd5b337a182a71f05e8defba847588ffea6673f7a4de1ae2a2732c6b93e5079e02f1263bf2c61bf987742736ecedd5ba7cb37164d4f9ea30c7e0128658d426025a37efa104e42cf6d284eae6a00e6f64d3385c3f8a4f4a243421009c2ab171493f2ff04f08a58d0badbbebcca69952a98ff2f8dd84b23244b51999afa1b1d3d628937bffd2d58860be21168e3a134aa8172b506cc522ca719348f26e6683a8fd26def7ea786022f2aff227a1f4aa35765dd9e633e5fe1ffe520314fbc80bb54a58d0a98634e138a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h6722a0a6b573b9249cd26b20989aa7023404079564bce41d4e3274debe5b4cfb42a4f0028e22bad2706d274e4628dbb661aeee09c25d817d503ec0dd47a29b462bc5529bde3ca022de284cc5adee16400bd98de3aaf08623ecd65acdbf67251091f2a8def5dc402a5fd3789e9dc1e900e1a775684b694683a90b9023f098bb9df4da2eb60e473efb85e2085e62f2240887c6ba39c69575ae1d40656075aa59ec24ede31c6adcbff8e4f4cd8dc3fab0a6e8bce3facf9cb2e7c71eec604a641d8eb0f39761ae57eeb03453f0210cea1e6112c119d4f77796f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h559c6a2576fcb935ad8ccd502a8a97ed6a1d9fdb5fea3bfff7cd205b5b78a73ff8373b485e2e48ca2889ddc31de944e25ed896e05a04ae1fe556d3d3ccd92fec24d371754be7a552ddc55fca8a7a0ec6a11dbad05257d4d896eeb73d7877b9d86e60f5a8506b9db8ae3ced6e5bef1cc81f9825e04a5a22645eb3976a870215e04c4077a2dcdbb36145881ea44de5819954c34eee3f7247c2e520c74d790e1a6ce12284307763e2c5533b8023410dfd8ec3a6dfc59d9116d7cdf6bd2fdcc3ffbe5e71066e5a1fc1323e9122370fd780af9309f535bc155879;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hae933ce51f932f4fe86835ccee250ca0aa659a1a3eb1d10d5a95a77c8103345bb40b793d0fc8cecdfcd03bd91f564d5d6adbca86a328f9d481d8906987709803e9176d39d42165c6b78bc424fc75f7ea3278bd0f3c3309dc860d7b2f47adc5db678f182bd4a07ec8eca0d29acb2eb0bf7236d0f4184390d1227b826b03ecd6f279d3eef526c98b6f57b575cc2398b44046637a4bf0c39ad322e79ad92a75d08067513abeb2275da6defb77c598ee0d0316399d29c814f689d5f9a02a35392d230861f144ef162c5e1e856d9d840521b94f1ba812b179574e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hfaa612f19a7f38a5c2652cd2e1ff71360d3a4a60989888a03cd45dcf3c8f7c2dcfbeba22adf84a2466c889cbb38d6eaba46e607fc093e0f36e2dc8bbb29351537dcc966484183ebfb93435ddaa11a99c4e84b52c6bbe9511adb926466dc712e34a374d57b9b525f549d0a1ffec08f9a791de531bff2c78838b0ce7123e60b074a9c7a876743a8c7df4e8c526aca1b4aea291fb41faa10c28222f48a9a05ad69274fbd8533466a4d442e54ba2d8f9f748887b7d3d24830ba27c75b715921368299bee0c492e416b93515f1252fee8f475856e2d10981cdc1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h7a13b778bdead0466273173b88c9da3eede45335cce2ae58907a7942b88b12118b78901835a22e88b22feedb8784cc83e2d214464073bf90fbc681b494dd93c0ab9b88378a7205a337b44b120164c6365544e88a353f94dec58c4ce7a8d1f88c227a964accfc41823a6635c53c3e268da394b9060270f5446a1c2630252f3e8663c0ce95a5411138327809945cdb4abcabdac6ca4d1d69385307540ce6267e0d6b6f6de8d3ac80669416fb47a562a652e521c870711cde70fca71324256fd0741c1d28d1edf7b9e43467c540489a32dad5f1012d8bdfd7c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h57262a57c39133e706a1e3f44d4eb153abc31668393f12b91ce1875376ddf3538796ac490658e66f659f482daeb16af43f3980ad1c61d90852f1c2a204acbd002c08c3482231816c136ea0aeb8b8df1cecb3a0cec5ee6da5e166e7c296a74890c700333ce32335d146df8bc95f41ac45d3bdc043abab3e7d28e169dbfd02b79d9a761ebd2524aadf6f461e762149b500d665671a938618fd0c164d7bb0cb054e0bc2d8cb7ae3966d15faf079682f3fedcd94cb000db55281923dae729257da434199ce54dcdc3a4dedf9f93d427b3ab83c38e76151e19ef0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hba0cfdacac16f51e9a146382339e74134212b63652cfecb37d2f36691a1419d48093a1ecfd8d0c2ed398f77af991b6b14ea5b1f3c00b41d65c7d1a626ebca97894254860858d80fd4e8deb4b079723ce963b5698b9bf349cb5710b85128677640c1e6853492bb0c19ace035e9bc7ec5c2c92a88af987b823c473e9fa3354b6ce38d5ef7445e1ce3dd2b07ae8408f539b6978446fa9ae25923829d121b3e7be6fb51d0c6ff001dfe55c9ad94c389d73b4454ad262a45370be5418bf0b1fcb7178079eb949175621abd73dc64d58a02d5a6dd3bed7e51d229;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h1243268d9883301c28358766e8198fe06760cc348052c593396edce94857ffa3f1a1031f8f20e43cc656d7db1d5eefbe2d1a82f8cb2b9dac406c28fd5b2bb9785282eacddb9c5e85fe2e7800a37d6383aeb12d57559ac75c2cde476f8c56581a4e79a55a421853d901945e63643245de02094e1f614fb8c8678fbfac58d494909a5ee583f7e6c336653f0616401155595d58521122964c45d15272c4b41e6699339061c0ea8a3f13371c0f0b4f8d153923cab72336c97d4d5cce6eded38530181f4126a3fa72283ce7e4821db50a3f0f7cc979fc13e193d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'he635e4e599b20c5c4c133cbb08bb6771253f510173c7153f0206c08456b7a4623ce5b72448fc18794dddd9edb539e239f96644d1626285b931d7c30379c7cbf7089f07782f2b0c0fdc8b8c2c80cae7e3840f3bebc408d5a62730cedd95c65b78912194df1e87135ae4a1df03a987ce9cb815a99772aaa5c73fde27712f1038ac85875b0878c9b0449ad1b1b13dde512f3fe881ba7a5185aee33977d1109a76389e3b9e5a3a7fef2d239590161741ac7e73d3f0e4c0eb0192ec4174596e42cb6979b9614235452b89e7aadfa9c172d7bc1a9f1d28e63c1334;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha3fa98b40acfcaaf65297f6221c0bb57f21554de58633e74ad887c8ae032f800591795114d549a582f2109f514b198f1e28b48312f534cea63490c1d8de91c832cf65faa8c3366625bb05bd0eb44b1c96b2a98f0e2ae9ef66a87e856cca8f1e6da1d1477b2271ec3b03aeb25716201d98a329d857516cdf1c636bd86f9834c9e96e12a93cab36cc043e20bd2a6938b232ba5629dfcb9eba883847ce58d7c03d0f5509545230f8604687e2bac457dca8a96d3d93f09cb400c2194d42b6b591eb097a80565d4711786152b7063ac5986381034765a9104665b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h9ff8f4f7bf724a5c54dcf8ee90d89fb957b3a2c72e76477f6f161b8044b8c89fb797caf9f26fb6b7771665968a126be3b48ba0ac0c8fcf7ea85baa5e6e7cd3f358bdfa6cee619650594a2e13f255e26c8500ccb4ee2ce29dfd3c488d9650d8ddb2b204e1fc05fb10fa4a74c1304b8ad9b7d9dfed929331fd1ce7a1b2dfb261399b1c687cbaffbbac506ebfc21f1e9250c2762cc063807054ee30c8eed839244fb26729cd9398bdcbad654b3ae3e296e1d394deaf1e02a1a1dad610fd09d3eb0742f56754e29c59a6bc623fbfce6fce7e693d5f0fa4fe2c2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hb539dad1bdb703e76cb3aa4d3aaf40aa164c7297ee176cc0e811a4b9f041ea454a42125a3e953dc276e90cd5f38c3bcf1ddc303357e2351f4f6ade64e869481802a4a850f2a82cd8f40e42b02184177fdedf0c97768952eb6cb9e24559f0f54a0348102190ad2aaf5a2a01debcdd79ec14d1007c5c9d56fe60f865750807ecf2736619a8a0a7ddc86eb7712474a63935633445c0f191643b2d44572c7fe03fe4b4d21e2117b86215e73f17b78cfcde55e63c4cb156fc73a6c0ff74638a6162734e713a58ef54ae94c71df5701a295813a813049fc52e9969;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd2badd89512156cac656c3274c75aa62bf61fd130e7a806930934e96dc3894ae4bc2efa9c77fc2fc6f252fbc2a5fd1b50bf64984200f4d7bd60d0fbda9a2713d17eec94f806045fe7070119e1899e8fb0fea0b3c94d34b4ca0ebf8b60425c312b79f752a3321580ee8d78b961024b1d8ffdb5972b97259f33b0a14797343025388b7bbd27222e6cab5243f3b522d7f3caeb5ed1c888e19bac865aeaf5ee8573536f51c6d994472db806e0244e3fc9313d8a6239bd6ab86a7d209ef561a928f2de91f37456e8d2bc2581483990e8a50c8634a21b40831287e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h1dfc0d2736b112dcd435fce901c75ef31aee5659c89e555c3229fd274dba62e05aca1f46c11cd59ffc42d50368c01e59338fdbd5a16831882d6bf0e8ccb9d195d2c2ebc12055eeb73c41b548ca35db22a29b813c43317c7e136e539fce36b1bcc6bc8b64992e93fc441c0fa05aa63ee0ff90dffdf5b6f5b377ada3e75e4a29ff39e8dd39b76da22f041ea7dc620440896c6211a75aafafed342500d57c5f9a36b2cd775e4c5412a5413cd27c04c12e9a574a33f900e0ae4865ecd3bc8f1e96497768a011cccfc0f5c0e61601af0285d6ed9da77ded2f5be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h59962f025587246eae4153610d4eb6640d2499c832b6ada91c9e664c408ba29bef9a1ac897d409cee6fd424e1b7480b648675705c5feeacd0aa6464009482511ac8c4ebed8633f898e236cea4caef9de324a37f5e4b3d36869d3d177b44256e2493ae35f6c4b8111ae0f911d1ef6ec8de655a82f3a677c457841f72146cb1b43f7435b82bb45545456ca04685c0d01d405921f4dd54984f32077969b95fcecb45702a52c61ca116c329b22e7cd3502a5e9d6b9f8d64de98556eb423af7962c84f5552f9b4273a0710244e9e6d11d8630f21d717180eecc17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h737b5eef23905b474f96ce42403afeed17ed979504ad03f5c7dc810cd56fb9e106bf7b24f456020e868da6042d8e2763748f65754d459fe2705cc4080bb571d0315259dbb021d8af8ba13794f8aed69bc2c27305916a467207725bb25885e41720163f12e24e2fa2d9597a45cb674aadc55492b88d5e7acc9a77f7f4e793d8b0b78a156a3a8064ac6f43916b0d7649bd03434b661bf6117314decade29d25dcc6060f313393a217f26767f975b7de6017b5851312dff5e14b7dc1f727db3d2a721b85ba0fb2cd81cb41e2b7fb0b45de39294ca586d22d10b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h635e19661d5e111ee14df4c2a80afacf5a80598da28e7d3ba915999867c013b32a74688615926e51f92fa59891f4cc41bf5211f5c80986e461b8b65cf9a74d82e194562eb0c4f0727e056a9aaf711d87c204ed2364c77c45cc21bd3ce683da5456213b961d3198a11a7dcf0a6eb967fb5a0698bcc2c6ff55399bac8f6ebef010737c2f932b9fcb3ee3ac74c6c95240e5e32991d89c1f1a85916c4e883e952d9c3c4b9933edf58678f466825f9edcd997e51055599ecc5aa02062918edc08b7d3c8bd10d9ccb5b9a909a200bdcd90b88f9811b1c177c9fa2d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h2a5c30d9c283b539cd5937393cbd1e668ca0c84032aef9be445a421b8d4e3f4e4acf780f8201a221610fcf479b41ba51d9bbbbcb71087a3eae85008a5d94956c648b53b0edac34c27e07ba233576247747ecd8182294a4f34dc7e136e624f848c056692de6d851708e106f21f1722963529eb16df7417da004e5ee1a41aa8e716ccfe6a3a5ba1020e6f887f5dc53b381f25925c9afee794ffb983f058f3344905261ad655fc768d3ec4314b5922c7a635c278a5ead441a096175434f6a81af956a4b86e487659c63c0d2b679d198c4876072da77d5590a41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h73d15ed1079a6330b1e88170d8f18433d091efb573be3a84abb8f118bf2187c6c6740bcb5d698b396aa06b9b9d1a550e6cf6d73b53650331378a7c1705f3bb222f8e52f34963d0835d2b33871c8d8b855cafe860cf25ac49ea087a7589ec3b8a6f280980ef7e13f34ce547810c9002a16e4f396777832e08bdeab7da533c8e956e1a2f9d6ba1d896d5729debbfb21dcffbe6159199de529c859309256b4a99fe0224bff35c7ebc2e6553dbf896aa5608da601e656b852ac1e775011c7dbbc3dc9969c59b802d5f0c17a0a2608d9bee32a04e38c756ea5d44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h1b4276311c16acc338341c9e21074a560a79ee34f973ef6c21738dc634161a3385389b4530ae9c939bba5a869b7c0ee357298f282b46214934ed5debabdb0f028b4f0423b7dbcaa11ff7045e0c45f53eb62a85e90a2cbdf949aac2d879afaf961149b0d3823619e3b6c6ca93e22932138838e4cff11a9b2dda0b642c61856e3f35d85ccb3b5945b90a5d2cbfb57b6a3b22b6cf6a597fd71f75f53e37d8ca3263d3d79d6338468477a0208d0d933527270ff94c123b80b71708b837420727aeeedf2f6d042f8a6a0b0f8db80afeff7cf39c8dd8c626d3b521;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h872f19824d45d46ab865a6461b543f63f8b78934ad6655f131119df48ac3f2592570ad75cbb6741365c13f2c4459c25031c92c4a7946300da2d0e38e4f59dbf1d4e52730bb57b9c5ce49ebb446708879c1c3c212fed683766495afb9492c76f1692ec73dcd8e5ba3670cdbdfc5a1348d36ed94dc68a8d8f612171ee2e665ffebf96b803605021aca5585af45f363fa527a3568566a6afeaf4f51e521fd64f933f5c279c9e7ccff56891845d0e1fe6a94dd51db1008ba07533f8a600c31dd5545a54e7f82f6ccb8877d6663f9cb08b632640f165b902c26b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h38c7d63feef76be465d0ffbcfeea3c160cf78fcaa1efd4b5c88fbbf154b50a2a5b767d63857a898d40ff88465c9030cdc2f4c3d093f1e3a7e935a6e6c459992d01885ae680dc7b36142f30fd83619de6bfd5f7446d4e6faed1e3fbb1f8fa42fc2224e014a56491798e59b8d2951db7ae4792be48d06861750dda4ada75da9541369f5da6a60d6dbb9ef1130ed388d6b94e6955c5d91a9928aa26e984234469147ca151a5ae14eadc4e8d2d89e3154846cfaedb78f807e2bd4a45cdb3beafaef9f59e020f5ad126e96111edc53a8aa3c339d2d55b45eec647;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha5a7ab86441ff0eef0a974bb608c708be76cf42c923980aacfb603aea7dbae5d577eaf2402b51a592db34cd12dc6e655ac2aa879001e7aeb852dee7852b6996a43e225e477ab71c7fda0abe309cef5f63854a49fc3c1f60be25095c5d3ab2f1bc0787cd77e45b30f9b5ce69966c9256e19f960b4354b58171bd0e94e3867cbf61126e73fd03f6e6c397e3764f4499d6d9d0a492a36dfee66dbf99fca808fd661ebbd1af446c050226f6f3d1ef020c87eed2985007f3ebd4559df1288e32bdfa5f728e3c78740bae9ef8db15ad2b33805b115723630ae4fe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hd18c70ca7d349b39f4e49cadf75120db33a21e5452cc9fce3e161d19c18815a885ae771d41d3457efadb76ec9868a7f08db16d04377994ddb60a90bdd3f6f4ddc21c88a5b0a1536a8a034985bca3e9d579943ae950b0bde22a06b5f9784d1f9f5d4f0ed9ed77dc0a21e2da6e683ecda7b689167dd5b133fd163fac9e0ca5918fc59e950781ab86ec07dae398c4dbd75a1b8ae82b9d3cc7acde77b46c007fd406bd0c5bdc6bb3b4c06ea9541d7ac22ad6a0af52dc24584b59072cca65ff5793bd15e0bb997bdfefea57ad2946dd1788079e1c7f204ad0424d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h4f4777c933e3052678976457276bc8b67e67cf9d75e6ba2578a621196dc2ad22e8b090163a0c106a7c4c995fc9e7c47651886495e2353825ed66af34279670dcf2b7f91cde5d954542b9721f7d732849ad4a89025e76665c52eaeee70091a2c7b03d2f4909065438f42634c3bd00d1ad74bbac7c04ad436c08523ff7e7af5f5bd4e6e639ebb32e77f331a9cb1350bda9219694dfdc1b8d07eaa044c06a0e1861e12fe8193427fa7c2241af1a8f37aa32a8ffed7b7d44dae09fdb79f3094da5baa9b469961a0e6b5cd1eb9ac278275c920ebd0fa4c6facaa0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hc050df4ff74e3a69470a74da3cb4357f148ce3c029df801ebb67f0b5db77c9404b82defde5da68a5f9d01c52f7a509b5250697e336708b9b1dcd2ac04252ea03ad30e186325f4b89f4e44cfb866c15509d09dd7e0676c43b19ef4e22645f39f016584e853294af9f6fb6caf430f66d5ced2ef21d193bdbc8cd6bf00abc69a29195887649ceffad1f6b81a128bececdaaae471d06639f4086bcc6993b4f7b558413928b2984322e4bc38c126140533f0acd82588cb2b3f1043a1b771aeaa565a44ee502f9192ed94ea87fff9bf84e69011a873c53484d43d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3cb4a9c19bb39f491a66dcf6af5bcc4ca3199497a561378889ada2cd5836b62463a05e94707de5bf403bc3367ee54001df5b403261f3b01416fe47f542a3536f5f3b4fd9b0d9d124a3068222c16a15b0ab6d59138c12c5040952d2b13c214a88298d50931abc26d7a8b48595bb185cb8754b771e649935361d07934ba62a74388828109efce12d4474298e4c25ac8a6a9c2dc376b55c5143b1f5d98b7c3c1b5c15c50e6d78efdc1ee1223a96458a18cde72b669b46ef5acd9f6c3d8cd98b43aca43f132941ad658f9333d4edb6ec648031ba8440df5f90d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h75c7498a4d72100ac3fbcf183a47597fde1e1f4af846908f56b81cae4aaa931c3b86feeee09c9053c5a425cf05a871d7eea2e2902271f41327cb86e2366fb34325f12862e5a1fa79006727035443d41ced4e4ec441022bc7d71df5eba50047abac5abd31d85efa04df77c98bcd7888a61a9b2ddcb4b6640ed77ab9a41d28833c2496b9f36eabb8663c2b7e8196c3561165030634d7167ad300f3142f3d454751ba4471bf5e7d28a55d968406e970849f9543670539c00ad0c9abeacc2b28b4d54e997e2b8fb4c01af1666e3908297abf65bcc37c890a14fe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'he0f529f9f11ec373bfa474bc37657df5644c31db1b6dd68e63533b7b4772d62253d88cfd629523eefb23f55e00df9a9d616847a56b1ca44bacf982d14a1de545fba93531c97a8895bda8b9d044def730e9376218b7c0eb45b41c14b0748c6ffecf26a02fcafe76c9687a741c7ad8991668cdcdb47016228bb018345ba06f387c1165bbbe292d711ee962146191f730e96fd50400e12ecb7ec429f521a2b6165c04c9d0ee0e4f5330b4239af14730907c508a7864fc3acd740cfe6f88e6982fbef092be154e315d63e8265d3fcda22027c8d4cc4c11bd2742;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h309648022da7af8c2ca622c5662dce84ed046dfde6ec67be478b08b1ce9e6db1ca210c3b887b436f4bb7a65cbb7688b7cc6079ad9b75670e49f46fa8bd568b34a3bcd6ecb9ed34bd1945c1b00e78f18a744a5089df2aa99858df6461e3d29e91a0b21805a66d279bf52504f342a39b249e39db3a4aa875d4301649e15d55281a9b0fc63e380ae39395f11e61b42d5f4422f4707332d63f233a7f2fea377bc3480c6ad99e88c53d40b2b8c5698d160b548b109f97c53c844799291c234538db98aca734664c2910aae56f51d021004c7218d3036d7da9bdb6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h452aec5bb2254c2e6fadec9c35c60f32fb1818d69da346962c1ae2c67d369ab643078c1fd421c2296d9d8ed7b70ea65c7387226a1648621ac0141d9fe86a3b43a980eb95375c3c21b0d0298eaaaa3b9982f67933837342fe8604c88051fead20e4ae6aa000c253893caa5e24bc41365585adf628d8126cdbe1fee1da5f2973cf3d0f3909a18a7c851ae6ecbf3d7740fc9e4d2a39ca7e160197ab411b2d8968fc551f2f2669f4f593b25577f05a7e609b400a0eaddc77b7846938a1bac3a90b10fa88bca08c1e294d390c2e4a3d3d3350b5d5bda244cb1408;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h88094b9c78f3e9546c6809fcb03e93a7e19f02614b7848142b077a5616c2a84c7b6d434aedc7c3139f3a5ceb257263a63e9ec658a5f4031b43ac9376a12e9fc354dca6dc515993ad363ff9ed8bb78911c8e649187fbef4708d95047acbf06fe96fe28d8dc9b06d29be02cfbb949bf9101eb74d889959236ecf9c577aed02ba3bd625888de64871d7e4d103db81586019ea6e74df565d0ecb59139e5dd254a94a7225bfc488f6ea2e06f5dc4ec01510bc6bb7e8285f7c8be3d83ba37984bbdeaff3e9d77eaf29899f8df6183ecafed41032b8da9d61f9f04b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h92034ef6271fd2f71c645e72d190b0755418da131868725a3d7b1485d6a0066f181a6378450cd81ad014732762c6a86f36775323a79a554fbc985208addaf97bc4531383e2eb002bcce960d21d38ee562a3a32cb7b646918cf4ad2501a6ec325a338387843ef87b180b85d31d63d4048dbafb2afbecc50254536436163c313f3a8b957001f2779543f29e24a419a5c48a9e2c0343a0e4d09e11fec1c31ffd3f7a89dfdd36cbed31b7c727c09142c188b4c6f4b6cb84fcf4f289ab9f2ad8aba6f4492ae854dd7595d2c3949631572a8338c997771f19fd37d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'ha4760612a610fa1bac40ce12a276008a4b4dad49c1fbbf633bffb82361c297284ab4b680393d63592c7796b28c0aea618845fec0370b08055cf7523d649b4c6d1936212b24d146b9710934265b4ca1acd9c377140a050041adbb1e922c4f5ed3a99cfeb836d25d8f9e1a520a85fbdf50de178e1d2c580c3f112776eb280584af70774cc3f28cb5698a86160d8c9354fc30b4177f2abf8811f76361707d69467dd4ad210429046a0c23b1bd998639382e4b16d6d2c4037e2e70206449d08a638b8813940178e55ef06c6e06ec5a33413067317762907c1595;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h8d442fbb7810c8eebc8c1ac172157618ac9b0aa6b7eb637788f1aa83d3980ccbe6f31cc781347681bb60a81d3d7d7071388c0707fc469d16fb7b5956e3b84ac27393441e55582f06653e225bd9f59dc46d67cd852ba718b334cb1d7568713d9a6655d939f61143fb01d6cf4a826acff1e6dfac01fd3e92aadc705f2c74eb5ea77ea927f93c936f30d198a1fd3cf744f38e00c51e90095d57a89954ebe7e80d8894a719f5a72ae00e0fa240d8d3d260b900863b11bdc5ea8e07504b54fac61cbb0de8e5dd0b7e589cd9396f6aab5cef28b118a7fde3d1dc7d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'had2546a0fef8336d4b5bff5900e878d35e0afde7f6257fdb1e4f742e432c0b2998e1fae7381b1fb2b901ed9f34363ebcb4bfad5efc21975831a344636b0bef159e44f6e62679cca64d7e75468e338eae6fcc05911a72a42b8fec517d2d25ec6b512128df4859ded400c661d9301f7bb5b2ec3951e1ec49e0d6d7f6805a557b1e37dfecf85794ae149aabd47762f5a1db408d702722ab77b5c265d96b62cf3b993887d399b3f0740b76a8dc2bf1a5b3afd4611bf7e5929e81bb37682b07f8c3bec516e6c0a24005d5b74bc640695324c7bcbafd505f1e5295;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h220a563786f8ee541450ce3476cf320659f37ca507c6eae856b10a93e7b644e46be40b240e04c47e24917a6c592182a7ecb2a3cc201e395c50e0410eb526be89498660b9a6291871b97adb1ed85386cc5e7153a8ac36d3dc8d40909cb297233cafbfe243d715b5b55969a04457e3e8960da4dbe6ff648340d6acc73d0483947ced83803371eb6e3cc44e2adecdd5a6424a302f46c3b19e00330ed6a8a389c025e74b16a223eaff8a320a71f326c08570f2b739ee6107a37d0fb5036faace122dd8bec594e81f05ee6cf9f28fb7ad0172d9dd6760734a47b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hfee29345a7d9ddee9a82cc3d9084e980404494bf9348b36ddf68f61377600682cb3dfa40c3e1a903805fc2cee6ec43f9ee59ab58a4dd5d0b78a6c4a631f3d0f78201b9d9a5361a3fc757d58398190414c31fc60d9a4ea49178b8e1044cdb5df3143fc49913afd178e1840e95024b6bb8119a68f283d3e1b122e5648c967f52e0d6039078e59eec29c1748d8fcdac285eb1f0865337e7a3b25b9c1a50a82e582860494b7eb5e20dec3d2b19cb70b6d3612d4b7994a76756c0b92ccfc33588d676b7ca035d29a64d5793be2486c6ba90a11d479ee8423a77d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h994e77155f976e7ef661d08d39855066d64c5910d3743ad1f25fd84570969144323213f7b08e48cbdd9b1f737fd99595a1ac0881e1a655aed984dfa98a9059324701f0096b44a42dcea8bb64d377fcb563ddedd9b7d4690d10c0affef6f1f7d1da6191cf6a7aa500fbb2930e59e4312d095ca653204ce7d9e7dc7196a81168958167e5b58e18f36f6fd5afa4f1dcfc45c7e3eee46736ee5bfc1153b15f64e49332e2d4890f55490faa2bf8cd4a684573aa421e1d85add38678865fcccd968558a51e74caf13eb6fc8d17fdb0d4328cd0ed260781eea9d8c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hdd2a9ed14bb2188e190ee890c6aa1e6f22312c85ee93bd94dffc6dbd719a6ecb82cc1e69002f78a40171f66cef3d0344fef77d10cd897da469d6b87af51ae6e2aaf9980858e2f39340620ca0f035c783f0f9c489a0b7cae2f218fbe0f7b3b5723b0bf200d582fc1c74da18a311adf4385b89b15d00b6bc2a0e36d4286b649e9aee9505df51d647894ba1337eaa65abb4950f95dcaa5a98a2eed74550a2892a9d8c877f086f1961da480b1e840fe9ab42c28511a831165bacba4224760475fb4feb3e6b4417db8ddd2018537d93188b76a50eaa308e1f4f21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h57beb5559e4e8f505d09dae88057ae53f676ccc5122e3b1b50cbdb6f735318ab2152acfaf9c27cd01a668ce726ed5842467640378537dadac2bf8f3ffc6acdc58701ff3f7805b12da757c39c551284c025b4b9aeac75c37d1716fb957d087ba34179e1472c697a52dd22939310cabe18aa14186830cb3f0265c3f463c59f14ff825698d24e438f15fad611cc4f1fd166e670145aa625c65c15b5650db3e981eaf5c462e18c9e8443249b2217f6b2dbc5af4eea4f42402318e9668410f4d4cbc800877b9a69ba28721e13c3e89e3114af09b7307a7f426bc1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'heb6850460872ce03de9a651bbce5ec82b3483f82ea554805c7b001dbb61ef98cd4085767a577c76a349aca949d28daf4694e82626cda7b4836301f93237d53853f43787d99793f246090646f2b659386ee4f9df2ba380e3b48ee4e5c81198de573a5ade7076f2eeeee6c9aad12a88d6ad16329d44445715afbc320f6105b3bf02e863274d3191c75a5c279f182156e96a1c04b0cfaa490706a16c4a34c1d589013cf3aef690171454bc7d9b6abea54e9a02910d677e988e00f2def61daaf0bf10b6b104dd3ea522aca6424ffde514939d507a6eba9e0301;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h49da34f931e92ae01e120c37d0915f8ba3d62cf0fe4e9a69c61b557f3045ba15cfec75786e0410ff0e808771f798a12324b4d933c25d7799f89f74aab3c6fb70cccbc7120ff31717ec4b6e9c6069f535db215f7266c6caa1a8f0988159ff144255d68f47354c60e85488d304df984663fe62fd248fe9796368ef52296b4bbaa3e3d226cd30a8ef66254257dee6b2f39ce7dadf81446fd2c5000c38d251947818985e4ab01f51fb7567e457cf00183cac586bf1020e66b7b645fecc29a1d406eb569fccfe38f817aa8cb9a9e861798a2406fee91dcca97533;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h708375531eb526b362c1d292362785c5a50fb40996723f66423cd4bb1df17de8d64eaf89e5079cf28798070051bc6e8dafd3fd316162cc6aefc69a8498fa4fde47a899c36f98dbc258bd27151a9f45aa719d3943cd83113f15e6434452222c3ee681ca9153df83623c2188b442d1e1022731b142666bf5faa20f6afc4041a316585b1c0947084a0c0b1fcd403edb283092800f612dd47b7089be6f3d361da54dcca70747934a91003799f54f1e28cc585563ca9e3d059b070b93638bd0bdd6c56310788c7bb848d20de68b2e27d5c22c8db521a7287d3b69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'hed215a8b50bbc60292482c82699fc1ece8ff99e8dba7ee09f15a9b3f7c16c00a551b23e70b8b5a7982747cc3f98be407a73664bfc6597554148f48b53d32f51a55c2a5c434e3631280d36c0d06ef0d48619f32cac4ee7e67f4512bf993ec4c08b48a52b7012b5baca70eb884caa3f685a3618bd782103bdf5647406ad483d0fc3137380e6288ef4e64c795fb0f17bbbc71c0d42c0348b5b42b38be7a5e3697c30b49b144025df7605da5f812abe7452810686643637f6398d3d1f110f625ab541e4995626d6a909ccddd24637a98030a910977cbef6bcd82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3303ec7fc47aceb5e275e4860efde8d2c1402959f198abe851ca9806344c2a0327708b6719824a33a79f23df63417caa41626ebead6b6b9b7314384c7abbe7696d4cd3170216c780865bcd6a7d7af25ee1093f7e51250db82bf05d76ebda18756612689786620b871645e2962dae732dcbff1eb27d269115ba7c7eef27453b9a7421e52f8a1394d5ccb47334085134ec572718b83db33fa70758a2d6a59b8dceb2d2e69a7ddbe72eeecacbdcef895bfbb74536cdd75de6d39d004533e2ee27a14c3763a90b71b9e122e387c79a58ff78ed09b283c8d237d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1728'h3dbf4c2fb82435b0033acaf22e93deaf750598df5408a4b5338d61ec8abbec58b776bca7cd1b5bf00003e073434b29ad505082620515f4a41de5b8e843ae569f2c34ee8c787adfe63105a045c9a5c3a0dd550e48f3ffef2df49d7bf8f9b7e452d770f7ffeb9e18057b19af594991805cc3b9933d6f3e592669235495ae709c11a6b61f28401f48a1529cdab641ea5cad29e103e5ca52c995ea2d5efce49d47283d8c22296c6967c2e741e81b09da0a992f238e4e91c0f96d0b9c05062526b438063564199aa204f991bc6db062756d13676ec00d10aea12a;
        #1
        $finish();
    end
endmodule
