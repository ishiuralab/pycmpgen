module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [30:0] src30;
    reg [31:0] src31;
    reg [30:0] src32;
    reg [29:0] src33;
    reg [28:0] src34;
    reg [27:0] src35;
    reg [26:0] src36;
    reg [25:0] src37;
    reg [24:0] src38;
    reg [23:0] src39;
    reg [22:0] src40;
    reg [21:0] src41;
    reg [20:0] src42;
    reg [19:0] src43;
    reg [18:0] src44;
    reg [17:0] src45;
    reg [16:0] src46;
    reg [15:0] src47;
    reg [14:0] src48;
    reg [13:0] src49;
    reg [12:0] src50;
    reg [11:0] src51;
    reg [10:0] src52;
    reg [9:0] src53;
    reg [8:0] src54;
    reg [7:0] src55;
    reg [6:0] src56;
    reg [5:0] src57;
    reg [4:0] src58;
    reg [3:0] src59;
    reg [2:0] src60;
    reg [1:0] src61;
    reg [0:0] src62;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [63:0] srcsum;
    wire [63:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3])<<59) + ((src60[0] + src60[1] + src60[2])<<60) + ((src61[0] + src61[1])<<61) + ((src62[0])<<62);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h358ff7c533a10fe62671ece87c0ce0ce01a5b2a64f2e0fc4349d960c40723b34b8b2f5dde0686504477fc482cdb44dc3f6661eeef139d021aab64119902a8b1831ee02ea222f62d7684790a591e83f05ccd5c364a3b0769a89fac416a0bc828ebc51845831ec03d7d996e813c43d7037856384e832a3937bb5cdbee27573883b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d924eb76d235d66e9fdf71c757fd93d41511586d07748b35c405d57c352a464f4ab3953c3bb9a5ebb31205d70268e4c69454cf598353c672f368d5abb9119fb21b026faffe2a47c25acd155cbdda0942ec10a33248f8744de752e5bc13715d952c8a196a676452b368a5628ed9a6416e39a1f6e1987e4f1f7101294873ae45c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedee9a03460a7b45ac24d5b300f63087efe701bf97c7dbdf78be6760219c64f48fb36438536b84a77a12155ed56cd345a1c777422de16adfb4fbc61839f5952b3dc960adf4165017ac98232285a9b66952973bfea2ba8cfd675d2bac6d4110e58b27b8f08c414acb8e751c5c6dde5c5b4ed748397b5afab3d587bd8cab5baa2d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e4734e0a1c860cef47930398752e4c5870b4cafed2ae3b417fd0b7b4f7c290d9f6a411c2c621ee9eb1d7b4e9607853d760aff593d3a9bb40d08884245e04bbc9a29708c47b617d10377df869a770a0744f75d25b0597e2782b82f17acb11574c7004a92bbb4979200ac6f40c723e00c25d56ca4c1e57cfb87075838cecefded;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7eed88531e59877499ae8ae5f4050e35e4a900a793ac60d9af4dec5cba8b7cab55ec939387caf8ffa877afa7124b8ebbe6c3746af5e83993616df7d44c40ed79a4b03a0f4a991e3cfcc364c39d06a06d1c6f5a0a267df6a6d659767d73632577fc78526d04b529ccbbae475c55cacab579934c3d2461b5d25c0b052e35d820b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee406ba98db2a4c80cb8ecba8ca9066e0b0c2cae6383c341ed5cad217bfc7ab8cc21863236a5ca143ab24b4f2267e14ba314e9418b0760c4ac9dfd9b6f19fbd51ccf21a753c860be96152f15d39ac8d970529dac4cf241c4cd796cacea5cdaa77f27b662c9e3945db0e520fde53d993e1d0604595a4a65e7f450909f6602edce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4397f84cbb13cb131cd6a931384dbf3968e4c0c48dcf7ff6a86456c804f57536b21e1c32efa4d8808f43be5b5534478a26eefb69e7f30fae872aa14376f63ecb8291058815107fb89bf38582d97e37edec1d46a2399e16b1ba103abd9d3eb9028f41cb168bd9c682f509979b814d7c20e8e9c6f6867bb475a84fb697d3781385;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h556008ee5968f9b5e2eb428ece168b85d79312ba5e336915be33471803a7b3243018e775c2c91334472c43c81c8b319fcf3b98050c2649c6bfca2c038c45274cbd09217ee545ecf1819b73ab98275d8739b2598a5391ebcb791742968ee0b21d29047ffc16c6dbcdb14da92fc38e40a4e59ca41757f0bdde5439f0e808eeac01;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff313c9096688f868a209dc98eecf02d5f7f750edfa8057428f73ca1776a18c8ad5ba5fa5c5e965fb608497dce3b41c2ae70c2f2f307e4e341c8c83ae8f4b5a021902589e102dbaa8831f2a34e9943c3bd6ab806e5e28d23ba3168fd57a3bb6cb2b739263a8d6b47368c66d41c6fcdf0efdf65aa4e6c4b548665099724e8e573;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfe2d3b9d523650d0ce86ce2523bd1673ed30261dbd7e9ebd34785362ac31107e0d5716b9a48077e7ecc8c9c875c502b04c26ada4f7e213ccc518135c6c8fe0179f4427c5dad41ae1d1dfb83358a1f4a82b01090b4d840ab0d90249a9c0ef1952409a94a16a86cd73eea6b2d1d53d21e31f5629bb8054b932896fc0bc5f9a053;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedb06a47217607dfcdc478a17a814ad3156103eb92d96bff2bade04506fdaac99ad5df7e5075832999ec472a6812e10ee6df9460836f4069569d2e4cc1d0f16ab292c9c17c1426af800cb5562fa4eb14391cefdad987abcc1efe5f34a0b53cbe09b866afdcc69b021b712167627c441505d0aee1e6cd9e70a25ad11fef18442;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73583ff78baac928b962f332b07cfc2f435c6f47192595e99b2e1422bec60f4d2faec60d486828c5dd5044a867ea0c5c5fdb0893bd6f067f1043197f16a883bf8ab2c9c880d31e769326d0276c08abc3a0f7a7a204e414d5d85862b025e353ad45714898acd0e86fba5a52a1da66f9069e2d6c9a695641d6a1a5fe4a41c0f9d4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1011ea0a749d783250f919a773a2f5ca504543437280d41ec2bcf73033cfca195a3b1d0d4ef453b350bfa749057475f660dfc1a26157195422922340706dea68bfb49c248c08aee019e9ea4a2f68c266a3705ab87ff3b9ef1075838f00f9d97b0f5ae297f5e557f41ef7e20321280839b6df58bcfc698870d2b2578e9a35672;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ce3b5fd8c12f2e2cac6b77a28f4e4aae9fa493b8d279c9b2529fb634b4d1ebd8b7cc98c74804bf352cbcad099f2f6ab5ddb7f3c00f46502cd61d51b431db297c74e75ff71106f2d8642b9f6bf7b5c09d446e869dc4858d67e996f7c2d926a0ac2500550ff54407e42387a93ed13a3f58b3476e1a41a996458b4d8ff5a35329b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a92637bff4cb51d27f14356e640d974d888acb3147b203a07f7910de2cbbabcd930eac6776f728840714747a24ebab32b39a7e479c8de9a2b6a588807e2bf456c63e2eb7c141978d6d47c48412c1c66afcfb796c0a857fd7079fff0e67a0bd7daa59a23c2bac0f65a448098b44b7a2c13530d4c9d4b0a38596b62fb20cade89;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68b9251670f6dd2c1e01f435dcac8f564fe226c91440b572115a0a2c0b90887fb66729d5c3b1844199af7bdd0188cf89570656bc616944a7f6f627ea7e7e073b5c2bb00a52d034c80fa3aa35b9acd3a20b195a78db9c795d0ecde32095761d7e872dd71a7d2b8985ba6f99f6a9845f4bec8c1fa9aa366c171dbe5fa01f576881;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb93f4bbb5566c447aff0c4fe8b8b42ec64880b3dc30638bdb71325a2efda2b55ea731ed6ddfeb2a8b589ebaa1fb6d808f973d5b3bbd0431c5a4366df7deb4c45e0079bb7d3a5cb5c910ef2cdc8efeb90af45cb753ace755edbb4b2ab50584f95febf3c1b2eca85f7bb203c7b1e3eab42887dbaf5d95a5242f05a5bd44904be1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5c518d2bf7357be56ad863edac9fcbca30ded53d506a02d64eee202fda72f5417a53cb692bfe6f09bd6b30a368a4755434619148b5fb78f720e1133ecd5bf24e99dbe41a198ffe006962730bb651aa70d7dc8fc04c098a91f6a750252f9810fdc94bd823153ab9d3b3f2e0eedf1c36341398c9cdbe5ff43461fdb4b4f9d8df0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb74e492d2123a5feec1e0a070c58c2d390059186736e28f8beff8e9dd6a5480393bc86d61734b606d9130b75cf6e040eb77266cb873d76f56e17ae05ac44d67fbdbf2efaf31ea42acfddbdd27e52871e94ca2de433f21245fb66ba68d7e0b315d3172b42e357eded97bc3efe95bf28e0b5d1043b7734034209cd0d7ed1c1011e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28672182269b47f17e2bb8454632638533ac727401e908c884a05a9c3b52421a236671f498fae260c9fd2e1358237e9d3ac10af40abf74cceb84ecb93fa5a758ba8da2eedda4790d589bd22baffa2f0bf1b253340098c11660668b4731900a8eda2961a30397ee16200e61290260377c94d492d09fb3395c854906a6e4daf2ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd2363e10ab8ab26ec0480575a590aeaed0d7dab12e1c0c86e42de103b3907e2eefd800f975de12c4e6d1cd5d04e93f6897b396165eaa57844220840548cb99bb9ef4ebd435591baf89b064f0b88a945105e5aec0173af81fc6e0078dba88303b8a5f498f1d700397088ff629e30a785a429d770042f82a9501265fbf3686bff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ce1d2b90e4656c49b0ddf10bfd09ef6cb2eed73e42f3ead41fe6d6b3ae3a838acb12bc76adb7756a12bfbba741e1067ccf20aa88b8de7a376b385783907176effe8b6960c84ca02bdb8784123655b266af7288890ec51edb13879ce81fad487e3ca3a69f4f28806977a3b3e511536cf94eaeb1225746a98b2f5cf978a980253;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18ec9fca23e787257bc7b9173b6611cec86cd4c542cf4e508dcd89db09c40a35742499eb8b16698e696c9825abf7afcb76737608b7f49e5b70ba55bd51b901ee855f32207460c267ac1c42abdba15d69e485a40fecfdf270d1bebe5ccbfcc420a93aa8fa6bc9caed4025edc66d8509dbed3cc74450ec111073a3ac27fd623f66;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bd573e2dedb5ccbe3f27a77a7904a7428468e2b5bffbc9d1ae672f66f15470a4c8d69d227f1383f5bace5a4812e49fe2412cc672fb2d7ad0605ac0882707ba3cfbf812bdd847fb4c0a7f62a14f820c74c63d4b7a055f7f1ce510d8deae164c564f97e218b51b717d8667f40524c6491f02a03011adc63972b48b36dc606a320;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h84065155a03e531f3d7c064bad370b5dc5a628df54c206894fe903c98a4ff81d6c5561abb218fc130e734acd2ed82381fffa29a34ed8a71e85839ee9feaaf6dda735d773e2bb374ae03c005f282f54822c769675b06fc6e6c6e064ff1c4af1b94b47bc8a8cefa174da1a009dbce228bfa515cd5fd0ee56fef0c293ebe868e342;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ff47e005d5cc46ccff0df5d409c3217a81285b5ca0fe799af9856e63bd8fe23af0784494845f65e950d66c755ab1b14334c13aef70785a0aeace61cff0139d193a6e078372339fb6c9a2d57ee0ced779e32b3b9cc6389f78b7b82b7a37d2cec6f0028573a0c2acef1dc2dd833abe712e4150377c457dd37fcc26349a537cd6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8db17a650772a714d5e24eb2097e4ef37a2181acf838b51a1ed214c8900f5a6a51018446e618f29d9fae96fe60dd84b7c901f0cd33cf94ae85546070f9f651375beaf4d9df7f37472d81af5152aaf13181e2a08fb29a2baea7d514bedcf2a750e56e25aaa655ab87b11387b7a7023e87adb846f2cc9d399f2fa354d1811740ea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2c50360184e7dae0dd130e71b0ee3a3d766616827f426489731d23faa71db45b15298be77969c04b327fb458709e9082257f04617bbf943882b96736a3eac45742e7ab76b1b766841deff7c31feaa50bcf1862548e527d1a68a0c5cdf7112680a4beab81b591824e815ad3ecd7dd5fe80e899f81f36e97c416d3f57d73497a9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e23b284f6ae37e3396d42676b0f95b689135548be55f03461279dd78628e51d4fbb59d9d2e034b76aafce0d4c9eb9be46d88267993df77c97c2aed704fdc4fa72f25f430b4cfd9e0e3ad6df1bf429c2d69a008b68a9cac4fcd2116e594f1a2c5a9226ddd601d7f19af97e95efa59e9309d135f54f51c77690259232bce22439;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b8c4ae6fc8e2ec0cee6fe00ce02063a160bbdbf979f6407af7f6723b13c53601705d7a7ea1ba7ae95ee3e40e8ee2d6b7865cc89f588cc2947c18cbe84f517577a7e1a5597d3f6fee848ee73e4b3146a0ee0a654f7c55d3e2d6c25e2dcda242753180d7176f2bc6f1d2337a8f80f0b37ccce4ada52101b1e60edfbd81f9d0475;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf401f60128f3eb3c38f8bfd135be900c5e3a5d9672e038ef189648d64019382e137f53b25e85070e5d519b2d7b901c7df86a12450dce992bf1a1ab552f1348f793067091294d445e6eed56a85766464473f166f65b3b763196d45da0a0aeaf72561708c673fe667ca4a9935d308f9ae2c4dd09d9e05be5b0d68540a3031882eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce3656428af508f98e76f8d96d6f91291ab38b005aee19c9208d5f6bb8ab12111faf6292e8ead85a19526b0a13b57ea165b6d1dd7b45f0cd8df4b294aa941d9f7c16973f49eb8757d17499949a633483c267b185234141b195be2a8adca3b51bfeae61ae97c43d189665183b6fa90eea834cac7e63a505d3bc9fbf7defec6486;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d10148249250c9a81c130e00255ea3b333610230e8b22ae5e2f23b3b4d95283416c0a02b962e5af1fed7642b695d7d592b465b3c43e6d4a1cfde16c0fe7d15f6a524cd4e1fc99c680aff929ef34cff0d115370122433e532652ab0057743b739d09e1f0e3cd06e6366b24f455740ed8e7b4b016f8aca0ad6cee2809b4227c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea28ae49b2c3fa609bc39f6ed73f12e0fbf77aaa03213a3cb8014a1e87466418720719c9b6fc6510f97c8e759a527345fdf0c201ef39becc6bf34e9a70058626c15905d48d593a91f735672be8bcdf3e96bdd58511ac49b3cc520c6b277f39292e249e8d37090b5e0a18ce54473b2bccfe3c9cc277edee857e6adfe22e446d4d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7dbf24fe0b633ed4a1da65c6cf7d5d0661a955b52c955082a0c31c5fb0ed160371d820ce24e6466a02aea6f9c084495874ade286b6477ecaf0a72f3af57fa121c980e2e6b69ad0ce04ed0ac32b74b9042bedc612f5875f142a1c53b60ef35c6211f7903a48a285ef2860962501d6afe4b3e18b981ee57b58acaee06bc398d1b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1dddb379f65f54eedffcc32117a34053c0d0c9b05620b7aa160026bcb39e7ec9670acbfe2004c0cd9348342d44be73e829efc4988a956850d1ab3789de8d71fdb5a0b0fbc514faa73543ab62c6803dd94a7c6503ddfc857b7f3045fecad8579a7c2bd02883a695c3d6ac07d6c36fdc5c3c56fe734046b9b38f672a3bf4911cf1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd985ae55474fb225d4bc08b31beeaee48dc3f9d71d805603510880e517f95f5b00ac05211507538ebeddaabd0d5ed310b252fe709b60c5b0ddd97c1e1cf625d116ddfb6bc597d84b47953ddeae138aa501aac23e8c9b52c5dcebb13a17d5861e775bf670ce4ad3a29ce5048601977efd988945ac2b3ef6cdc98d1abc359a4cd3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9be6c2d3aec937674a22f3e3e764cc878dc7389955cf0ca363134755200c1ebf97d44424336b414f242e64cf9b68d745f2a8b4ef3cecebee8815a70121ea54e75d8a67ddee8d776aba476dbf725edb3c7fd4211f2b163bf25f8420a77deeba28da0049d1759f8320e6db490ef2373c7f11e4fe68bb0332ddcbb003e3a82367d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc84c04180771324c79660c8c9d3e6d8a4f56a181e7c41f7ec59f03ec855de50158b24409fc737555dd0155586daa30457a01b4fb1af8577b9d752129d8829a124f30ff19518bf76126b7ee081f001126fed0af3d18207e51c988d2ae552a4a1b95d946044fcaaf70fbf139ab377ce14ea4577aaab8d08e7f157b2be6732ed5ac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdedd447af6c7ebe76c85a805ab68416bc1161ba899c97b5bcd2dec1a2b936e227d12c1f860c9899809e6b66616ae32d999d9300d95882dcbe09fc0e91b10020d44504139d698b56d87978d4857684adf88e213dee0d4364a38b4b669edb91a1785e1954642b362761ae84b55885c04567c1fe2d62f10c2467944c83f50274d89;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha36f462fe50587e6b0355ab1d61c36a030d83f318553449fc77862aff1460277459af451b01c55a5f77b9c938e0bc95a163b38e77253dd00cc088b509b341cf84842d35d46e1bdaf76bf816057aabe319acb2f6c14648a3355d991bb04901d748b54e6e83dda68e28055e77477e54d73e723e45091f16b23b8959bbac97dba1a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79982c56e758ed72b75cd83360c19cf1ac0773c18faf5f7533402b4bb31f894617a6d43b59b3c300ee2ca968adefe3d0d7381610bd21c31e8e44295f0e8c7cb31b00f1e279397bb9b6f8225cea23fdc753bfcf1fbf17c050dd55019b8d997a5ea506d17a03f6fd57934c3845154ea025bb8e84ab01f608ba20e11bfca8d72060;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e914c8f5c6178b890fa49a79d378367b3d170c3b26b3610cbcafb77469c15cb5a7db064675e6aba487ae307069a39cc73abf7f7f5d5682b6dd176b8d17d88bb5ebb800cd7c3dbfc24bb84b782a7545f58b4ab9a4f75868844f4b258e24747a31f7f9c90a5fc76664264703cb91e2e2b943dbde625e68e469fbf8d357b08e1a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1abea8583293ff8907a1db1e66237cc3503948f51ce14142c535e4929514597297e84e2dc626e53554f04dad1f5ca6d51a47bb39016e727ba6fbb6febb9f52007ec8062b9cf8221f442f4fd1d53c91cb9d2c6b4d1b6f014ce6c6b524fe155b337e952e2e735288e557e0d70672fa9115c5d4984777241225eac36b4f5969cb9c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a1e92144e8166150a6a1fafccf30a94437e2e2efc6a74b86a8870d75249337f4a336c2a87096c06b2f0a8d0b667190459eb20bd9f9174a82a9fdfedfaa3b6ff78ea5e3bcec6028aed5c0999a9d486da471e7a6f2a599c9c252f2a1ca10237ea1b5b23122ecebd157c5d69010c90553a32040f59dd66d0d02fdca1763b23b836;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec9c1d2912b92fc32d5464b052af251ee65816067a097ad820b6a318592232f90065e15aac4dcc59bd5b941b827887c12fb19d09beada5039145c285a727546c15b7f058b12c90153e58bcd45d174b515fa45f160fde6246d033e4aa1e8e7b9f72ea5a43101d9702714e64bd0da7f7b7cd2cbbb007539239b2597b2b1d845716;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cf8b586e87539ceecda3e31867c9875bca6ebf53bf00e9f44a87ee76855b25624226c8717d1f5b9b5f48658f8d7c1fb2428867abe5de1a462e65f4352abe8f6d4a6f52a70eac5205d6e37ca0e8699556467d9aee39fa985e508d80c4ceeb35e103b028118bb533189e8fef1011834c4477a8fa39f4035d22fb0a8ccdf314498;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f95bef6935a347b00d35c90a3695493ea4da21a94661c3f0245a85ef7662b4f890514fe1e0c702820dbb56128fca1018357e5b7ae3110678b5b88f67da9d4e8c357d31ef6148db95c2449bb7d9396887884ae259c43f7d806b92ef34a52bec45d2a42c5e7a57a1125298dab358707db4fe8f60683f0c966d64c7659550bdb70;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d4f0f496e4d62236d67fcccda85a2ca73d86c9c6a41968e914d88bbfd7b17039e53baa93f0e40999487731c672a72c068dec822bf3abbac46779e4fafccdd19f616223486982c0ddf82b6ea5d43164a2f097e11649b220842fb1a7040ffd7ade16aeedb140efd2077968135efbd0502de021b804d0e367a4199848d171fa0ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc31c66d80c8ac081bab6741c9db57a1b1e26bbe080aee5b35a8f1290710eed82eaf776f4c926004595aaacd1affd8e5ecd6128e85e15c7a90c42c79cbf20d6500de5c9f2499a7a16c2f5d4aed19f118515fbc70f35bfe4af6c19892ab3c24574f77361526913a10290d08d6d50347f5635adecbd0a082a45fae2896ded8afd2b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c6627935aedb564ef0f0971488fe98a56ed81ed91b02e7cde792195b41d0165c279de75675dc00c61c8cb8038870d4e373397c526dce2d4e32b1d933e339e5d66405c5cbed12d5f33038e75530f40fd7672b3946530407798c9eddfc8f2f0df3a9bbc5037c20a6edbe58e3012d6fac56f5b5df8db715af4879b3b5eb6ee9eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39ed2fbb966a9c2e079894f7cea12f65807987243d35cccfdaabe52d7ef934aa69b0f02a2bb1b06463b76fbca2fe36ae5d27c4e294fa154a7489420beea19354757ba98c52462b705a84a7cff1e350725826b5ded6de9791dd17545eb444f1076d58708cac53b77cbe053de1f47ed4b48c14f1f95fae8ffd764ea7c794117455;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a56bf3b06b829618aea5176dd001ee218e02d526bcf9ff7356c3de25823f48b4ab363aeca4888580e0ddd278e3cf471eaf6b03e09d62e7d5fef3347ccda3336665a55d2120c9442e0b1cad9ca8c482e2b9856239283c332f6216cae139d419a723886705365e21d0a0bb0d76899aa8d061c40dc102297daa8c04c2cdc0ce06d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3f0d3d2d8d6efd801f1f77d06740b168f13dfccee07ced38f2cd01e67cc18a1582a6a4633df340fca46a2ed4f37dcd365d85f3f3313d566170a50ceb494b4c27b3c2f3c95c0d9795a140a92f4023f58544b20a7ff45ba63aa67739a85a0f46b5626d635d7b81d248e2c6722e7aec49c791a55351e2eaeee06a87677117c0a76;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cbe8c96dfa35056e2481e891ffcf55659f066ed28abdd2388c3f05af9df3e44fd2187d07c90c7bd663e1700f6199cfa48f5dc529b676a97f03d5ff963536850aa29d9cfb66896c7f01d7cb6895cc0e77aa320be509298a820ff868ccecd3eb9ab7b8418d0d01cd9582aad819c9a9da90a22b02574aa9958463731e6d3b68fd2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h293230b784a2b0928bf2c60e35a5db61527dcd89c4252a5f877d65b87613cf256f55287613895109dabd9c1393436babaa2a6263ed807c53a381e8795dee2f53bf6591161af309e369c5e15842930715347b65d36839197a8f05eac46afc63e8ef8af1e44fa19ad5018d996246c287155abf07b8c3b28ec4fd1398c1508ac8f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hadc78dc92ed905088a358c66e1f31217276d837e68feaefef8006fd1f5e5006033ee930f6e799de02e6e7c410b58acd1ede9c776b5e87cd4f2201f886900195d214409610ad5862da43dc9a3a7c39a5ff3c49f42c89196ffd7631f205fe10eedc87ebb3df7fd2a721364be4afdb3b6be79e6309abe061c653f99eed313e8ea05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88c02b8ee40a9a3c5cb5f1e703a1d2379ff7de54f591087f616081ebd686eab02f9e516ec25f6368b7c0e6ff13f91bb47970e2713d1e41d31ecfee60fb7ed7aeea09aef9b9571aa30ca5904f3123b77434d57e5530ae6ec40fcfc38cf48941398879fb5d398122033828439369ef292f4a783b57801075455bff82e8df27d018;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h353e18f246976495ffed6918f30384c0490a0db2eb30892d89155645b4dd84b3e9dc86e21a5b848c8ca234e583990e1ee7ce17f41deeacf77f336f615d08ae211c31a61bc6826d92e83a84e87ec5ea7401c58758c747df925c6154708d0e7c058dc84466c53365a483bc4cb2384a41302017cdc4f1b11c3496be441453af07b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e99980584dd6289c658702e33658c8ba5384e2f13da864bc43a821ee08ca361656297f676ac103f456424fe2ae9e2dac546e210b4ff15cb8ecd790249be611dde033db3cfd1abdd4fb93871c407ccd8c5f0b09934ab0d127e4f2d565691faf41839684ca2830a0de149f2e3f4ff1cd75306903df44ea3de6d8dadf5ca8d2f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b21f3e9001c83aabb441e11920891bf1e7fde5e3d3cc714cf4a0920bea4bc6b6d627dafc318640348f96be69542615155f2f6302cb3d1698ce9c549555d68df4d66cdb0dd813dcb32d8c089bca02bac04fed42ab67a514dbc8b9a7142f4b8532eaa6a53a97934ad0eafd763232ebc8de4b103cbb0c4944cee01f9270d440edd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca4b1ea6085b5133f10d6577d18cd21747c526edf2bb51b59f1e1d0d870f168012537e63e667643bb26cce555b06256e1eb8a025033e1234c103834c52ec2cf8f3817922f87e9abd63c53a6f50487a5ac72ba07a8ccfe817e6987ea30d548ff86674f1e395ab5323d2477a93a77f2060cd5ff40125a35979a44942c31ec80876;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61c9cefad1cacf8240bf19a7fa87e99a7dd388136b07b1d713c5d4c02335ad8571e56f25fa5b59db490752f294c23a51237d5d9122befa28ebeaab0c634c03fe263bef01a11045714f7c8604545e2fc8bc689435447aa974e10af9a23932d0d77f9156efca22af658d99a38c89188bf322b5db16d9e354142d7f94ca4b6c5528;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1df27c3d1b1975d61c9a4b2261f377d606a44fe641fafc391aa7d69898311762bcafaae119c66fcbf04e21d0c84a720aff61ca771125b36075d5d2de0aa136cc9af2d85cb9434865a130ae5ceb837f4e65a00a73766fd6fa153a44e7eb21038da8d9eebe3095dbe1fbe543697a67fc2275d104de1474d68b6153dafca64e15ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he216841f3b3e275e9b3c3c3cd85491584fefa7e0e39cdafedc4aaba8004e3192cf6548de2e77827cfe59eef1701174406c8e47e788447fee901c9f9ca1a0580ca9b89badfce245966bdb7437301171a316572158e14a972f9762fd743a8f55e5f35158fe0783fa20c92f629297986102b2fcdcdef2b8d860f1eb393e235fb149;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd51e008b473211e248d7e5d88eefdb860ef8f6e35eaa86096082b542b0e7de5608cd57972a7ded760491dd27b2ae55a5f2e831c5d1914b3af66a30f6faefee4269859573f981459ff77d8aa67e474f8c605857e80f031842e51986974ae651f91a138586cb5e514e72b95fc2975b111b3195ff55cfb8b13255b6e800fba74dde;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b6893554e68bf936e7fec0e788beed718867f05b3e53c2c28b9e2d3b6c431e58461c65b0de4c199144e43770ec9038749d7c69e788b7e577553a45cf76258689de527cc162ee000d9a6709c6ee121c6e55e0ad6acfb669c66b65b2ecaa2a03aee37f9f8ca58e49528a51016683d164d64c8ef293093c46ca333b94450433a9b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b81fdca5afcdcf06ec1dc0d6a14a82f20aad91c51e4a2621194af651458b5ae79d3ecf8ffcb5980afc93daace9921046b73864421de29874de8ead53bb13daba816da2d10f85a2ab2f5a14849cbaf80c19caab7e7d4b853df85d0154d2502e17ce1c8feac8cf9a931e5a02248db65d05ba3ae8654d72f230981fcbc601eaf3a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf9d00808ac0974e240c108b95a082469afe4ed13424d58c4a09468814be496604a61c39d75edaac56bd12e63fd7df64ef38449148c369e4c8101b3d6fe97d8acfb68654b457eafa46c04e2754d571457149633631d351fc8c840d7da7fc93c01ed1865f3f5b7c11a4cb745c9329e3aee9f0ef9c406c4205edd3c76d0eefd004;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19110029195b2a79b09140990ce92e48cf61f94828be7597a410c4159253a4151d453e1ed5ca3bb834b6dce78994ff8f873293db38bbe231e542aa3ed6e6ef3dc82fc072780c200a237a5432d3ed5585f2b42a6efeffa20cd3f58f9b3af01bff0e698434bc0ff22c3481cec4ee9e4464cec6bca2ea1e46d1f3452634165c8133;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7307fdbb6f0861d7ea1f0c7f7ffd914bad583155ff4443bd4bd9474a5dfc910bad9920519e2039d45a84dbbd8ddfa5d4009cdfe8dcda8f5c19b8e9dae2d8ff2107ea234e6978facfc49de3e4a8d928c7edebb28028fc66c55c4376e2b89a65dfb998942979a80f8eaeb8cc99c061afa47076f00d38fff40a1b3bb898326de80f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he10a669cb40ee4c2d0658245a9451ccd42dd60a3007993447d19dd3a06203e923778f283096cf3d7e24538bc600aa80315cac36c72d69afc0f9831ba40f5aa028fb2dcf6b6e53f0fb8c216a53e1d2186fd2a2bc3e247beb4f1773cce766d3b8b1c652873e91137b54bd74c588628537f439fbba57f93b7eae61f6ef2985c169c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28529ab57b97eb0877680d411a45325d0b6e23d6eb3c5b915ac4923c9890ce85878fe78f6622603eab70eb150468aa66f216c08178c6bc3f90518a7f24f83ff50d8a9d6e46fc24cfd80d4918d99ddfb0301d92141b4df18df7f78d979745f61cf382347f730195fa61bd1e9ab0e29fa43fc7f0eb5f1bfcdcd352bd8a86f2b1ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3f016caac4357f42f9e5e53111ed2cd5bab8e57ad540fec2e0b4f5f5647da74fcc449012b4e258678dc0796c8c65e980596c3d83c773af5dc73fb7387bdfe4572e55b4131493c2f215254c3bffdfef6f706b88cba31485946eed3c1231b9fb3536e0dd23234bb9711dbc430a246856c3a88e5b065d557e341c9dcbbfae80ada;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6e128bcc768a0ce5563d12dbd2ef6406eea351f512fc58e9a1f02c10aed38d5771a5143d130688d1e6abe63dd46c81d8fc3f4ee1141e94e0e9db29202fda0bb05dfaee201b51a4713acac6cb6cbde2b0a7b487dbdebfa0446d2d89f551a4d905a2025bf6c7d29252235355caba096430b4083ed7fc1a822cb5995deb91fa919;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb4d7cee482a9ca2fe73aedf83862fd149df36642ba046e8ff0a4d6ef556292fffd6b12c5304079eed754eb51138b69d801ed65034dd600bb700bc9e778edd89ab2ef3b74983e7168647df89c034ab00ab26ddf26ae8c9925e958810f1f13027083f40e99ec25e2290d2b4b829660523900a64b4895aa247e1fcdafebf52931a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1771d3c1410e16e49cc5f0c65d769dfbc9b624420585501af96662b3be383a40a4c03e914aca23f25c96c6174040681ff4681eae6dafad025db503c4a0510994b444ec416e2ad4eec943c2b068db33f517d0982beae51e260e522082e77c454bfc21d9a0d6510322ab055e8261d8ac287a80f97889c25ef82540b3452139baea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h271a01e2abb92b809366e6ab5531c4ff2411bc6738faf35da35f61ad791386cdf3204079520f20904046c07529a0b1c7ce70518fe05ff3ce5950ea1cc5c7732e67eba31cf7e8d667a0d29436697be6df226754b0894900a8fbbedbd11155fe7032b8609815f98ea5c0fe918a8f3db1802169e3a91b608c99e00fdd52a1750406;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5ae4cbc612cf5cfb267e101ad48c9d8485cce77a9d8c18b3ff49f0a98cd33f70a3791ddea0555d66595b072fb7c5705774c5679a0427a7abe788015667c888eb5fe9e2751ec708ca8787f65b390011819a4b1f96838653e3b04a16cc6a53f56325e9d7f16760756ad3d7ec9a70584d587857f7a48dbc9a6699a0f513936d2bf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf12fb31954e2ef8b614ee342f1e7c230b577ef221475e967ae9170d0878c76eb8f408f240a7f80fd897200f78690d5f0ce8a545508c12742176465482818e54e568dfbbcf3360beacc2b03ac02b66ad6da7e45a4b8230a45b40ccc712d7b2325b827952b66b9f3a7c8a05f2f93d802d4eb43ece8541abf01322f2887b102325a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had6a262cfcde9b13c1680ce69412cbac2a65ae80833a39ea8c4293571647eb319d786ab5c243eac533968241f65f2e6d42bb84446b8fe19760a43e8a9010817319fa8f031cd088583a83e832be619e85aeabad1665df53ab8bcc6750c9ac869b04d33029f4cec07d657b30195931409cae0f2b522d83240093504e737385f939;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he13f879bfad43aad66f3b926063a5d9ce12cf85b9fad5413eab60b1196f85a6bcaeed698f6ea4d1f0e0ce38fabeae93accc6c4c2b33c44a25e2d185aaa6a7a43a9026923b0a28dab7818e6d3f96bb5ed3d100765231e805c9bffcc63f2fed1851f3292e4d80d6ba8c030c9edf6ea36705b6e797fa464fc10cc454f897fb1d02d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cc8ddf83cca5a26d9f82c4b0642093a749d4303420e1e49123fb1fb9e0783303ce6f5036798e460fe5210b8223f10339c626b9644ada3e5fd56ee152649796183e16bb6c59d4267351f71307efbcb612b176072f37ab6c5d3184f9b8da19aef4da751f920a2b83eebfc21c412d0026e7904353416787396cf80139eac307e2e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf15d8f6efa845cb699612350baf24f51ef0e06634882800776c2bb064b4c2b9ff65537cc438397e71022dd56c85d032c54655715807e7c4b747b8e462a5a084c1dfc990a3c72a6997a4ba35a6a346f4993e4bac67824bab72d7a72348d02961441531a90a6674fd584411a57144176418eabc2fd4b4e91cc6ae4e7e3486c59cd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12b14745c9cb636645872a8258ee766c7101fe838e5b48da2732113719e0c4bbdc1f41de25f889cfe40dcda04808ae233a8bb9ad49aacbe9c89610ddb13aa227a1b3443d8245b36268c008ce8d5d0b3bffb59879629e1e1ff68d3e7a7e4ab8e32cf0c1090fcd7fb5fc258246eacfb02da85bf284541dc5ac8bc8b2559f9f7710;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb3e5b9694b55e624faa85a28b90f9209655211189ac7dec56586cd194b5941d2e08a23884172efbc9f144b4c6fd3b20303960edcce2535727ed02ce36c3dd820c63334cca55b66607ac52bf1a5186a70c60a9b735a49592c5368d4aa97c3aa1ccb042b4b2f2e461d06bce059aa7512d46205d0581ff26b257a951798bcebecf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a99a188ce80f5c6cd8715cc6e2d6692321998f74f054df50247b219361e4abe7ba27c7c6110c09f2b8aa7baf87ecb66c00090f6841da8ddfadd1d3bc82c518a45fcc9fefc01c0d8759ba394cdd9d662b9be49c1414b95f57e8700bb9c71254d4b6ce1c5bb0515107ea55640c26cd1a0490d16391a3682c58e14aa8810a91749;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12ff36823e15dfc96325eba4a8d6141b97f168db1e620abd7bb7bb57a512bc7fd17fdc96f30003eef7429a28f7b5c934438e5ea18b143dd878977b9b5b882e4c8f49d851893630f2425abfc5781f646e3a73b0d1e5fe97033f81095f33c408190114ed685ec75c0d4cd57e256c0e840547981357e853fe09c8f7cad2efbb34d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85a717ef1aaec756e65b17149cb83ebc8887f644cd58546baef1255bca0bc6cb47537afcae5a374a461958ff129c8e513613cddd3107b561ee087db8c1d731d47d6eede176cad018ef54aa8df5534128fa11d0837934780fa409bbcf41f5bac6ff0c66dfaf8768ce1efc7e55390b8761fd09dfb896f35c448887f0ea05659258;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb01ef5823f7c7fa04680c4009fd5a2ccfbd56b9647fc67d5589e5915c704f22a540873943dcdd46d04b11cf449be19753dbbedcdf8ce2b6cf3f7b53bf61e1025a4eefac55bb7650aa7f2a8adfbaa92fec38ae6d0f9e0a237f7b47d39f4f40b945692c087ea6b5508993b686c0a0f0e39391758aaf24bf8c53e1fdd9b4ed0e42;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76ac83781c8f1b38e76e6032d7ebdd5e0c912ae01b7113fff12aee2a047983c713bbf4971e60491937361fd28a550f0697351d887a4b221232bdd0f19303c0596f28494c8c80a78c537a31b3383a84ea112a50f31890e9fd30170e94d2a359a7a42c62f5bf953f8654600f050af03af0e155c9dfcaee3a36c530895c29744b4a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64c19943103fd56a7ad01ab9cc1152d4b87a0061c68e60fe8bef859773d562d88074bdb4332faab938c923852de993900fec887cb8245bd61dd42ea60feef013c0fd9f55474d211753d58e232148c04e30f18c0978dd27ee665463c56ea0e59fe40ab9084dd3a88fb18538147e5cb7e2697a13b54700930e2e534d1383dff277;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36ba5cf6194a79df3e52e461bff31816e5892cf0190dc8ed62f9b482247382093f828e3c521b471a6def501786a45a1bba58693638ba3d230a73f9af79ed24616d081361c8baf06cc0b063f083346a43df9e24107172db8b11faa9294b919b1cc78358a021ce832a158292643f272ad82994fd509365b3576c65b6ad678dcf1f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h134d8e34cd3d82580248e8c33ad28d44ea13e02b48880f357c6fc3f2470c528a12551546e248e95790a9ba7e76e44e93ec613d391b6bc665a0d581515584decd2303ea6c4c373a97299ece9a94174152cfe8f755157d2c1c2bd8fe0bff139a432e9158972deb65b1247a5a757aeb7bcaa87b7004f1cc57a5f84f7dc4e8a57900;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3f49f4d1c188e45d75316e94ad91fd9f35268315029a751a771680f0a917dc6e3e6d842e7589de5a28e5fdf74b2fb1c1a960585e32cc0b4de44580100c1e6fbba5863b81d64a229cb943a1222dcea44f4409dee089d0a1f6ac52cd5bc4bc2d29ceaf62c7e5d47b32e37cab46f7366368a4af34e9f69f005c7db283c5093f3ab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcfa44b677ca14fe52f1b18d947d875d3c472f14b1b797ee4510e6c6ffb5f3f43a906b7352522e168745c061fa4c5624461412bc2f714a4b26692efa9e107f57097031e3a515ae658c3d089c36f1582f359a5ebcabaa12deaeac160ab5eb4e4b50d0fbcc520ecd0b61da477a3d53c222eaf7665af714a28340eb01936a9c35bf0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h173a9101d8a0fd863e60ce93684058795b487c2dbd7229a5b2832466a084bf32c6e04cc5225d96d4b0400e9571bb0235cf6c1f9a919356bfd8f70e55d588fd7f7a8aa31f1092b93ae051d28c12d46aa1a7e8c3b053a5d5be5299c6ed68a104b19d6acc9b392180aa66c286bdbc4d12b510d32cd865af11307b093b773741946d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h768463c272d4a6c7d927dca0da78534190a460ae1ed1438124d74b2ac613319799ec4a92aae05b095138ccf0f2455b18c311e4b28284e2ab5adb6f7c37642651489add85c4672b332a1fb1ccbca4d653903b5c757264db343004182e7eedc62b2ca38568ed1757475947dc09cdd0fbf1f406a0381f30ce3b38508249eb88b3b4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb83c8c130a53b25d06f9f0ddf4e2609702b6b601bd19af035d5eb9aa2293550fa07b4414cb3a887e079ebe5cc2ef6270f60fd4ffd13ae89cfe626ae698eaa21bcec956143b29323c9bb7757890e61a2838dbaaac256151fe16c83c6c486d1d291e9a492bbce6daa189acd8bd3f5394ffec5b439dee5228ef71cda86367614ed7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39bdcffb82c17439b588309accbfae0517660c6326aef0f28d265ca93369ba4fb797c063d4ee7cbc6097f70e31aeb712f53b2135978e24eda1858fcf4f8d2552c416c0cdfb665e464f8bc756b36f44c1884cccac68b2618116a7b74a414eee49fb38dbb88d8a6eaff361c0ffc0944dbd8729769e2e2309b306fe98ac2dff4d06;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3af451e98ce214d26f772397f34e5466abc529e3b5a7157b4bdb15e2fa2c146dab18af7d7c087df2b93fa07e58538631736e692a19eef629bd6833e22a33c1ca6502dd0bef3a6f954354084f9462dc625c4346b31b1b940988248b8eb7b8988c080eb3a38d70cf66f35ee28a9244337bf9920e1d60e77ce80322ce0c75f2554;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87250c12c7162eeb9af143e9774dcf16afcd2caa22a09e8449dfb0421a347e1610a2b8b2d5d3f8c586b40b6efcb1563e69127a023f26231e227446242b817861f930412b20ba81cfc48c38b1fae0525b3107644c904ad7ec67e70d2cbf5b210d50afa3a6d2b68705e44fe7ccad77980c505b28b69deaf2d96795072447311130;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69a344bb54aada1ad9ad98ee6c75748043e5633488b2dc8ac8d1fd30d3a35d49584955dbb1aaf35f5df0081434b1e9979e07c23caa8f0fef014381b1d915b26455b453fc389e45889ff8d197e2c2f3204cce6cd7e00fca78a1b1562d3565a4bca0b617657d8bb3a181647ef313e6d8c3a9d24d56e1490e7928f270c563fc59dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8701f3735ba28ae06cfa737854f6d02ec4422575e1a190c75137d4a77e157492880d3d09b4f328e4d4d36ca6e443a4058a1fdf62c12d59198956a7692abddf51e4186cae65f3262b48b131577fac222f225047d84b3df853da26d096a266b35f159151a2e439a3f7e4db697af6027e0142e44cae82a91eed5d7881f1bb60a02;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf94500f2f9b899bb4e022e1b5ef24e9dfe5f5bd4974bf57943be83bc43a633c944a3e7f4d407771180c00a844d75e7267ba8a15f299f32e2fde708975f31c0a5d0c563e7c707bb8bc8417c2cbe5fae9ae6c63afdf287384202f68c35990bb1aa964df746029de35bcafb0818728b6d7a217f55fd046b94fe0d5e77bd186976cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a489054ab5b8fb51a53c6292ddb1eaeaf941bf9767fbb979436795e9ca0eebf83197274a74a0f63c054727fc226add854116f6de2675c7189904523b84b4ab371ce817c6adb071af00bfdb42bacf2b28047be0bbb710af3648cf4a351922cd54b101991255a2b892c564344683d2958eef3327213d3da5a566216ebd2662171;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26be54db094e5dff1546cc315e2750f83bff0b8bdab1f5cb23f5a63d1755733c7c36447f65382d9d086378ff9c02b4a123a1dd964269e5073766d7fa46ba4ef8113412d923ba800fb8b22bf967fedc90aae9aafc22a78d400f41f1bc25bff0f59d403d114827a050af0a592f2f84fc4159910c8cfe496ca03e21aaaddd2cc96b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15959f33853dba99da59c3c4030bafaa697e70f20586bbd9eb16872f90701a2a1902c51cbd61dbd8ea9ee3ca0c82135c1a4c46caa80c194bc45eddf7ca65aa0e0d8fc0214ac470dd179c907f03fcbdc64bc89e770be42b486027babf542d7a07f77fc85e8bc37689d17204f20f735f2d612c39d12462f4284c626155a34f2917;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcef2b258542a0e68abdb500ee19371148a55714f58745e5c4b82b8208084312583a83e241a724b035a24aa5edee4ef08a518ed49bdbc9d98df39c851fd1ab8ff3ae1b1a8174704bfd3d05211010a4ad6b9dcc0552999947170464c939dfca23850b691a478485010736871130196e449971ce2490929ae8f642d58f3658c5728;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98d54f482d2f8455ee246e7fd18bbd0b3464a9d696f0fc4d89da87e278a720f995819566d994d9b296ac007080bf2bea677dc92bc4793c0036c2bc479541cc8fea741f13458831b8e600539fb7adb351e1b090a95d926ed8ceae7fba2e9ca54c5d31a98ce290bb702be0b1a6c1fae3bee00f3847f3b27c2240b694f1192a229c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3af21c5db9470207ba948bf0aa5331561a73e452655155bc90ff2b41d3b2ed300562f9bbfacc87df380f551cbd49034c404317bd0ba53285e05c7a21774fc833c0d770ce57fe447a6c150ced2a57fcc68f8577401b396514af8a8011a51bed6fd2841baeeafeeed5c68e32b6b7ddf73071aefa82962721b003f021de753a61a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60efbfd2e815c1a989641796b69d736dbc81006c4f7d3cadd153ef105235ad984c80427db1ba5f8f4e70d9fe13773be728707e3ee2db2b7231c4442d40d39e716d0b80074500eb5edcb6e5de13dbc2419e4f210fd2f38af0d97f2413056071e3fbc3825cc93324d139ddf7dc700087e7e72ee60c7fb23489468c1dfd33ace9a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6d526a5a2e2487cf53a3b5459e2e679dbfebbcd3de207f031243ef19f2ba5c9068c9ce2d5ffcdd1944c64a3ae8bf8500d85baf0e21e669f8739284bf31b09fa7e1c7e7d1be7e3538052e7e8119525f240549524598cbdf645ace4ba2dfe98f70ac01b73360c204da0eec0ee876edd7a63a977ed2097b8c17882d421ec7cca06;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d1dcf1035dbf6c2be18f8730340d9d3d20f8f7e6fb58012f26a6b8d1ee55b5a96129a69d8ae5d06b7a79310397c7e9b7a2cf690a9f62c7f08125ade93d89909ce5cb45566a496863650dd4bc8fd6eb08a04231eca76bba2bf878ad291b21d98e4a0ccf3ef657a5edd4c4099c03274b25c2bfda3e281b8948383b677f063ecc3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46c56be0863a2ccef08801c7e31d93f07320b20d088c494e376d310c518d146843f46d168de56888240f42d3ec78059526243e704f644a75e339e7e9d16fb643036ed09e1a6ad45dbf0d9d28f9eb0913af6952c93e3be3d25932570fefbfaaa802b135ac707f1fa149e65320fdc74d4058dd90cf939db8bb52408b3b306b0d52;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5ed26310263439c5e51e88003f6d928c29f37d8f64f1f03b80a3360f0c0d8e275fb031918bc54e6e6d51f772f5c18ad215f9db8a1c358f47ced972f43ea4bb1f0c0c173149d4f74dd4fe0bd3fe9fec446fd3ca9a8b5d0f1bcb070099c2a52a25e3ab4f129780c6bc916277ccc4c727bd940b12c8589d2a279a4dbb7cbdd6dd4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h872282b26f67aca169ff9992e5b8c96875d337b90acde011f7f6351048cc91ea27cc5158dba6500a083462aa316c5a8ae11865e3bd72285d4c8a0c608dc59adf77c69e313c7169e4e1d0152caa0e64f6fd1bef41be10a8959871b7481bb0e9814b08cacea3e198f7f2cbbdce43871491872d58c457f7c5eac1d94115941e0892;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e53d5a444571bddce4cc71b867750fe3ae424ceee1c10c157404bb70488f21dd1afd19c1af0ae358ce668a30d93cee71d5bcd13751e0d7c1b1bae37c2f909f3848eac3fd3be116d2d1070bfabf5a3b325b689ff38baf6066973ff90b3218f1f628d84517fbf3d6b6302082e046b074278aa8b9a69ddacf163a8e73ea110e628;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc031b3971c014c03b773b1f942075adc12f851ffe12aebdd6d61809fdff8b47e91751298fa91dd26a1705cd48f963f76c81d47c9ca2078545f40e1e34ba674f9e36492c5e96e846d63af1d56495c9bb4da488432a0515488bdde0e5fa9c712a8bd51b6bf42e662a030de1c93ccc50a3138c7ae83da84b07b0781133ea5dd691c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e0515334fbadd636a8d1b5f5ad862a52168a67593ef2cf78258971c41560b9c561b01fee10f18c5aa661594b3f84862173fca33f81490e7061d20c25e6162c346cd0691488c6fd42e7c99f2d67f0135df76d1a5f49d4d1e35b1905d2c2bd63edaacad7517bbbb9fe5850c175b01572eaa66c48dd234645bb217089da1e69307;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf806ff591c1ccabf71cbb2b3903cd7bb8a162cd85c5638090f9b46c83433892f3a9b57f4f5391cd93878acdf73183566f9011d4603f655b897557225167f40b02e61c37e644810d2746c0a4ad081be05d125e34e3a767fcfb374ef57610cde8036a2df751b4c4f8c90ef53472efdec0b235f525dcdacac599e98f160aedcecd3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd17c0cd98285af72cc4504304e7e26880ac29838502f230bd223e3509278f9698c95d485946a0691c7a55c64eb8ff0b8be6b49d6a0602df40bfefcbac80804cb1a6acdb172e95f0073d66cf184cc970113981cae37846767a096fa06ef2475f66987b5f7ada346b273b285796e3fc78113d3de7c5c9780abb945c989d9fd4919;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18cdcba0628f6a2f5c66de86bc4c95cdddcd467e5a7e9017e7489f081a913948e54cc24eb7d9d7fb7b69175d0c5ea6924490589b92e0dd1f58c3784c08d0759e13481c79e012c9f4079a7cd8dfd17fc1eec474138ca206e0246087780799b85e56db1e29b6c8ab5997d4b8532ff6f8faac138ad82ea7fa48fc77d423b87b6127;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3052f0d33b02e042d6dbd8c387351b4bac561d7892b27dbb4dade9e0712f1ca9fd2944716c13f161b7dc5feac2488fd3ab0c6bcc32f96b2392f2e1e7ed6c0bb8250b74e4608e0e28766219e07d93c606f98472ee49f13893f28bfa480b25a496569ae5729de0745fc6aca111fea9b77f28682ddd35a852ce9a56bf7cd5327d13;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3211fe237ef03de066bb30661a6a4192cff7d0b89835f61d884ab6347259f7a931b9cd8287497f1408b9bf1cda3bb0b29103475c9f200c88ea2e038c323d4b48ce4bc52601387ee9b300064002d9bba58c9130f8d917baaa844cf06af2d47ba8676148e8487c582d6ebf0dcd17fa4b29e4b20574517d979cd272c2c8b2a23acc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b8a365013e149ca4ab0a2d25c4ff879bd932690e2a4411d06c33c4dcaa8744152ce18029e762dff53a77088afb49c4dc0ef35b2e0b16b7e4151679b66a9afd3c29457adc40247cca2110b7b7690cc7e8780395762febbca09730f8fd5387285dce15582a7275b269bc824314bd12d9b4e1825b3ed1cfe642b091d5fae9d0bd0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h234cb59036f0cdcaa18955d134bac738b33af30a7a538c2239034883f67d15cfc1d09c7e2ec7d7e1f202ce08b3e8d172401e7dfd06f0dcb7db8bcdce359cce12c0a8e3b746ef42b515e823076d62e2ceeb085d2857581a84f7f08d4b68415872c32235c52794337bd230b02798b1d7101161840bb2138ecf263e876bb6b26898;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd26ec233a723aee0f99079acf1845172da9ab8c6d0a7629632b674498c4a4ecfe529a926fff1e1e907c553fa1265d27eda1266652df076a4975b1a83816aec18a3a243d9af7d1bf140d460babe80a5ced1d1f830ff5b81cfba4fb2476fe2729bbe96f75fccc23bbdc4d74d16b9cd09239c22424c32a8fb20cd3c7620bce1f7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa7dd750798fca6507eac4e0363616053a5336b25cf1ee4e0acab69e30646637af2d6cfeaae5ff30112171a98758bcb6a00b8d6c327572b7ea3017b8f462599d5f2101ed160865a4077e810859dee8cafde066b5330fb82276eb12c8acff9f657a0d53f484a5693ab1fbd6c69f6dafd5116bc430ad566ddd237917ae753dafe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e4f38a470cbb51c5f1c15b1de4962b37a2db7c43a353dd6aab088cf9afa58c409265a0379204a7a205353da3181f90bac31cea72dc2b8bd77d9a6311626a21f29f2c6fd02ee0c350dbbf730182a461b037efb666b50cbe2d01a62a8fc9c168f6414138d23de89ea6ea1cb34e305b13b2adfa075a3c83b9367e8326e2bee6bf0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4dfc5a3a02e18eb89359bf1d7e3a671d4b91f922937a1a7030fecf6390949367673d8b47fca600cc113790d43abab3eb665e91f1e906eaab30dfe97e659010da7968d3577cad571479f36a7153e07f6b3cde013e397e58f4912718a90093ccd0087979d08d8521e05656d11d89206b7f2d2536e862b280028e3053b987e77556;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb85a156ccd09c20d74a2b04123332a8301dd7bab558c218802ed1adc2ab1ac0c74120927fa2f73394b2cdea6a9957e75cf309ef2262d8e650256d081da023ee0a02904412c3cc8b8c1a03eaa30a8470feb22b3188f6e3ee455609403dbfcdae3c273ddd38f9cbcbaf2ee9fd1a4125e7ae00934313e9478a58681a457f76ace9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c92e20d5dc1de9329a2d88c05d179bd7394e664b794e4e41f72c898627aad43e7942ecc425072cc173b2d602270d1c5a5bc526c742b50e29387727989f0e923a9575facb68304f3c1248b379afe9c632a46b9256e61c88d38308d7a262f06a5caf09dd7578327b700c46f2016c1f0c4105a6c545a2ce89151005dfe91ee93ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae3ee9c097896fecadfa122f15815a0687935aa36ae5a9ad80b118fc08427695da24d9908d97c0893d2ac682be3e02f0584a01d0656c3de5549483db4af1ed3c3a9f21d7e7b9648efbb5b24099970db8d984722da1a189571f46f6ca4654a9dc575022c83429dd592db11e555c913352ae3f282a1854af45e179f21cfc679950;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bd96f154fb3a9062379d3154429c790a4a5d4b1f39cee3e4b021922c377fd492d865756b7069763e658f95ba09c97cec45cf174614f6e9cf2e5a01cc47c74bd690f4b986140f25fb13fd485d28924a1b9bfe4782bb6cc08502c61b828c5b8148fb805f8efe9af2400cd0dc944130aa9a72d59d505e57958c93e276f0514f012;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7305662a32867192e8a1b00306bf762422fc737daad9d3b2983ca101ffd22d6a4069afa9ec36bad413df0b44236a9ad2676d35dad4089215bce382c800a90eb3ce87b288be061e337580e427a969fda3e4319778359ab9d809a094cb32866c4af876ed51d189778a1b70d4a151eb1c0f2c6a90c59062142aeb8b46457d08f62a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cc91882ba90334d89c4cc3d562c4589317b77c6a76c4d38a01fb34cfe562a73660578c9790148e6e6caf91dbd59cbe4e2d799afab7c341de91b4d9ca99dc17cc71b1a1f0d45c669e8f024943b267eabb58af1b14791ac68c2efef19f0c4792118fcb4b038a999d75ba420cfd72ef718736f080c6773070e1d5af9763e0b6057;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba6efbe5438d759a972504956633afee40fefff773c87bc189455778e49a917ce197b86ca9d9467bfe74d941f428dee9e45a1296be1a1f51e6a8da622ad58b686691a45fbe7f30991707ff34d522b2d7d7f5088f97949f7913c897a5d777f0db382db98a468a6afa09ae1b943a401f23ab45630c549b488c3badd885173974f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb66df36317e1de8736d7a4b05731106a7fb67f1d542786b0c89fc23b10d0f960e1de368587bdb5ec48296a58ab9732de0135f16e30198aba7134b2c9083a400fa74e680a64b60c7f70624372c751ae60650247ed3556eef09725de539ad4f5eb385440a7ac4f9f5ac089d0129a435a2fe07e6fa6f5a7e55e01925f89da00f4f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h970ab449b55e38bfd63388e2358db4bdc1b2926a9500393dde23098d14772916ef9f6d8212eafd696f59396bb0df9ff1d3083f3a0d54a263bdc1fced952b58404f2b5a1ce4ae5c2c81395850a81f2c4de1e4c4de10280b5e75b5631e731e906988f7cbd9766fd588005af9b5819aa311765aafdb93774f1246f70030f4a9181b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8231ffaac03a6c5f931634ed4d27d1b10bb19e118e0000687e153ac7e16c41d197c1979abf7f03a03dce6a4703f918e6d81e98f17f073aa89c1aac578b7cb592a58f17dc65e45a382828932c4dcba33f88f381d20b28b3095f8bfc255d43ad93bc8ff6c8e2728f79b84ac9c37404b22303f225286c92502e58af41dcbd791f67;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf9dafffa9ca56fa2dabf61a4520138854adb6c7af21c7a86174496fab8dcd38d48e032f3f6d551564cab36a47c396eabca32e459099072f8ac7bb7fcdfdbc13a099c7bbdd2ce5656e1c2b6bacedacd09b0e605cd4de444735219bb5916a8b13282a15570ef0865c25ee8f7184534a797e23c6d9099ea30592d5deb095cf4c88;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf1585da825e53c04080ccec95b5d76ea2667fbd4ccdae478f9e4c24ad5e7d45e0026429131af349e760f67abf997b15532be486a04ebae0278c52732991c567fdc5fb72728e9c1c5af32a704c126621034df385eab0cd12b49b748a8cddd1960d8280b0e4880b13487a37509b1cfd1ec2cc8bbb9a99d421e5d6355b1f895431;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h220e524a7a4c1419b1140b02f089cde53c6937e41bcfd95f96cf53bdf761d7a1173595b57659c186c3e0a8dfb3b6261450d346fa7d0164a525edd0918319e6072d0ee4f1dc5cf8d631e49d0ca2d42eb50c33295679e526ed66f572860188909e277705d3d6f33bb932a1b5773caa0628822774acc32311931cd9f2745647cf1a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b6a9331a23ffe7351c142bdd3e8c0a12f6637da025ae42e82c14e38e6a6642173b46564d04d404a45b308dfc5013f87823e98d9156301a408d0044b81ebc3e0f5435c06acc8aac6a5dabed754c6da5a84ae4e68e4551516856eefdac48dbd79b8d8f58adbdd79e98d655454533c413378fab566c4f6961c5182039b2da81492;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h698d7be327cd59e1d3f54d6616c587a40397bff9be24e1e410309ddc90c4f6ed6a57db0c007ffb346e73d11477f5655a3203669144e43f46f85c925f776ab9cb734ea8fcf735c8c8b61ea00fc9c87d9761895866b7b2f43cd68c3554ea595d8206d043c2d4c628a9b44db1ea9a79297699ee28dd079ac79649486f9fc7549a63;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb344036b1ac80fd8d14accbc0c5475905edb6903b6af0db5c5c519239c0d5d5d70075f25e1ef15cd2a08511cb89af829899c6d2ff3823b166073947a46df8133e74d88678bd5f6824906595c6d89b96146a98290b36a85b883c67607bea2acc610172d5b54ee440f70b95f674c010139b51a2bad183babc55f19236475cdff10;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27527b7a297cee2aad8aa4643d473f897646aa3fafc86723e8c1b38c6f76c1aa7ebbcbc15658ea28d05a39d468ddd27f9cdbdf90ceb0361978ecfef5563cbc5e846f5cf5f0151e542187abe465eecd39dc142ac7d56773f3e977b9a1c2afed676d147c12d7dd3995457bb4b3ef3be21a1af262ef2120953ec5ae3087ed40ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbd20ca3720d7d81ed8bbb45f2d2a8dbe7c5ba2f7d378c870c863567f49ef766af8eced1dac55795b83bbd88cbf944dcf732aaf52c7440ccc866564a971c8bdd4553ec1ae4ed06d02c597b2bade91ce960c7d882b35ff30af531ddd86ae6a241cc0baf1e3ff0ce2423ba5f225f0572fd8e0326ac994a8328f31db7d244eaf759;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c596d7a17a20a2528ad8ef8f6ed1a7a13c86d7717da271026982243bf5c04ad6ba7f576fab3c3bf70b23bbe3db2be3cb886a8833edcdcb5ac6da8c44e43c354a1b93b8345bcf742ed36eec2fbb2b1b1f9345b0984345202924ac5dcd30fe883492825dd2c3e553c7a189d88c20d38408ab7386015880d7a4bbaba060ad6e46f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h972d8edabb6f7961844df4589ad3ecaea68f2f04980f11c9a69532b7b54a23f86663923b3258bcf10254cd161b9e93e2ec111aad26eb18e4db83ef3043428f12b1da5563047a464961dc6e4b7117343a8c3e4462adbf54432ee938c25a88bf4c988f51169ebcab832e269b6e75dc8457d19a5aec54d6fc6d72edba8f8f3632e9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h492d8b3690c4c78b50ca1ce6f2a5a6b60adb239e05ba796223ae88f034b55b28a836488d3508767379a215007b24c21fce69b63237a11be16335e2130792612081448e92f7429668bacbf5fa48d929396f3b24e5aa0a53001dc9458bd7310b7e1a7cb4b532095225c5680b7308a148146c6777c2bdf82109076badde9910fb05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h166378e3687eac13d6d9e19b0a01c9a21f9ce270e6699cd97185a27b7d86228525cbe38f5edd480605b326d8969d27ccc3cc76f55836054750eb50928d2e3ba9f34c6fa3dd24bcf8ad8a5f2bbbc782d6319e4421a48920dff9316539b4111d5a8e0091a0acdd13ce0a45d7dd792ce033c62449e88335861d320a04c1ca5356f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe4967710e8e0daca50d15896ae3df3a259f9f426e94ae1f0dcbc002dd096c05b0b8ab70754a4e581c3e5acc746b91dd647a4400cb9ab14e6e75806854c60ab2d57ce00bd56c8a453db326f1a512d1a3fca6d045e917f7f27b6a2475ea71549d403d8add92fd8cd07556f9247b7c929217f52a0791e174a4fc86785194aaf4e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc5f6aee123d800da552321ebe3e09aefeb54412f5bf4266c52925f871074623bb5860dde5c8097fba3f78fc9d7dfea73900c315fa2b4c7bd6d511780efd77453e33e2c7eaf78112d347c27260804c629aeef962fd9b07000cac5cc9a34c881d8d5b02079caa5545a97e8c4586a60691804cf5db905e5386553c4df1aed3ef67;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33eab291aa9935d9f981880da677e8d33b0793242e1fc9638f64e96bd0b361c7981fc2f93098141117ec8a83bdb531bab26b82db3442a875f4de0424e23238beff5ed3822e1686b1cddd783302030741dc8559bd4ffcd9c807dade26cb1d0cb495c7ead09ab212689b11553d47eef224aa0b19ff2a37f2dfdcf4524280b00b6b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa88237452ac8cf1f0744989ab0e2544eb074bd1d40f2635d3868b1f2eb038906a0f4f1dc1491bc19a8fc97635bc475f2980bcdc0d12927db7be961d81ce30d0bde13237128d2351f01687e7080691e5bd059adb637e84c71d0ce9f1f22cd1cd157b6e91a4583c973d6a41b7b477b3981c0c32aeb27c013316e863f54fa9c89e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35b00dd0d00114b6ea0bc48ed32aeb05679721779c7c506c48afc2edca5b23e599fd46fd0375b83bb76472317e39fa8f266ad50d0be93c986047d4702841a51f8a46631a053af15fad84bd4c7abf377615adceae81873cbb6e8276f5b49520f63ce1b5aa6338668ba30a342b3d46a66e29d8a7c122a0a4b0701c3de81284e815;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f2ba9237b702856677df19b11a5699dac2d20d9c79c86aa503196efbee898a510de6320eddeae1c8a252996ec60b09ecc1a1f1b49c433d9c085b61f3b1c813ddb91f6b9a99ce4405ff7a6f7c8aebfe42dbc134d03a4816cb38da6360d3c9a64e5ebbac1bb7f6e2b6ff3c404c6eedc0f02120036decd5bf88d80e6aba8852632;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d746096247703ea59fea1e663b0249382508567980cdadb99f9879072b27d16abe2944da619a679316461dd81f92a32d09866a533664547f3fc3150bb0f07cfd805225527c0f00d2dc925ede1504d8603bb7d3eb797d27c91848d4cc2ac02eeb4ce306bb1f12f2df7763b8be550caf4bb988c22d91cc4b1988280677f4508f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99b53ec20b111a968a9068cc7dce3241c61b1dc4c3fdf7e6d71a209daa4920b468b1f4b1c939b9b5829ca6a75cdb14e37d941b9604a430f5c55a8e666c1aaeae15c6c25c81727aa8899cf402fa4d73712b72a8c81aa9d6db60f3d2223e7ad16b9494e9c2671f7962d32bc4896d3d4fc855622e88ea82251fb5706e59d88fccb9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb75b6696cd8318ab09e8101f8d19903bd40e1c34c5736c0b19ebae6d398f6354ff93e0cf704e870a92e50f74e8998f4c8dd6109b13997784c1d9d5d1f150d61f37cbd89f00bb05b27ff0ee7075cb4ded07ab8b5b3f12ea4ad9b6288be921ff850e6e907d2174caf2b992eef76f51c2422ca2862c915111226e24be6c111f2a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21f18b85d59e27ae1f2f1538c9cd4a7b921095f03d5ae8bd004d647ad8bd086d2539bb4f5a1c5fd8413cdcc96e93f04b8d0eced00828db1fc214496ca8d831bc2b420ed319c6307560084c8b58ad530c03bbcde6efc29d8a6be86f8007eb81dc59ac421196541a9036657039ed8a1bc637b4b4ec17d2e1ee6dd0562e3582a0cf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b00f772b5af689e79654b78f65426fd8d762b9fc037f8749d7a50a9df6d667839be06d623c313a36e2c18dbddab85f8fd86e3926084dacce08c9e891568e362ca8104881cb6438c2e51540878d5413250b8afcf2603f947717711f7e9c4b7bcebb4285e436b370fd85ab1948d04c488ec3543757adc079ca00677c48003cc2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7267022e68dd17162012ae8258025e818e0e51ef2e7757ecfcb89c336097c60b0f9f37a00083fc842747d623c871ed896450cccb3d9545ef2f6fc64ce355f6494d6bbf9ae8a2cea58b0509f7cdfdb7132982d78211d45351142a542bc4c01cbf987d5a0c6410b806c0a02ef61cba1416c7cca0f5019ffe677a9ff98c85a366b6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heade48920023c9e2ea2874f612c3c1af9ee519b1d1cbecb133f896e7fd8cfc3a22d784dd2c4623ff9cfd2d2e923914683fa438ad6e17efefd9f6577df2abf81efcc55e261da197ac323b2fd42ac80c8f32eb1bcf79384cc4ab02d97afaf55814f11f22a22cff94f5ef6fbc949b4ab5776c97498b37688bdbc12df1fe5f40e72f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc610fe5c24ba3ac46bf84598f80f9bdc2bc0c470da21a43cb4de2d013433ba4a95d53a409cffeba22c069315ddd4d2c32a2cc32a8784aa6cca5fb6ff732b9986b021a5d1f6015b89e080e3242d0cbe5002b8e72f3e6e5a3889658281ee9e114330fc34e22d5035eee06ccfdff46156ccbd387f33d04ef9decceb25a56acdaa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6484ca9eace340042b910c47bc222a34f4fcd07507a8549673d01a01f134b8990b7e5bcbfcd65d373eb7c8aa08ee2e1d53e96142e1195c30978783f7fed5939cf7222f403bc2daaed4b77e370fb3a03b2edfd68c13ba5ff7e202ab30ba8e6452b984efc98819561cd2c9ac30bc1189599859ddca791f7d3ae46be8b180854019;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc7596169e3f3de00ad4c68679c869be7dfdfa574b1772956beb18c9d84cb6620670995b333f1a9608e7c9297449ace460ce5cb1c71d62f308a66b95e2e321a234a52e5f3f98e07d5886ea1023e078b61a468c8fa6ecc1e71b53e0c7f3ab8aa46295757d2751575886a2807b3538130064a4aab71d8ab7cfce7d9a7f28ba4dd4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6de616397ed39bf1059a4c6d21cb416ec02b676fe0fc56b82d8520abc65d2290364209be67d5bdea9d31f0d3195403d88a6e40a9487a6d8f00676fbebc07f9e2b91055839d240c51971117f44a78d792101435c0e0b5f99e8bcc96e462f040bd6de9eb0262f387654218aa50729f293e9dadcc3d992f5190ee55a2c7a4184a00;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bc54363d56de215f7b35dcc75bf2740fecd0df551283e8fe58c1f2f8c6d4c866c0d1ccb33bc2d9ea2a6850916661dc7f94cb72fdab0c8d704068f10f634835700d82ef6373e0d13626bc0eea12d0ebb373f47a802ff52667c5e860d450a275d22b389d42242fd3c3606b7f68c5b7e7cc630a30351795009f41a3adf6d014778;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae38fc449fa1bdeb47fccd34bd62d88704eb1dcc877512268e78f999a7fee514ff34e79f4503aeea3f80653b8e9ba612fa1b397bf93f40dbbaf106d65750a5a29b8593431c061b87eba3c3bbaccb557a9855090b1e8e24293c91f318e7405a4acd2228fbbe8c8792576ab137b2b955cdbb84eb63a7f0ef41463963b573f5b473;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9b73388850b1049faa0ce9c5bd04947aff4ac8b01f8593701f0e63a17d9fa9cdb63fbc89cd22ed22054d6122493f8da12278c9c6772e560b6a81da3b71508319de69f5bd8761ffcf57ab00a6386faf73f903e9b4dc63070358ee2e509049dc0d06d81ed931dd3e6c9259a3914cf0bd700d12f2bce9643b36c62d362c8d46c16;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a0367215318a9e0948ac71df5fa5dc85cd266b38add50e0003e2dbee929c77024d63cef35e1ee547c5690741ad50125795059f6b2d759a9a0ebde7c00b9ebd8e1542f30ed79cc474d498ede72bf352fb7d69ad2d3ac16fb9b0c4d9ff668ec76199ed5e1266360d9720e877d6a41afe30ed8a75ae172aca053cb0a7a4e8723f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10c2c4cfe30dc0e6b12945d5656b965ded0e31cdc6a849021d2a7d73ca417c94522d439b7ad5c898bd1dbe37ea7d54c1e32f46fb70096527ee1dfded930a8c9c72b0e67b1212ccbb9721f0e0d118d76d63d0f49bbf44f976bba99a33221bc074500c5d3af2be60bbdd10aceca45226fa9d8178737ffe86b830dfaea25725d0b4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefc577e610d20550de2823704b2ef2814aadffae0235c56fb00d3593c04501ade6ced3dec2c9e2a28e345d9311ad929ced4d3575bf2cbde4a2362c57a19f1318e857e0750a1c030e1deebc08997475361a288fc0767db2ffa15ceb4a5256dd3dbae7b733c966154aeb727fe2de7538813b64ed4587a1a0896465bdeec09132f6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f3bd723d10468044f7338e7784b408dc9056c7e597e6bbdec3fe2d0dd8c121c529302b8b861cb3580253b85cfe6eaaaaf479f1e887efffd85f2468e530439e02f3ecad866bfe16e90fac81b233c1c601b8b8a8fa974ad75051915579f8380a8c78beddf36d9b5ce09010fa76d28046a6bfeeffe31322c2896f59e65a60b581c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h221c349e6bf8e8ceacc42b33cb52b50ab30bbb53ad75707cacd3c5623919d486a28c83c36c2e4ec22c6de14128db38b0ddb2dec7534c06d6308f77afcf6e931f358f3afef23e8f0236f9de8aaf5d14b1577c59162ff49126bec7a30a9d0f6d76a9eed6cc0b00bb85b1fdc5934f24c47a6df7b0faa207cb69734b79b772a0596f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7583f5c63c4ebaade9042234dab6beb5d77ef518590c853c8c8a96b9ce070c4e6837d3b1ba6fb2d00c77b9d4f62cdfdd7ca70347f3e766e1e5c1d55e3e837e2fa385f2ae087809b28177314fd43e31c3b46add7dba752000e84b437371329fb9898b9f84e0da39451a3b1028b1ad02004151666848b1d14be1bf1122f989835;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f5e010259344eb9303e27eb403e414918de5520a88a4428ff6193323a225a159e1d97684315044c80c23b86bf4cece19067e8d986944a0421fd48b1c751be8c6ac40d29841af0d4a2834f32cfd36366d5961d2c37a1ec46e5647310e441104a9d7432e49321e3cd289dc13705992348c61a34b0a1c61cb4368e2866f68ac48b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3d73f31961ccad3319554077e0f3a30772fac476ba3dc9bd82ee8d00fbefed824a27f98d5e525abe5ca37fa211e1f6af34fb2cd081c0bc56b62fb8480580de28831f74ee28761b055a3822d43b15cfe48b288eae636c8322a5d6d37f33bd1122140f1c2efb5dc6e61520550c25b5c959943af62d45ad11bc116d71473de36b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h584ce54f52168167a273d44e72985e25e71958b744a4db7e31f817941a070fe306f122637baf5fe83366903c0f2c7c7dc2a4a739eeee8b2543a2dc5016167662b3333e98bf3a76118a23aac2d282c8d477cf093af892e99a555a67788fd8187877969146f2cb1c06d5d68cd266e8b37700b593be99c68a6d67aabd173ad731c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h288c5fbac538d51e1dc17c9bfc6d86f8adb16ab88d13d1569b7f5087f15e5b79aa093dfae89a455723ac495dfa1a60c69dd9a2ed037bf2a2b72d8bfc35f12d9213439a59e55376e9aa947f716f3b4ffd962901e5336048d6d8943688a17805293629a15d263f8f3d2e61537b7674f3bca82f590a1797b5f8554e743c9f9d2b94;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h645da25fdb9f814d8f5b1320eaabf94da89fe25627cc00f2697189377d99e9b5d444a0cb08c30513e3810a4c285763d31c9a3037ebfa4848b1ae69894daa553e5ce45c04edb46c8e56c14d929e29a3080761d13f1a55b2f0d4c1a1720e026c498fe44668938f4f7bcefd442264dfafdc41317f1bd89a20835ba89b10ced04e06;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6204867bb01a5036f8e8c57debaa174f11f917343e20e3d01bf0edb36b532f43639793bf4749a43609f7332aa2f26893111832b0856725041b29f78cff9f407db44e425f2780730cc1a6bc37b963700b2d91fb6dc302eac9c66fc5cb3cff6301778b41781806733b0c4086ab6553b3f783ec3997c887a678b177292a80bca3a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12819c8593c672c8892d3e918fe12a8ffe4541eb8f88260dea429a99ae88701419990a301c0f5bc14566becf3a0a1d120e8d6931b3848686567e0bc8fe7a9b8d0a995adee1c0bb8f090fcb6ac5c1d9f56b07861667f6737bbdb5ae372eac8a8baaaaf62f0dec1c293f90c90e416f90a7f7e2d032e29a0176b490929c6193944e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he58f39af6732dd0518d87e9f0e094934876f3130f8c526944a5f978c4a1c1ef64e2c2869601495409787154f032318c3bf2f27e3c3eada3ce6ef6acead091d76593e60594f3d3a23ff491786751fa35e841103b994b9a595f2296414639a08d45e804b4f85507ccb80aa17adde7892318beb4c6fa0a72e0dc5effeebb108cc44;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2682a4baf8012d7f2e2355d7c82b7d04e206c3102d2a4d32babda918a58ee0a88b5466ac3e1a102b195d9a3084bfd924d671df09183b5f796a2f2fea1e9ec136f5311b3e71a9ce2a287a0053150be353401b4ba807d4b20dc3d3b3cd283fb9d7220f7d8a1f6cb0a90989dc941dee4bddb2ef825ed1863f30eb151a844b4112c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67f3791d5edd68f7a950e66041ab2412131c31fee598172f2b60cbd109b948c99bc8c2e668b4f4bf454ebfcd8c4c5cb1ab8ad0b4463d19be8a7e4e3ac2e7ca67e70b9f683fec7ade2fad85a1601e23568e7371f95ffdddc224e1f015a14912257b1ec04f02dfa0fe2e2cc5978c5033b2d22be84a21d586c16b99a545c18dd06f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6dbfd00df0a398373a3899a26538af0569bd6ea238153e855f5d44ef244be6fb9bf1caec08a2de08cc0be8024a5a3741742e950f42fa99ae93eef4d251ab084f9cd425a966835f81d6c63b13db05061114d467c7b393b3b32fb13e7aa94e002e629419e617350a0763e8e0a70c0b01ebb0704289ad1061f462c0afd038e9ab2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90f80f52dcb4462b82c79fc1a1f5f4d2b8a6ac77f8a318deeb35b2c52059b992b6f4c76983baa8ad6d7b5b5b77848f2dca7f23264f4f74e7f54fbb851d115e4d7d04db45ee132533e5f732b7713e9c939b5a77669618f70d4c333b5af081767cae9dc5ae36d6f2f12f4bb8cbd3592325259e4be746a5c44e49aded2a3b3550b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfeac0e471b09adc67332232317421fd323f7685af6cf109b01fd7096211f6ca0e458e70cd8c74064cd6c8020b2dd52a3b305ccc8caf2bff819337cb89715b8353429d69b6acf147b0f4e20c8d8548d21520d396b23b79b4aa4f2ad161ce3a53c67a26d2275533e34756878e4be5d507fcc1b9323846b93891de6ca6dc2b58044;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2655653be38cc3a977b0867b56c0880d71b2d012e4654e19f0d70f8fd7cc7089b3f41c7a24f193ead9013ac36c849e7391c5cee87562821dc6cc63b5a458f9878091975e240044d080fe4d01ddde995408a78f381df3a14c4d2a51275e54184b118d7e8a1880cf2c472758e5ed60b0e10268b6369e83e8e56262dcc011b1a81c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3b8f3a2087cb36a25460535ca12784022c684b9ca0ec47128cb555400edbdd03cdfe791e10d4b85f3e82e8e87bfc61abe15e712d06588a7b2318764977914b1a54ad88f9ff283dd9c769fcb321c17b80d9dfdd4d6ebc4d7207e81cf88f76273a6c0d4fba19cd65343cca90889a8985798ae8308d790784b9f21f4ea52b6a87c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2cfcafc2470c011756b158ce1e36fe2987e161d9314b9b16e9db3452cd2d659bb5b1e3abffbeed02bb132714108d23ac3143b275dc9cd2d357cdfcbdab25fcfc630bcd219c3ef2b7ab1931a0dc519ea7c22348103b216fa3e9f5bcc3773b96aa097b43bc435be70df6bba24f93c41350b63116ef5562199a3de5a4babe4af829;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h126611a82fbf61938187a643166b42bcaee4e0dc1aafe08a7fb3d246deb28f72cb5482db9324f5ece4f8e51d2d438ebbd606c0ecca7680e24eec6a8a443e25c9b3f9248a76cd7375f2b2ccd19b18690da611ba1da1a1dee29986ead83d36fd854ee3b7748577aae92af00064a3029507f690d0d974846623d208f7d28340628a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h117e20d0b26915d31b6f7cb09358a8ce4eb8e799125df964a514e8ba9144ea0de7b0c63fe10bf798aff052fd542053ed3fd08f8d372d376e552c3705aaca221cfab284786e495595604486399618c9026a160eeb568e27bdc749bb2431bb6dbd9fa60d12794fa1ccfd58c3349a6d61acc7c9e11d3fee14c7c0beb4e5503d7897;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b021b20f913e30310c90638b8f55849444df25ea4a3a23a151f114cb558c0393c2019457c932df985857ac35d6e85ed5239d35b62d4b621547868eb96f3c2078b75dbf353a7072203feeb8b5efaad1d7703f9a3a90ebff2525cc5240641b3169e0e27162addd776ab9451d4af4be5edac2e06e1166eeacd16bfef74931ba334;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb010d1af886c353e9e810f498057c1cfc7683b0ef207d38f4f6f3fafbe5039c4317f705ade9c3e4b6566c030316b2eeefe86cd55d1ce46416d4bd015bd39a9f3e35fd9fab64fd91cf0afca2053b65f61a40f5e3ca11d86d4f6264e143cd7c5f1b7f032ad0a203064e94644d7a3b90aa62e2f69dd4866467e71756c8eccbf6ddc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f6ce50ebeafbd8b234a4ddcdf6f807409654f12e2b96d24b8dfd4c42d423b83dcd05f43368c9cbde4313a13ddaeb303cf4e7d6c99cf81559960fd0a6a8bb70b20a83a21163168f72cf44d1c047e7f1594f45deea66cae58b63c3cb902e20c59f17be4aa0ea52604aaea94088a198cfd746d0d3859c8d1cc21595eb528ddd3d0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67ad048cfcc1edaf27a6ab11537e4f882a74339d47dbb4bd2f28aa2099879f65ecc904180411a1c29884a100b0cd053a07281e15019cc463108fe861823ca22a3a0b8ebd9f45c3043d37441b34abed877b81f92b57078529c7708e6fc50128f8d244fef751274a8af9acad18e865ea45d24152cecb29e5e63c8b1cbbd8973b4d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c3faca1653c420a00140b4834f29636108c45ca96302b935e7f326ee4853a94f3316f9ea748a97c1a18db1506310e0c92321a9ad16ce9194f80036d58a05d5b61c5f09732cd5d4c2f50f20f4ad4265a1dea7981c1fcd72309e12cd02103d15825f1f66fa2a0bb37b7aa29146046daa6e714cae2d140e8fb62a63629c3564ea9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9c1f22c5219f0c4e36bb8da82f9270be287cfb381d558f7fdf686188682ad2f748e8b3fab7c40b97e84d691e44553b27f8d8e6d4aedfc79fdbc496518e7e4ad191de7d658b17d8016b725daf9b18bc38c2a3ab1921d28cad719b40db7eea491c2a1693c79a1f3ac7e4e490f53c30f0f4017f7880c23d84882b4113e1fc53c7c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59dec54c1db8d8cdde0f619a328cc109303cbfff048fe945397eb77cce20217d474a65d1d9c3d475fa4e3aebc9840cc3f64df235a95360ddcff20ef1ab370307de422b613d99c1cddacd5a524a704b71e85e42279152e023901fa3e8fec2222cffcb76903d917a4972c09177039f07699ce51590ae0e1dc0f02c17d32c15f581;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f1824b7a995727ddaae95d2935b7b5a02e9afe0d885e51a3b63561541ba68788d349a9c6956f66115c4ae52378bc638536dcbd439ec704072e73e2301b7020d5ffa7b8a283704997e87ea64ffbaede9b61224ecddde46b1f56d9390777c785380159dedecac9942c6c85f35c18b275c95d9c8978c592ef5791bdb9f4668770c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce0809c8ccee86a5f28b0af6f2170bcddd615166404e27eef7826f7150dc91ad9409075f430ebe2bf1728119635eb285729d7bfaa98fa594d09fbf333aaaf5f0e8ceecdf3bec0fa9fb0887b2af777ced77407b26b53ed656d3a221beaa64abed7a0902cca8a6021bf0d4db2ce871338c5230221c33e566e556f3558e85874e7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62e2bf70fc4ccefe907ef073145d16d4eb50493dbb430c357d4eb27431397dd9877a6a7996a9dfd1d178f4f5ae39d9004be2665afdc0341d4163e6d52b0453fbb383a70136fc539296dc3e352a2ae14b43b6ce0a4442b5e3167bf88999e67e810fbb7853397c3099957ae9909caf31c3b25f160159ace195340cf81747be858c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h248afb895b2c73bfb96e6fc68d0fb12db706a6fa71578182c7d1098dc089278d84c46a80fc27f1cfc3140a321863dbad9e1285cd392e1d6fb1f980fec0acf04698d32c556f3a6c1ad22a20af8fb852746dc401ca2bc768b437d30437406b36b3f644b8f0fefe941b63df92ea5907df2f7b11bd9e6c9e0f92679ac7808da743df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12fc54691dcd1beb4a21ce324585f259ab4a3f790d708b0eeb21a898094d2d9f79ee646c8f12a6079001b8885dd917e9f83139b2c69f83ec9c1d66aabf7aedb28594b35370034ffecf7a6e865aa3f2c8fa9bb05a408f088d65839f8f0ee64ffda11f11146f91afb3be3cdaa39ee903bfaff9a87086e6b8292cc74e881faec2c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h136959c9988cdf39d5861112abbfc114c127468932da78a77163f3a9a17e62a5042df5489c8e8db0f7aa10c0947dc3ec28eb989cb3eb91d2a83f198bbaef789080c026729977ecdbf1b1bcdfa214e3bc27434d6e215d6583d3b4b8255e49a6af65d661a2b0e3d53e442d4e2a0624841baca29d0198c7f41cc7f546edcf68961;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1a847fe23f9f1009edded73408d3891d6f5edaa3e79da9e6fb38f0f40dc80338b73226daecfe95e87e6afc6e91dcf9daa38d1e3d8914362791ea61bd5db4b38a88a19ff2cf36b31ebb86762e77416f90915df684bbbc1ed4a945e8db92c0760160a8f35d36cc162bfa91f3bf03c3e87845d07188edbe5a491776136f00a62c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce4c03f542284796a9cbf38596e74551cdffb1a7a7ce991ac10a3a660d013c244badaedf2ef48c5680c8e157b0027af3f4ca1d1403e04771681607f118e4c4ed3f87d8fde1fc76a51d8843b1745597190debb245ea9d188ed19748a0b334464721064fcc1d720524335682184550eaf20886d89a61b60a4d2941a58a310d99df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd31a2aee2df860127fa79f9e4f9be370792bfb50c8dbdf1a25b48d7dcec58c6d76032887511008a21660ed3730f952e44ab0ec0037eebeb2c419391ee8168fba9d28a5df0454975ccfe911f70b6dfa31bed31562a0e8f75ea6a51d1bc768ac052e22b9e1103ca2b84fa06907bb008ffbdc0947c6d487ceb965c39ed6c0650aae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc80e086f206ab51dbddcd2aad308786fbcfdf47b6f004d669d53de18988c6b0bc13216940636c3bb193cdf85285651aaecd0eea6d2a326370fb3f9d9a3a5df8356c2b1b4022d96bc320cca8a17b12fa35aad02c23a3fc9a905dbe6b42514ff8610603b3c5f8258b1d5655fb1a44497ab565db520ca0cb1881d4eba71867186c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haac5276841fc0f02dba9144b418a695ac4b3ad73e9499074c01fad0d744029fcab0da6853806092aecd1991a60a7760254bae1f5a1ad943b6b11af0089ef0c4778d575475ab8b53b5fd91ac57bc0cee2a155cdf507716a5e46fe75d1824077303e42957ec7a8a1516cac078441f719044225a0da1ff100b004f403d80c610f34;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d3d86c60d88b27cad607403b3a074b9f5387db9dd5aa61c528393e4c15c67f935d98f47d6ad29ec41f9c99a3eddcc89c0d2951f0ef4f6b37702a98630d2936f4043587e9a8e139654390d02de1473ca384c2a9338553d7a570c08b4c4b92a8d7021a28be213223fefeb00282170171d1c0818ac5a36d4ed9a500f6b57455688;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h177e7b55c506b7b6fd17b38dc4990191781fc41db9affb42f5615f513f597f8c269a0a24290cad6961d410b937f69a91d059a04a172553265347d0bbef9bb7a929dd958542db2ab0206f0a701b2ddffe880ee8ff4ee67eda9ac811d5653f8943edd877a1d305e2cef9ce3a368908ab55938d4b944ff4e1d3f11215553c97d74e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7f293e84547dc4cb3b56aefc0edf15bde1d10005725d7cb9e8a18a2cdf6c24cb02f601376d61bba60e73c5d01867ee64d95f83fbd77ff4a872616473d4004295b2af84e0b8b2cd1a58c3ac0cb3668d8d36dd444ef56acd4bb2f926ea850ea6b7977f04a0d8b6193ecd306412af4cb5ca639fec352a86159304a556c312901b2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6338e86eb823dd8262ea4483e749a237d7d226859eb9dc12df4407935d0298e7512be2a3f578f3d16f798a6bfb92e39fea9f824368f07003abb0ed2b5378794bae880625f8ecb302be79fe8f145dca53b1d25e34f844da99771b7f79cca457a29c37f0480bf35e196d553914e45398b430577a7d930c1ef995d4e6ea96422885;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbcb2677459bd837918a362677030c5e26d913280d8b7b5ff9b40f4886abfb010f8095b10070d0ef08c7cc678c46a279408378dd72f9804b2ed4dd01422fdbe1e9537c35e78fcb6709726c7eda860e43053716fddc920bceb0831cf46e488bb68e34c04dd792d8c26632299dd7d6eb1f4d06a0716fe9904b68f283f97bfd908a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc25a91da9d6d78ff3e8bd68fc7d63b44598d8bea871ecc97ae9ac4b9bb93883e1c7c996e40673affdfe911f723e0df40f8cb51b9d33f04801ccaa7e589a4f7532b5511438ffc8f9cbdfaac4b22b0fda7d2af4950b120c6f5c8776ea04b90ca4f0393f9390ae6e2a3b2806f983f33e1f181e17a3250ff77d05d93840f046771e2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf3b866bd1e48e199ba2e04922fc6ba3fbf0ecafca2c285114f0a0861b1a9cbf556222183261dc736b13a725ecf675bb78be0b9bfa8d7aa6dba17c6af529c9569a951c4fcbbb5369dae4d2de06934ceb20c78de866ca96537f7d971f7c94fb2d2eb62d0d03679f7de2c347ee68d07dc8d50a06319ff81a28c47fded4002c8780;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2b285894dc45ab9724e0e645bbb13da7dc076d6929144357df8b6534e324662ef2ba76d0c0b9d76417dfcf3fd426516e1910bc111f8ed2ba021092c91d03ae6b149a8df8b4d12ef202851cc8667823501035b7c3c8db34598654b0ed7026b67e1c19115bd57db43044459522193ae12041a69197d2609f997828f5bc8601fa9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h291e9da46dde9e0d4ead3036b211e9744b5edb1c76d858279c396dad9815fead6b4180e130ba9f1a514b12829d0e2b95f88127931e38c3326f72ec0f2ce89db10c95abf74aa3c35e8d97bde03406f92701f4d3770723382c79b118b9df9f96c8e04f5986b5ac83f726c71d1ebeb18cade00630c2eee5c34cc7978a7f635fbb77;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85d424bc0f9031b9869572b5a5eed1621f4177e38e3c9621537ae65d90fed4d1ebc81bd98a6818508288621bf858231195c64925968963dfba3514e5403ca7a83ee76e7b6b8ba622c0b440a0ec0e4d0ca202b55df508a2b34c4306282d3b5aa24b76081bd9ce76ddb852f1c8da42859a72a0b3e79aa99558318f17665cd85f9f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18a14f094b744bd387e298540f5ce9cb6743089a619597a4665a42dc5eeb3c72735e1a55c2ee2597cd6e05494aed91faf6ef3690a4f5a44020bc27cb979bee0703b3c9bdef7f76148a69ecdf09d9eafeb1689fc86b5e78a86faa524ddc950ec6bd40edeef0758c9efcd20f3fef949da42204cba391f8f1c0dad18d49debf966;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bf143d75088df70a0f65f68d441adf6754704a42869ebeb404f1eaff3ac97a0866a8f190e834650580e2551f7bd5246f1bf472d61bada38894291a8d365e722c06bc05ad2c618e14a955a94568e8a00be4ba3400e88dd6893fed3022cedd5a70634bebdf26e3f781d8ad4a5cc27a767b09c2f8e216aaf711159f40d4cdcf560;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9781f02b057d6b65ba7a9ccbc2555e7505dc5c18d690ee656dbcce960c3053675e38e281e2382a82ef81e007ba728fd0b46b03238854aa341605e37e00cbcb1b71170f919dd3517f36b6d58211d665190eb2cd4ef60d70f60170272c49bf67934e7c98eb380dacdfc6845507e9a952438fd471cbb4d09c26c5b916a35b42949a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafe5f1732ce7788ad8f1ce3059383f144e1f950d300368dace1fc316163f906f8f2e81fb34de59184b226a8259a9f25c1cde5159e1d220799fed3b39c8ffc4f27ee5078989d7a9c379c08b169c1d3c1518f931bee5983e7fa51218d85d1a69032d7eb644351bb977f5c02a13f07e300c47bd0cab19b7ebfb8733c8a38ebf7d5c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h902989667e0d65538dce7441709dce1b0d9004154338dd2e9286e0dafb4b47721a2a37ca0b279f329f8389141571fb2580c7dca370c43c06816060fa9a17175011256be1c219de5bc685360b38c7a425ea4745974ee7caed3385b190206e77ddc391d09000b5adc0d46bd257e129feccdaddd04c5d1a63eac02ae56dfce60512;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2c4953091e435a7dc750f9d8e49a7d857e29c3c968afd6b4d18e1c5f30cad3d121c46bf61c70e612be5160a832eb924eefd330dd2d408ffa8ebab2ed1495c27f328b08d7263a260797d3d4561c3ed964b21df8a7bdd891f66d57d5ec6216127887d99b964906ab9247a5dfd77e872ba5dfdd4a8077ea3f8f5d6832e8b196cf6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4fab405e92de6afd38e153cedd146a0cdc6c7ebe44af627ac5153a5b18abd6909665db97b313a9e8619e04b4f098b458e157632ef1b03b84eea8f68d583612019b52046358e8dc0a7f874b105c5ec9d39f2ff3625b7b84aff6f42f2ce1166e5ed08db75e3d759318e983dadf3b1f2a80e69e18f49efd6d8bda76d2ee6cec0e0f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had3bba145de75ccafae9b4e2d7a8ea45c09fedb2b5469db6af6783d84b3ff3cc97446c3427025730b2b6414003076b11b28ea863a922c3845e25836af41b3a0ce791566f021dd978b9a127a340a6fe09b82ff3349cd4df20eed1d738d8aa0bb1613731723aaae907b69fb75b6d7286e011d07df7526ea97029716f86a5849262;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13cfefcdcd9842c5e937b176e174cc4178df8667dca3bf166c84ebd2e55bc8a9e27db54e7b64084c4cf7989983615ffdf6a397a08b165ed4e4364be9ca59ad9fda56d8d065b51a7a2d96c5905c156c833325fca58e127c41a4cf99b799e3bf5714e3ee3a2361a376830bed5839ed9370d2a6d12c984f9ee8cdaf5636e9430873;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60c7705970ca577eae78669681e205d7cb2aef0f74cac2a739abf099037cb30cec2f5beeb190d35539f2855b6211d2bff2cbf742775ee1d5c60f0a28fd81b3b49aa442a0ad1c8a08a65768bcf4a79a8a69b5803bd0c07d80a25030054f7dfecac867ed5bc1b9e462c3c46a0c2830d03ccc69bed4ec6bad98f3183535f69c9395;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89d81f48953129307ce2c183f569dd4c13b8c5825ffbee2be1fc1b80e01c850c1639bb463e6c936fabee1ce5e4d5045bdc0d6394ac517078eabfabeff4993c2d297c8ac3eb893cb5d275b50392ab7cfe3605f38583fc8b1cf2274d5aa05b7580025b0bbdd12ebf3dabc7a270a8ba7beb32fa321e9548efb025bafd8fc3ced29a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96abfc75c08940296109c06fe3fa3a31439a9f6bdac707f24d923ce927e728f8d952d8d681c49456de756c10faddd42e2c832e3d2af59608d1640455d4c30faf3a339c5ca170c5a90a3410c6a614e43921c8a8331efe649b72b1b1e0d053945c5978bf033b9c8e0e55fcb141ea1d6f6c6265a231415f46a9ddcacca304c4713e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h675442098c794bdfc57222fcb6fb34c183e25b8c9b6789f55b8615039c0e2216db263ab6ec7d9d7b64a498cdd9d0a0c260d82f52a4e2ddb8b639eb808e6ac37cc051c38c5f769f746532071b90f8c89e80b6794d52f9b7d95313ddb5d3bd411401d1bd829fc631a421a5e30fb49bdf345bc40f622ff15388e5d05baac2c23937;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf32f62dedcf2df332051c43bff16cda1ba53b3caa91fe71711b8cadb6344fe12add12394c8d4896806b028ace79757139e35678809fc3f7f4f3eb468db1b1954e081e5b382fb360d54864f663ab712278bfd897f22a102c7307a1b0d58c9701479f7a99bfb73dcc106bdb334ca9406af4beefe5aee6649914b5f1698d3fc976f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1b70cca3052d06e6ecf6c656e2c549ea5bba99a33523a39979dce2ff3038f75539b28908fbda238b95ba1fcc0ca59adc37ef7ccd0f87466eff148cb57791c06bbe18b30a98d900ea3edd2ca93efb529c443cdaaaa4826d7364e1d937bf7a8cab0ff868b4f1023dfc18d251ed2edc105a8ddc75383eef1046ea3eab4814d12d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17e1b4e09f5382e821bfec8f071447e8943c625328f61f935fe56d5050200a9bfb1fa51866271fc8315a7635274aecf14034316e738de0c63f301c919913708c2b4f40279acadc972c7e9dd2db5e8a0232b688d61e4eb90fdb5f28c454d07ae766cb23ba410700d2889694a8b1d4f8191523d9a440bb7af5d7f73963ac75beaf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47efbdeffcd714dca6d03212e2faebe3836dd8494d8432f77708de0c9c4c017ebe7c2a3faf2ed86e05951a6d339ea143fb47cb0cde860bcd778ba7932d913ff6c8a95da5b371c8deebf013b58383d5fa8016d341476624e07200e240feed6d86114198feba7b8e9605c96b4eb524e43795645733f4280704db84ce6042d5fff9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb0a92a4475f9ea436127edc78e625dd17db95cf66788f7b44a9ed3bdcec49135ad5f683b8ec78ea1d4dc5680929a587e9fea7ee12bda9e0dca2c84efc87d3d0a44cb6738c94f20c339027139be2aafdf4c10f9d953ac037a34c0b9ce6fa71155e943387de638ded2e0cf69a77a1a0b49f2dc616c16e5652418427e056adc288;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h950934764a960a658889d5bc9ef8e9cb77828d309bd4fd373faadc334c342cec3e76860298aaaecfa117b072373e4064c79c6c64a9c950465c01fec3392da17a5ebe3fdf88c9a96a53e48eeb9ff28d6e7bfb7e2630c08aa046d830a0037743cda6ae0aff49759afd555fbee7e92cbd0f40269a44ee5c71bb7dc5cd9a272a0701;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h525fd4a5055cecb9fd3f38ea8d1b0388a800d4d8fb3d631a23e37dc576f1a2d6f9b18185fc38a6cc90582c44a0f55c431ecbfec71165383f70bbcdfe0ea8bca3b2c0da95a7abe8223895077a39555f83e920f274227e5f2adcac01c9c85622f7836f9ea562288251622e5e4b56faedfece7e8699c94c490428905b42ad0396f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e982217a016b5ea6cba330344eec018e82f09750adaaf4ae09a7abe2b9d5ab95aaab13f52c5e87e84318bcf5588564b559d245725d717002320f61e7f7e7947427c6209d02f70eac0894ac25801e0749eaeeb1eb2f81652d8f1530d2ccd6b5d80debb22f9e9f65f496009d56b36ec325181feeddc929dd29e82a65a653abd29;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3bd92d877798de20f0b86f60913646d55aaf906b723dcbea36e3256c8987b3ee111704b673a3123ebef19e53d4b23422f4ea83f930c08086fbdbabc4da1774e8b699a01ef11c5003183c8fdd1fe3da20e9a69a2bb377eba35ea315761543f45035f577bde9f5e84424343eed426e79f3b444ff1f30531882cdbac6d3ec036fd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82e7cfe2c2827b2638a73bc29f1aaf69dc8bb053e67dff6ae839debec7e587c7bfe83bd9472cb910dd48e77f4d34f8b9938fd4f2ad6127b2267ab9513ea47787097f074a7505bb3a999bf40c7c46d422e23183b48bdd4b658164a660d015792a752fe3ea29e76de0cfc0f0a45404aaaffafa4c24e3636487bc2fbad0c78dcb87;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h161ed954a4b6d26eab093dce6b01027cc7a1ce91ff57fed11eb5176874b806082336a142ba1a11c968a57f4e4190500945db1e24955ad5b4ace022c50e0863788085123bac8e72da845546d35b0ccf3e74efe715cf92816f7cf79185f3bfdc898b6f3b3d708ef46bffabf08cbfaf794295fc3941228c7fa43f6536c04f45d72f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79a740ab60bc188d1e2d864ac3ce590a8a1c5fd58905770d2e2e3943de7b3c05de53748bc16703fa1b5756c32257c7b4b18a27758139db78b9165af4934e9874c0df4f333ebcb681502d31871ba33156a5a42938ed6e9bb926317f326df7ba3139270ef168b9316525347ab40069566780b2f7dfccb3e3b89f5b06b0b25259e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2457b907875907ea4367df758768e08307528723ea22d8242fd5447656cb4f9f2cc45fc4bea9ea5ee5ceb559fd65f1104bc3de9bfd22e591d349e944576529b2c3116a35cf6fe2c6ff05dc56e51ca36f266bdcc32909f2d6f389b54a2a662a4f83c08c608e8dd02568c89728f8de6c5a732bc681a282b598f24e28e2d97fd1ba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd39f7803d43154ecc6217d033781a346bb67c0a94e4d0f32966391ed026cfbf104b248bcef767d533de031083dbd164dd67c7cbe388dabbe0426d5c2d7880f466c31776aec83c6025390bf6248abc6f46d59e1078d5f917c5cecf875c512d3e0789b9bacb89c483415d661c5e66708500cc0bb15e1113c217ea2519bbb31e372;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95909f6f5555b57f4e0cd8bf4a0502eee9a27b8fcd43de963af6987293e2f748be457cb501ac5a0c3f86dff05920757e14335fdbccc71a4d60a76f90ce64da5a43d52d31a306d6c7ec5f0ab1e5fb179fc04f7382a9b2c4a3e30f12fdb278ce16b508aee1dac004c1b5b0c61943cef48183a6638781a2d7db7682c7bb2ee5d85f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1d24ccae3a5dc0eb0aa7d86dd06a562e8d6eb80404e27e73018f9171b419fddf7aebca6192d4a382901ff7d904cfb9a27c53d7d0d06483451a782576e1599f54ad46527c2c3c2aba8b888b0fe5a61e89b0f95699960a1afae1c1c290c0a3a6e6b2825c0cdad1c758eec8d5595606c3bd340f5f0d2c7d4e787a5d2552fdf77e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h232497607380639219955672ec5eb7822d6d3681020262d430c2fa5a8f9233dabd70aa84542e067a35884ba89c794901af956e4bbf9d9a27964be56bb873d1b717f98bb1be2c61c4b078114c6d7fe5d03d8e2e6c86a1659ecb31861adfc6ff2a7718e0044c6a0cea237bfc389ed0b9c27947607199880c08372baa3970889eef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e6531d8d36ed56bfbdfe520686fda2bfe9cecf90314e943042f9a21bab91dd3f9206c0164cb5a0d6463752b3cc10767a561685b24fb2b2a948dce24d11227f238e6e99c956b2edeebf0f57c54e24efc06d2ebab87a57607dbfb5603005cba9eee837c9de169e6286b661362a02cf8d43efb108e9ccfb9407655d8010c07e976;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd4055d9ab1d6f8c3d9aed7752c11cc0ab562c734d02d1d82230e74a4b381f0d863dd1bf486e857e1ede66855ad7192c36e31559942de42eec88296812a281ec36154f1639fe50a44547df8ce0878f35eeb6ef4ef5f70ff5ffd0472c6b96c4d902efd06032cc3169241c7cafdfbeb0a7dea41c4617fdeea0bf8808f6ed6ef7ba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d35cbf6ee63ba571f9a78b4666a33afaa9d0d182547a5c0f374d2a2377f82149f6f3b240f0040fc53106d46987b10eed387a2da8579a5ce5d7affd5cc4bda50bdaa497b48fa3741e024066707fd4fc5fd1475e3094539e457adf0a5102810f400122d89456d1d851a435d388b9300d1309e4394a221bd2fee12107697a9c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he342e4852ea8cfee944fe21c01b34b2cec2b627a50f16689ece671f1b189c02aba6c165057cc9cca1c51c2a0c2a8ad14307ed64c8b723afc122b69165c3c79fb3d18bf5e317cb09251ecfc1b423cdd4fc34771a3b9705d58f56c94ea335ea1fa72b8ef2261e3bbb32021814663736e9b37b36361843d45f9695ce64a38b37b89;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cc1f778dcc2f97df5d85c5eae028be0c0a77fd99a60d830882cceaa6e0bae4600caa0be7a18ceade23f068c5eaedb1afc48a2ddf4199d042ee642a4a483a3d66e714023b8d137c9b9d029f2cc9a5446feefaec57eca109fec42a71b29ddac04865050f4d39a4b54e549d446ad93d2b4a4202cdc9bb2c478d2b40075461c780f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39f0d23ad0275ad083557c47c265aa955f01b6f361c9e47b662ab191e8fc04dc67912182661876101dab7b3a5cf5017518df14b64799501eed9d546cfec226bfd0c2ecaa04b8b4b49846b7b3e5ed1e9fe33aa591604770cdbb63d51b05e5501bcdc7c54f5bfab0c592fe6265d6c302225f8927d39afc3a4d382919e94f20defa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h355fd4a3cbc5ea943987fee800b748368d2cdf1a8e14cbfc5883f381c8d4994176fc5fb7d7c9678a5cb925873c7b719fbaf13618a872d2f45264a9721327654593d8c35a25554c0bc57c6afa8669d1cb694ef2da4666e28422af2dd692a694ef184c73f3346415c5a85b11342941e9441c7d5fe1d3ea00e944b7552038b36834;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f61eaed98b49c90684d8185b17c1ea5b7fc35a24ab5f553cac6701cb71a01fca78ac8e3b8e8f66790e2544d35f7ba80a2c218053b111d8b859edf35d09b768bed87acfdb3ed03d60d948a77b787f9f4c2b8a4ca6529a90c97183d44118f91fde5c79c43907f6027b9404bd69259c501ba3fbf781116ffc478f489a4132ef547;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ba1deb666b2ebc7607f7481e7d3737cb5573bfe3aa5c56e7d52f5217a7ab0c4aaeaa95af528bc65ba8ab4bc247b5af973976644f9fe0d018154a510031ac82866ac2a952f61bbde71e9a5143063d5fda0a41afa56586dd2121483123889a63fc28dbfe65b24a3927884859f93783c26c8b5b3d919e3dcbf4fb471052e8ae05a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd10f275b0db3c6541c22907addf61cd241b08960bac81b32e3d9e9c0684e847b2d9d38be1b2e4c9f153440ac47f44a3a2524b7e5b60da9db008ea7c6fba763d0188d0ee2aaf04e55570631bdafb45058c3a6032f9c3c05056810dce6f0fae6314788d1c27d3090b2ccb9c71422caa486eed94ae242b4498314cd381924151a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h851ffc8a33a93a3710282c4196cf85f67f91d6a9d594a5ef272be70432cb7c1fe0448aa0bf1c7b4684d4f504619ef41094e2ed780cea69c1ae9390538a43169248d5e15ec5692214b4b24a8703083036eb9672860c60107aeff5edec4ad222024adec38044717d4ed4e12039e20e8be80763087655cbb2670fd2dbb4f75dfd5a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h962a75bb0f69fd70a46b4a72d0a1d1120ad7e2e9e88ea95fa8a1be82bc762d9768eec053a009294718a63863bb87b9acb925a032b549646b4c9ed4b89721ef25b43551c02b041605be637d61602c8d2300c730a2dce8e8ca2de11f7ccc262b02f5373e0708aa4795c8cd91d1ec9d617e49d72f8ea3f07b5a7750391db56b1f71;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7ff0ab5949cd8562ef91d48b15fba7126cc7fd831dfaaa25d39a3191f3bf7ccc6f0b9cad388446e8aaccf77fe2b97609c58eceaadac7a1df1a3f2de9c270e69f53d299e4fb2226c0be35c8ab267228e16c620cb2c791a63169968315cd8c9d5d73c5516e6dead9d660f55c8f7ccd5f064edecf14a1ea322568fc346b6e2b04b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e9727860411fe22c844ea6c616219bee84a26e0df8ea4432aac98961be80a029b6b343f2ca44b532140adc5902ae98cc4854e314c2de0a91aeb7f92b4adf49a531c4e91aadb3a2269307b1122724d1c37c9388d0b03a98b2a8b80957d1bb0091ce67dbb3e866f50cb694119694dde214de8826704755cd33b1ad08f993a8663;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ad118d01e9822caed9f81ec69f4e3f0182a36bf1dd0a87820f05c4618df67337fb14629231a965df38b69c2dc272bd046168797485c1b9ee5092b12101677d79f893414cb734594d3aa93e814f35815cdf889bb49ca5398d248d1dd7434da9302ef4d8abc49886f0407cd164b15959218891987e02c9c90a6609a5713fa32ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d655242bef09844b67328f6bb33621284a57fc0d3c011fba0b332e62cefd258a773f326ec53da612da808425d34b26b661cf872bd6d002c8a540dce0bf94c89fe479bf520a9f9df4f05f86aeee42c32de73aab6cf74852099a8712ea3a983566c11a004883c3f143e802dceb39a0342713a99c5d36e6689defd712050aea24b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa931f21a6269458adf6e004af309cc4a5a05eef38b23c12e032b931976ce0dfe5b6017a882372d8804142568e1b7630d294a870f29a6fbcbb0497a0c1b4ab5e79f2dfa32d019286e3e0927f4c8a5f7122d994c3af7ca1807f86e3ebb6ea21ac9ff4888a3b9706bed839f683e87be55b2fd18b7bc168058efbef9dce4c0ff832;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65e404e4bf0d26e7585f07eff1f3f7ab87ef3494b86f1b127b30f1c33538c09bfab26b1c7855a540128db1793c617f9512245a04dc9e808ca45b3694f86a28c4b911cf12ed815863c0b9ab65cf738a30381fa2ee560c71dfc15b6e2fd7e2650a70debffef658042bd93195c9baccfc3b3639675dd2c7fcbda54daa134b0a2a6f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7da603a955cd0c79af8d52d868c7c00d9b99dfd4a770d466c17ed4dff04683ead50319d5c76cb6c55133b1ed812b0d7764a67ef82c2e6fdad04e4b6a19cfa45a516990b78e18cdb1dc71683b4fb9e320f0a21c11256a26acd72234e0b4446a0500d17c8b22ee654194e5f1459cd2a4becab5990ad92e39a5ca57e82744054c1f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4bf0d905f650ff1715318d6ec1e3ca69993fcd8734e0511ab1befe5376325f4a1fed34c832aac6cf5157860621dbfa1edf3f37ad79c047c50cdd944062519697adcb57132d96e83ee0e3dd787c83c16ef6b79db32d1764a15445c2ad038b1ea5818deef19b52dc41318e1b477f4cf96cbe22557762a1b10290ae07ee3c2e0e34;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58b89a7a4e0ef47225225e71e83802a96227d10beb9ba55e3c3f3ca57f8cbaef3f210bf3aa348576a674822380d937f2e99ca3a76aa3d306ffd4e98dfe589e04e8202d57779316755e987d49d154f81077d0fb8a784c6ddc499d5d382ed165b10535c146a8825dfc2156d13351440a8d7368aaae6fa35714acf1492efb8f1a4b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heec2285ff94f82e21725c80db0130b38fcfc387cb46a88c29b3f3c6a7dc9790e255147a10be5cd7fdd4b35bc28512913136724d78e5c5bf24d74e2bdf4f2f3c7c1552ea6701ed1bbf355ddc967c4a7391895ec6e594234270b6fff94d69afc26c5221ec902664e571bfe38c4b19c5b8cfc8ee2bdbeb226eb32d83b25703f7ee2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44625e28e7ec731efedc86dbdc94fd6892eb487498f2e488158fd749163881d8e19901b63b5d9adf5a69cced404fed672b1e2a401be0d250fe890d4a7898cc3c1050ed90b8e029d45360effa379bb69e47169ae6d4d067c877cc4de78ed99e6bb7514f42e5727622729f215b955201eb0726a9566a5213f299806f30ce80a9b4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b0c1aba3f03608e1bf3d78b9c1ce704ab107a06a848ea2d9f95c73d64795a9a18a6aa99d822dcc4ab09ff5010afd1a0b80eff9ac8da9cf87a4f4cfd0f563b87741b68674ee01562b478a978893b9496f620d2ea9be3a2e1db1052c5d8610ceaeee3f7e41cb494957b93fc7f84c7f3a7ba17cea3b19e11509bf70d487a53be1c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb907f8bfc1c06707446649f4937f24e4022ec42782e243b4f98e0153930b1ec470c44165c8b549d4f8f92adad9d698eaed243c52417b16281d238596cd3aad357453339f7998888d170cb94ff58d605127dbde14101c72d6ddf2a81a68de14e6a3c0927af9e320e2f83b93cf365019f877e9341053948d025f78c8e5d1efe60;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a24825f7c01692e13bfb5c061d5e0afaf978ba8686c11a463c569d6dba23bcea37b361682efdf5c35e1c27439e482d6dd083ae9c4f67c8bde131dc58790e71d851111cdae00d94a54564a34faadffd7912ab3a9442c7b6816a53d0e1f3a7275b9b7dd043ba687e2508837b4be5fca7a01114a516c14151f9473a24dfdd077c6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4702cc0576aa0f3564d0595b295ced50584caca006f28bcdff17ae856d2a8daa26bc88a05e09aa5e0121a6eeaa025bf97ba98e8d242c82e4a0cb729b160116b9f0eeeecb96be0649918cd962f3673645ac8475ac069a96d52fc13bdddafb9c19e2f6edba707fbaebdd3538d38457bf7243cebf64965cec9d80ece544e63de307;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habd8ac6b4da8239582958a0bcd45f0f25be3e9314889cbfb45d296605e8fa13a2a355ca8088a36ecb3e538e58aefc8b0c27d167b8d20d585792cff41cf77395dbcdc55f8639a5c1923b57950db723fa2b05cc15f1f92de9721576a265881d75c367447aa49289cb23fc325177425de83bb89eab44a9dc0686ccf87496de83d67;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76f74aa9bdeffdfeb7d9c934081c738a457e19c3b029e0d1c4dbc4c29d30bd327d9d16ddbcfe3a611f17ecee2576d9a65008ffb8200e488bfb6556dbfdd55c77d03683dc69f107ce7729a6f54960ad9727f0f8dace1acf0c4b7a686334e6f6d2d0d8af0a9e9640a4e1eea16ce6d2a22a71210b084b452a58f9baa195f7c1e65a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3b30011ec6834a921b8497f820ea8e0eed082d6f8ac193f0f08801694b3b9896d43846108479c0da82d96c01050a3454ecab3521e8935f5f73dfb0ea56e68374db9b9a66bddf19fcbdb25da4700b85b3f8f2cf8a6d4fa6f9718a30dcf411703d434d0e4a4b7b45682a6d009d2e7e65bd19b0b9b64a9c2823d93e12bdb089224;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha662386993ff7aea3c395c40ac8864df72c5049d1e63ba2186ff1bef042e4a0c2993574e93c7e569129de22529f15d3cacdc1fd868bf588de5dfb85ade8b16b2ed37162bf363571c487a3d7c824ab82b4e3fd2b4f57b8bcc623a880764dbf62ed370a6a611bd58daa71cc881fde01811e7e8f33e996832c314966322df8f619c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10ebb307c59e5600362ed9301cee4eb3f2378adda2c9391b7938d35d6f0089b4933d239dd0296463d4052c548b789a879aecb7304b7b82c660770539e26488e259e37aad554ccc355e4b57dcd5b3c285fb1cc13500c6d24871e98812717d3e0ed15c81ee42113ed0bab3902a9f9e67a648a0732e8730b42169927bc636ec46c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfaf43ddde1edeb62b97379c664f111b979b975a66e144a13e4bb70f20092e6bff9c7afefe88769266ff6c60eda25f91d36ea9f99a94e37946bece8875c8f9bcd6dc1806a1af65e16b35ed8625dbbfdef89292e5b5a0cf523d612f3847154ac3228dc8b0f256ce735d69ef7772e833649aa7051602a5a7b0b0d7bfdc23fe0bd9e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40a2d8ee2a73e4920f23e02e95c937ae83def0507ecf076af3e6ed0f55008c37d8bf9d887cadf3a7edb50561ea40bff934ac4e7ab558a238486c37e3886398d34e35cc9463c39320f48f625da5204546d1fc8c93890c1150763bb865fb58b207739cc524bde916ea9c5626ec898d11c92e45379b5d873061ab67cde33ae14c54;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3937d9d464a0b7b32991c508f291ce0df689cf6fa8e4bdb1bd52a65277985c98723f462ba01f7f8e62fe3b8f56d630c8185876221eece0a0a7d988fe6fa1c8d4dcc14dbf489f6be59ad5337882215e61bc2dbd27d3e2df86c79d2e9190a3de961515905046ed1a884bcc4c15db22d4742b2955feba7b18c1f5444c3fe92cce00;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d786c9cf5c283edef369df615bf4456f3763aa2fd8445baf4735f784269735f926b048a45bb0b1e9eb6bfd4163dcd3a2f069e238aae438881cbe257e456dd60cb6fa5b142cad08565afcdbddd690ef021832e6e3859aa8c26098d84650743a134bce594efbdde4eb8304ee1ab34a22a978b8bd48f6750d577b46455e4eba04d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h645dab314a42601c0417a6e25c498ea6eaf20931063a6cf59b2de0fe4b79c8ab13bad16ac92ac22cf5ae161e8433aac93d562827fb55bb2b9fc29a724176ed18124f1cf0309efd2be8bedefcc9ee1bc21b2d3c14db6f6af2f4b89cb62fd4a969bcc214732b3e5a11ed256cc9f50aa6eaeabe5bfbd36c98fb9501318baa4ec131;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88a192faccd386d8298ca55602afb28fff23d0f3bdb39edf32ebd9b389ebf70a69ce8de02d58f64d99c29ee93cb969118c0a0df91a55132ed9f60b8abd59f27e249787c122a69f3ff1ab09adc4ebdcd6efc111735e6dd8d5638ae4ec50fc1808b1d6ecef1d19c1bdc511670b4bd1ae15214e95e50bde01936593a004d8236148;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h162f17d19f5f49c61f383ec128651c032de7ba544d224fd11692825c4ef21cc4ae33cf04a9967aa3ab452a74e58d3a4ebf27ee430f09497d9776bd57f1f1f68214d5dd38d95b272a62f79825c6bff458139d43fa091c153b40b9ddc9e24be922a3a18335bb581034df95d2d41d31fd806170952281c83da7f2f89c451cac4a7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba7b7a19ba88e8d481affd874d80027d908a8597bd1c154ee720b480127581445aa74d7b7ec446c4be6693fd427d1ccd11e093d93cc15766c1450618e2624e7aecb9e8ebfe2673cbae77faad1b049a44b3fdbe6660d3d8e200a5725ddb1d294cb4c764badf8d88f42ea5f3f3b83deaf3cfdd0ae108b13a7de901c35f73e1f226;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b808050ebb1456bdf69de2093fd1f6dd9a69b544cb1390817a9712394e41a993584cde366a61803fe229ec93472bd69efffbefaff143e31d93d54d9f9feeb1b9c22eafeddd06448b2ca422cd444be2c27692ffb628192ca3396894de28e7dc0eb981838789f28d8b97f8f247833adee086bf99edb0b48d2ec2087f057298eaa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h808e461a30d74de652c2a0ca2ce304a31d48e1f71989f897f3cb02464b52dc013d21e442e8e8dd03f7e50953a8a6ed02d64ed491f8dc0922e6019af5c6ad707ceff77d76add3476da978e48939e07faf10516f94f67a07bc1958244ea7ba0146664d1314b14bfe713346a37a8ba77d3e7dd4f55b64bc6da9375dde813f6262c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd29c32eadb9d58bed6c8651b19d42bdd4d2bb1afad8113552e0c7f7785d48c262012945baac914a72a7c3b3d5f7055963231f3fd1c6629b0b33d6c375d7564f429799f14dbcc0cf17817824dea793debbb7d2f1b5be89aa9a01633485cf4be0400344bc2694d329765a7cc7f5fa8dc7489a815c98554c84819ac64fc7a8b1ca5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3d20cc36f097750528999e7ea336759954bc14e2b8f2ca2ed764902bbdb2e4ee3d380906daf2be3c1416fe3fd829bc9486d821333dbb38355e80254e57df0f113177c91322cac74c4fe9443c90d5203bbad601f79a321a670f957133c89ac97965e537438cf35024aa451a0d8698e785b88ff7534ba7233ad93a467bdf562a4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67ffbef97085a523793beb281f58836f676d1392fd6bcd11b63c0b3824aeb7bbc750590da0419a364d53b673db797ef329b267a1dbbb2a4e770f8ebbfb670c66e27adc4a07585f015661c6794a6a38099aa46252c15147fd486fded68b9c8993a2ebacd35c1851f58c27c5a14f5d3747734de7d82f52539c612b39102147a84e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h403171186242653dc1e9c36788abc3d6ea9b9367891ccada06ac3afde98ce6df3776471e1be31509014671a6814df03fdfae2fe6da76e30cda188ff5048e2c970c971c077b7c273ba1662d6c1d90d053dd621e955b61e0bb21cb9ad555cc607b2742c80296e681d5d108287d5a6a6f7c9114150906f2156860b50e81052b43c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h77ae275112fb726b2279694c25720038b89bb5cc4a9d901c8f0432ae2be1adf8b2a2c2544eb4628e7d71db48cc062e5191b470cf9ba8aba74a9174e5687df6dd58fff202d0601336228397813b2624e36b52f77d2d1d38a51968e2084b9fc6e4391b91e733aeb436583cf286d66a2d8ba41432aea0a345a12376eb77b360ddb2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55ddb17f6ff9a4543dd727547aff24341ddca993439cb50cb6e8ca622a5c32b05cf30e5a47dda20d532138b5d23f6dd9e6106506088dab26c5eaee264a0e97825d37009a5811446103d755aee1aa9985a47a7b8a5aabec2ec6228ed19539469773d30cf18c6c0935bf507015cca58040a83ca17153e7f08c356853c678a7a7fc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cf1910ced302ebda57f1f9c52ffdf908a67f8c6407680f50725e125c1e6c7cac356b2d9f1ad747a454712a436cde5fa51ef41098cf5894e9de150eca6e5eb8816eef2e722d1451d825de6fefc96cf4c7c5566b975a434bc17e42c3c4cdc207efa9fe06761b8466827ef8a20881d35c6dc6bb942877e41457ff4fc411b8bb004;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d829da6cbfcee267285da8cb40c7781b27d7358ff4254cd85db3341266a17425e5c77609ac63ad8962dce42f8dba2e5769ba64ebc436c566ce371f4aacd023a5a940d3ca7f88ede634a9e3e6157af7cfa9c3510a0fd979427a7dbff3af2cf42e59eb6cc8f42eb76d62aea0c8d5b607d4188f86e5d7eb310bf3cdcb1e3e746ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he82f39c3c378b1088d4992c180f83441c8d94e11bdb94cfa03718e2cda8ef0513b14169181b083e10641b237b897d9dc4dfe9cf805d2c887785000230585af5f70423e7056f1f3e36f258dd00ca9538c40179cfd32d7da1aab0e04afaba52e4a146137964fc8345b83c41ac23ae6faefc78d900c53b74a1637ccdc62c1f3f5df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h279e32096e75254072023eca7c0e5e86d4e5b59272cf412c011c3ca138652b7d7dffbf4b5951ddb4c5e88a313736085417b77e99b188e05d9c4f16ae848a590895fad21e27802c1e55fd32bc41ac1a52ff21c08ea70abf3b99967ec21aa4d11420f65ec42ca8303448a409e6398f5558e33d56c8db0c08a1f6777569e4345524;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44f531cfb4cb472579a4d23688f3b2e286a415b4795abe57e62443878ab635838dbd6343be3108f6121357d718183fe709f28782ca5c8ad4fca3dc705795c4c5a3156316f5a5663f1dfe2e87f53403aadddbfd31bcc0f6fc0d05cb3c7ec8e2bb3d0e016b020df4d55ab2f7fbecedeb7fad6c15e75a4499e7d908bcc5b76eb107;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d55982be035b149518c80d261a2d4fe0c1d40205731290a3f14d2b967b888f86bc87c24de4b2323de5c027c645fd610c40d538a7731c135e96766758a409f2a8826fd734d1ca556acc7bd58e21399580a745a26e9b575898ae97c8c2a8355b596fd86c994b67809fdbafcd178ea90766025a962806e7a1e387efed5833693eb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h281da1821eabe3c4532af09f4d540a4c24d6810308ec429b7817459ea4f089824f10fa2422a5e1891a251a2e9ba093377811af010fcada1e45e2c177679c6062877b22b3305bef41b6abaab4c1aa3cb51a24a8d5f40b7d6036e763964affb762d386a38a0c761ba510949a65085ec8af1c494e99bc50386a5615414bad62952d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c5f556e89bd630f31e31e302c40aae98528e4187e5d020d0d86c8b7466ef2ad1d347ae1c2ec571e26bbfa290b9ae9215059ef9515c1d4ea7872a9de1caec9761e3101e12ac9ea2550ad13d184dc7e6ff930a5f7fbcce12e877f6c8e1262e36804368f929252dd65338c174708dc700ecccf7374b14b75953d01edacf734f003;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb81a2c744f5485c0fc02740ea536879d11f48e3c6c24625fc6ebe62ca31e85c82d6c033cd92a71e8167022430ac5207cc69b3026b8fd4d91db80776e4166483594adfc94be77896cb6c96dacd4b0aaef44a8d18bb5331817c4a5c28297f11effa0fff78c0058025623ab70f83da2ab8ac33878188d82691fea82a781315e9b6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h373318fb4f13b2e994b86b299591ae4b7e89db64e799498227bd599c6551dfec7146f4289d4b7f7025afe3ccd1fda5901dd080fbc61088ee1bdd44aab40d6bd2459a7c8eb99d12eaa0d2696403a799fa9177315b093b22a4a9a17503d6a6bb7076d58d6ea653380e837166c0999296d539c8ae80baab880fb36f8ffd0f9d30c5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb37467e3c87f4f6137e7d1fa80026e1ae9614d666a3ecbe2ebdb763cc455ac5ce4979e41430bacdcb213faf1343fd4fa55540c232629a769d9963471e87538a483bcd74c0badeb44fd5b76e864537bfa95961e54fb1218a5f0d037e3adf29107b7ba9eb33993c8899827399ebb87235b258f5e6ed7fbbfa4580c228a1d93d948;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8c11077f3d167b50f83f2adda3cce52d70f4483bd0e0440ac7164be8827c8a4a824f313a901b12b31487bd2f0fde47caa8bca8870760c86cdbe21e43ccad8515e03a5fcccbbc19b87c0637ad605928c9748bec3a5bfafd493db73ce606fa854a70347ac873a56185f0eb8727de1b73f868d530de4dfa5ebe2d7f7c7349b7cca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc090a2e03f87ad96602709f2b3097bef77157a05d1e57731602b926f35174b5ec00b9705f2f83552f0ca09d8b77e0be80f4e149825a0e6761c7099815806c20fd5abbe78531373ed9c01865cc12a65e397166f192dff54e9f29ee08e035e2a5187031315b88e744e668e16dac91d125325ee9a51bda773aa2e56c70a4098138;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd861794c6f224e6b42465b18f1e2e9c6e3e6320cd2d3a27db04862326d21e8d7efed055e3f60d6e5ccb943a01f78e7482415a29156fcc078d1fdb0d08caaf5f039fa7b8321d8662afc8e74f00d17a9377d9010313765601d83e3ef4922f6acb5a134841b19cf98a31ef747f4129fec3b881677640689325ae0d0adca92b1b503;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82360e3ae81a4874312fb020fe206e83ca2a116bd7cb1bc9bd1bdb97164cb345e3eec4529af522ebbe78a851e1b39501efcf252b4245c5db317cb6b73014354e443d324c92c256c7659dd8ff8ef1322d4c9b4a57c9e52f1a99ca2551c1be13af06ba29605bfa2156450aca0142e85a12e7dc4ad791a73662c1ccae9d8f6d9d30;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc20c0deca5002f7c9a849bab8d70b728c7af88a033e5a37445fde028c33beae3523eb5a584596d168fa696024393acb708694f88424ecdf6566c2a7012f2b57230cf9ac28d824798266361ea82ab22a8678b3efd41c9e0cfd460f9b6e80881aca1224593f16a6ddf4bdd2432af98e60b4d0ff656e19bd426f0676b9e2c78451;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2dcbefd334f2748cff04d009a7d98c1c4dd8f8f0a59fa709b69cc2d68e30406bf22feb0716ac2100a30dea50b684a83f0d68ab0a22b85352b8125f2b6695e919a64709366768a14c29e4d9d47a0c989ed8c6cd2509e09a7bb7d6925ac2a77d5080d148418089758131d87a715aeb00140fc0a2d1a98dfe1481c95c194be1e2c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2d193a54005fa8c807ec17aa2ffc4e6d9d66f8e06d8cb0308c1741edb85fa897779856755736d4b301a3155b2ee52f285a0882d92c3bcb643bb0cc9662ab10e940c5ae7062c9b0129b64e836612741d0d2de96dd073c93431204b932af1e99e0b5fced88a31c95a16b1f18a93ddd2d49ca6adaadf20cd3e45ba5db2475d7dd5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68e3e66506e1f9d9a135e25d0e814a35990a81a30bb6c3dcb248ebcf33ea08127dc215afac18646b8e6d62da2a182cd31da6bad0339b3fba27e958b5508afea503cfdc5b0bb3ed4ecb55598f935c208d22e6b7f10ffa1ea6591f868b62e0eae25d8e37aec517a9b1d7a0e20a93ef47dc23b9c9860e923239c6ba1dc941f10b7a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde9e327d71ef7a146b04d9a1b83a151c12f82b6dcced16f75898e860e191253f26fcc51edb54d99ae1e14cb008eaa02c895fb703b35e2f8e707029480d12bd24eb8a30e871f27da0dafb1c4896947357b918d94c0614bb7f5ffbe4eb8fcacf1568c13ad0a7af404a6cf08fc072dcd2e1e3d16009bf26d7d367b3a22204217fd8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74e3eb2f5444451733c42d6b6b030765112688f7b11ab6c99882d2600b9951c8ecaaf3fad0b67efca704851cedb7332723c555cfc7591bbb5a36d72d3a93efc99985df0ade79769ad75c40f2a81c82eec8c12186b172fc949b31e9771fcc09197c9395e8086e642120d1e7b0f83fc7428626b05b13d1ab6137b364a9f6d6c146;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h157ca60b5dddb596f195905a1d5733d3d1c0baf2ecf4111c6c1398abf25eeaedf37f90152e05051b540a3459baaf57c531666a1b9112eebecbbbb092b21b6cc5e50d7912bf6659eff2e554b8b8e10869288dc23246a24fd985f18e58a256954d9b57573fae7c9975e7ca7da30253c63aed53cc04b826ad5c46f99bd205c07ab4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6fd2bb6eceab4d586895a234e96a661ea9ba9ccc3de2ceb9592d6cb4bc5e2c843107c211a4167258170d4d3d4f2b62287b129811142119ace103b09a08485ece4529201c4faf4dd2445d8a9bca8ffe1836b24b49a94ec1e3f924a1ca836629c2104a29e57e388888a5c9cb6c118e397b736edf8775d8b90d5b959135bf7c18a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf70cd180a05f7945c20d8465f4adfcdebf1d1f85d8c327a24188cb608f628f2e5bf2e2f96ae0711437fdad4fe38cece01e43df9fcaec08c76992f4c53f6b7ff8a8c9b33b55ca6c71acd48ca5ad16d127d255393d1578f572a61706c69e8ace4e445f80212dabfccf37115f68cb1262fbf6f301f87df8e4831ace1c34dae8a3b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b3e99ef6c86451bcacf4f57dc4ac57186063c8485c78684a6c2bb9f3c53f3762d5f8cbaf1ff34a90a4a8b07eda46f0b1cd896af1c89d2eb699fbbc946b96a499e8f5a0475dd151612a43400885f2d9e293c9b14bd2ed92e1393c911dd717f833b9b44facd78e851fb2d59bffeda160559e0444e5ab5bb16069be4e17fbe0cf9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5c37b00e41dc6358af42f5c985cbf8c33c4084cc72503de23554ccba03f32f5a87abe9aad64bfbb05b4da3d905ccb36117f5a9d53be8aa9b2aeccf8be4e72128bd0cf00afe9effd8c16fc7b899549ac8e5268088e8a4088bb72ff99d0e680209d1e461be47cfb7c2f566ff62888838594f93910b0886439232277283cf7273e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3374f598bdee027d11d763c7bf09a72810202b1b393f299ef623fcbf61ab338a4d15db497567fd8d4fb16fe28503b9357c04168748dc5437e67aea0b6361881b69c5687893c718ad4a072a852c83c71e7fd92f97dadb6a9a8bb3beeeabdf6a3ee2059cece01e63e0896a44dd571ed1d25c57aa3822b6282f877a9ad2a0650f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fe3885c43e995ced40519b9dacb06b1283bd8ff1e89b3e92dbd9918bf275f8e84a5aa911a3a3fc2f9f79a16092c3a0d3c49427cbb694c238a08b44c17d8a8a00537a4bc76fc17befa41fe25c326bf9455a7fae5dfcead59deff10db544e253400a71c941752b5747b71767d1181a87f27a6a2f618bbbcb9fa178d487f326023;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd689e1fcdc56b133db19d194e7c383c2033f592dee400ff0d02b31276f19b0aa2ec4fecb39f7ce81e6ad276bb70997269b059d222a0f355657501862460bbf8777637c3bcc1323f4520a273014975c16c40c902af0319869fd37f5e31afb2597d8a158deef23bc733373041a03ca3c6de49123dfc71b11e4cff4e089c14328d9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60f4a0d6c0ac2ce56c10d709de0757bfd95bef551c2977fd64be7c725c566a8b7cf2ab2202598d6db1b9e932887335454044cf8fc5511999b075a8004ad95e521f8e40659521318405ebed904441f9824a015ab3223e78f6d4ad53ed3c54a51d72b405a87a434ba196dbec36b9e7d662d88b2e8e855d2bb0e5274dab7ed2f209;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h965ecaf9392269f2c8e5087121874aa023c415685560c9bfc1fc5acd91b55e48dbaf852fc5f3e40fcc7a071a1dd45d97fcf5b1c65cd465eb3585806fcf5bd3171a0bef6c57dcb7f2b7db4c8069e8fd99419d8ec42d0eb7fef086ff7d05cc51154116f5bd0b2617dfe441a365c68f08eed37ac37e1e5e4091a91d2e36dbe1d311;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83ba4c7ca669a3526da302ccf284219f3055892b76c70f2d12125d9ea9820e8dc6f60541778cf121f999e854a64461ec90ebd0b9ef75a5eacdebfcda5e0dcbc08f7833d2c57445a9aa024ca38024c1123b977cdffc960aeb3c16db478eb9c3f12ca5c9d7fb092f12737070a5ba3ad4d0fd3f796b644a99c406a495b6a6872c68;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b75bd39ec121df68d0a041a5ae7b809fdc3852a3b00ed6550e5954a5785a968276ace2ba7013067368f2ac9a20d6fa9a7bbe566a568fd3bbe7033ef5dd834753ac72c65b4beeeb705ad4194e5faf9c9732a67c0e3427e3f39d3fe270e9ea221dd92c36aefb11030686c9342f252f57ea0da47fcaba1cbdf15e3fe7a6d2dcd46;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c17893f74c0c184fb76819748a5971e6bb9b5acb1cb5ab04195f2cca3811724678aac3a185364f94b49b9e6f8232fbe60b1a0a2159a8822d6fa94ed9a4b1b35cffc38f5a48956a17cb449ad96ebe03d1bb0161986d5521561d19c8ff04a22cb1d0669cea4eed94a2fc1c72a3457e8e6b332f4d07dea55ef1829d11c5ae3d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e0e3ed763289d1b2e21cfcec96e52ecd34e699d17a47b4f87f2805907c01e3e10779a6c47e8cfe0b61306da878f5431e042d15c45bc8184a38cc086a4070266ff5c889d9a96b815ace597ec1adeb2ff2365e184a521c5fc604fb6d108c4bbe8ac831b5532ce0dd2bd2a5ff1989c209e33eaa9fa86c1fd346d4b32492e3efeac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5dec8c5fa75161af277074c2563ddff013522441a9f2600bd1c4dc9e77cd221b3db0d42a80de306b32955c215380e468bf2c8d53a66c2aee1c7163f86d900bde265275a11f592c806e0cd06bc21e1bdc6bfae2c4970248afbdcafd9960acab50ee33fc5d48678598d285801b387d882f390439e063675d382a7f181abd261a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2689d2eac92d108642e15a582fe6e05a29eda140ce649244186a33160f8dacf45576133dabd65a320e4c18cd374f09204c006a0969dfb47b88d001e31ceb3860bfe65be55c331e6b123f2527cf15c4de4dcfdf40a65fec0dfe9d0daf8062fa7781bfa415c6b92f6024a97570426208b7fd079e97bc0f6087a49bc19ba8e2c31d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc65ba058dc36ed69988b2418b99dda45562a51fe7f232965537138184f5a4668cf5a2cde8e1f4d938db145e10703c3161e6d6b7dc6a90bbea9f014d875afb9bce8100f6f2e6875a3f89d6d2c10f8885b550002209a812209e8da60e59d468e3eae98576419cbc96ee3594723ce934a4d315f45f60e176754950d4ed65a6713b4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb13883b297d374aaed3dd2da9c0792ad8023ef29e0ac6f137cb66e3a4c4ece4de93a5d4deb75b5d67f967d28634414c6dad5542d88b597359c2ce1e5353d9cdd0ba48aef4ff53ce650cf2f815a1ee4ca6344cfefebe49a69d00b3c0e97c53cd843ad859997d285a118f965df18e5674afd5b4ccf2d56fbecad8ba30b2238e81;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39d14d45ea8e4408f4b54b7c8ce8d0362bb280a3401af9b70263581c1ae57e0ed1f23d740e35bed33ed7f6c2b9d51d682416d37092a4af22928318c3c9318e47ef88996eed9468b2b9e0aea854f0dea97c13928a7fb79ad3b9f7cdcba41ca99b92b9ac491883cf1d748555fe30887d6bdedf5f1907562741b1607621781867de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h661721a969c9e93b554e3ee29999c5f7b7c816098d92a94c4f3255bd47471b98e0cb28ec51f2e7cd986f227cb95565b43f5431b4751035f203efe39bde5c35d9de9e184e4ee1c9e38cd41260878a8752a50280cae46f3e4237b2291d2506a9df43be576282c4ccbc29b5a052299f6e8510baca768cf6a4d178b6b38c6b95b062;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2f70ad2992b747103013b413ba598d985afe9ebca1f4d078a46d556d8e71da8b011729d50f4f9fa8ca1f0b3fb38491ea89fe49ba7c28d8155074421496e0a035f1bd58eb2a0a4aaf4b8f96b2984a9d36d6a06594c29f03c20fe76b0e233ed0f26174acf299c40add76d0bea30b02cf2ce1ec361315c340e549bc97815d6b302;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h783894e3b1bfa97cee47e6d959059b97d8f00f00045c21c3fb8a7b74e6e7e38af825b3d00cba0d11027f9022850d7fb098e4d3c052636ad6323ea137665d3054cf32996e1e356fe95301cdd4611bcdd072c68db02a24a4353036e2b98e4f1724ead8859a0a46e9c630d79a0fdf477ab45fa010ad582439fb10ce9e6373e7ac2c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he212e1b57a2ebd705e33d83f3bf28ef789f615351107d21622f8f7ae37e2988b80b26da14649aaf81e58bff6372a7205fd683a3cac33786f811cc52cecc22bb60301d35f7c3a47a53c76f80d883bdffb6be31b3b511c1704c695f3a36a5d897c3bafb342bcd0abb89da647702434c478ba2cc51dfa86e88cadae10be85a8a1c9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he202a567085a8ab37df572e226ff9be85e923ade160359a5bdaa6a6d9975a433c0e399e986372587c58618dd89d67b5458d346ef7853f53b8f15ecce098f38762d0092293700ab448e404ea350ee780755873f8867ace8aabf31e49743aaba7dbbaffd847a074bafa94612856b140e7fd3d1da8dfb781012ed2bcb339d9901dd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66920e52257075969126169f217966797d00ab8f6451fcf59a2ffe995c441c52f3b478310e239f7358dd9c9d5043b5774cd925d9347895229b3637cce3e168396fce0034098e7a604602bf92ea84d49c6fcfea76953c9c4c9aa9dcd5a4da10eb2d00f66dfff8e3fdbfd039ad006aa828a9fd1dc1e633ad71bed4b117b3f54703;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26e5de48e0824e6e5228e9e7f2be306da7d40dc3e872fda45a94e48c475ab13c73bab0631eb1e1bfe0360a446689ef050741a293f6d155b197b0dfba2d31ec515d5b51f740812ac3b42ffaccf552d54900431d7947c08aa199107c978c14bfe40468465128ecc7e6d1ee9eaa92d1eb6c8d66162484d6c40ae5bb4a3a460426e7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he546e03d1d5e998286fa563ac447762c4fc28ea432dc0a51778ea374ba93be655a11bd44b45e111043684eb844689391a77050c5a3f9c5b2af7c1a235a585819bb021f43013600508398a2bffa915c4cc9817d39c6015f6ae4b3fd22a5664ded5692ea985d4303ef3a6bf7636f7aee67d301cf862edea12d33f4c627aa94b662;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e9f55985899a4d336b8aecb984176e933f9bacb57a502863b0393a7aaa82cac4fe991ca31b4553bdc231d4a70c50f1e38359b9731cb44352e6a05731cf75f258afc7697c085003809b173eba4544cadc47ffd4cee455ce6be4a29d6b617ddcd7b7aad3771a1db6e3b8c907ef453fc91653aab4846522b937c60a23a9db08f17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb8037b4be649d3588b41bb1b2fb7b8a377b72c5d7c7c91dd5eb4f9548504122ec17e3de9ff912f8d104629cf7f584f53c1085a176a67db820b4daa87e9ff53014db6f1d9b3c68f583a4a08a9b52bd38c23fc10f4c4c9663cd32b0c30ffda7c6b159c24336d732fb69e77902569fadc4633b3b5e40df72d3854548ec0f175b69;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f5f3e9f4530187b32a7e9ef764fb45234cf7fc27184c36d71e8058bfee57f495b610e2d193cdeab2505ad8e644c70115bca69ef4c7ee729b2f22a9edbef18921913038efee632d4912b9171119521f8ddfb5172b8d6996903d5172c37f7f925282fb79634d04cee4b37436ae4732d19fa3dec3f05fba764df3b0bc32c7ca460;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf375fbff76458e5500a6cea9bbe4e8213db37fcce1a311c97e15db807266df4bfcbfc904cc44839037f3306c6dda8072340056cce1e0a57b670cf30992a8775ad1ec8d151bd8088b41f51a4a2afff386ed6a103fdb97ee9592ee63f7d77ff9cd09395ad4146e4367fc15a8cbcdff2c4abc4e7efce528ea9a30ba5834fbccc69a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60bd7661286786332d09fccb961f10ba646f8513900e27d1c0ee9a406e4b3621676460ce08d06ab6a794b0f38d8b6a24317beff21c47ade456ff167678a76d44e7942a785edd3a77d4e0c1f6fc630a1e60d903db4c32f71fbf4f4dee273af63d04569254d0cc98cc535e74cad72b4b688f5ebaadea4eaa57945c55db71b883ee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56773a9134eb9af4c5a1e73e8369e8db409b69e8410c802d8065cbd88834191da441fa7bc71b1b759b8bec910eb2234a29e6cdee29a3ae47907bc3b3a2328a6c88495dce499199b54e94b24cc80d8dc04727eafb74ec72141114e9c94f879ba5c78abebfce36c09faa6ef258cefd4e93ae93b5ece5f7ec40e5a8b6af2984ff56;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdad0317c704f6162e529fc08f3fb0ff3919ef6a6e1045f9f99e0c9f00b501ca4810937448bc89bc65bd03ac65877121ed57eafac25dd5bdee5df0b575d50e54eb291627367b7e90f8193181152bbd9018b2517e71719a1eb9832cea974b79340ead1d45ffc55d73488d590becff7dfb92a9a6ea9967291c976872ca3a72ad81;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9288cfcaa85c98704e255c53235bee7ac80259f141e97d325d933e2a2d9c11f7ac9c2924b9690ce63d51c3f68f40cefec45fc69829bb28859965fb93ca2ee9a4f046da9f433e9d202593550342543d1a629fe2bf88cc85d05f5f5fcae4e84ab4279b31a48c407bcb33338ac33afc371c444136ecdb5d324e2bc97884e28a94e1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9ec1f5f2ce69800cacc032fa38e02274f448c8c21815100fe7a3c56d7c1ddfb95061e59e3989f0bbdac695c8d3170f4bcc02b78db0a4ab1836210ee6759e01ec863f484d7a2383e30672e42de03bb8386ecfb6ea024d569f63e1e3f7105f5525e6e239d0343c2706f6cfc9ef04e9d53b9af815fb005028be1c77bfdeb51a2ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3affab82aeabb2ab7f8676c58421bb9b740e0162d804a718821bee271d30d947dbedf0425f8eba08aade4c3767cb330fa4cee112c204044de703890a05a1ce30234c626c7278757d4231ae103bab37855501167f4ca71a303353111a6a4f4a2947755f8f48d9b93080a418bb01961aac3caf312e256d4d28b03042595ca02569;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5b1054f179aca98bd324dcea7e58c56f8273f7d3e17084eaf44804a4454c499d5e1c566e5dd405859d972ccccd7f62d63eabab16efaa94c70f9c2cc180e5580b5abe5fcb50fe4909d7cf0a3dcd0f1fedb279cd35a50980373f52205b0ae4057c2b87dff3c9035de1235b75450cec1cfb9e4ca7bd1f6e76d10fb4d2ac4f64ec8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2615c5c455966169b86f51242312a84b5478fe0bdd7e47319f723ec712958f24562ac1b067877ecef8f6315eb182c7db385c518565220637d09529f0688cd8f41d7ff63b42c9884c5e3497639e9b1982fdc44c7729a8da207aa1de5ccf8d604265f537beadcde72d8f3092e7306c58bb537f14a2580613a85203211c91386dc5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf928ca171041afc196813e5a7a9d23fd30096b9dcaf597a212dc2d94396e49832688d0cfd8441c6cd4d098f7386e22b16cf70b667e967a180c9b1c38d07fe8b426bb10f998fe8bc0216ded142b408c33a6339e78ab034ff2139324ba8e46190955b7a425e6140e93390c22d5be5a9a2b3b901b1bdd27202397f13380a737ca4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h781d80a921c201c72e0ee2e652854f286e0ff6501946945f0a324af0e5e7e277c12e75cfa7c731ae1002dee6e9944392348511275aef1bbb43c964668368da7d6a6fb8c50c094ca61822eef470c8dda8e196188cfb2a3062af5e1f59fc5c5594aff88d7273e467a2d6d15b267f1141707385d3a710005487ba30184eb04f8a17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfca2136171822a0bdbd31d8dbbfc274db85d5f4ae730d138e3e07afda59cc853a1e1be5826146391bd435399c879619ba474435bd237030f083306bf7d2bcb97521e9648f9caef1ee0d00eaefc160fff7b7105e9f9aee9bd0d867dfb8a85b26f03b5123180abe5ee96f8cbeabeb62942d787197204ae0fd5502833087c77bed3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85a71ad4ac1682cb4a143ac840c1d1ed1e0d6a6df3185eeb0bcb154a9d4995b4779a0780859010035e697c7380a6da264c5a8e8de42188f0996425147062fbbd955927dacfab434eebc0a0d9fe98c02d669d27b8750b348a546cbfbd88bba63580125c3ed276daedbbfc6ebef0379a11fccf0ba1991d55f33d7299d57fe69b1a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93e023548965caa7d7e2aae5d1d5752985e443110dac42053c38c252d411fc3862d8be3ad3e9d3b72ff0dd75e57bf4cc96bd8a07ace6268df3e724a00acc1b12dede3758db78aa01f7872ef4c33155cdfe8af70ec8d6b6fa1df90376066b9a7765ef44b78af65077f574151ad90c2e5a29a95bde557a59e65643f9209f3cbefb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7ed747665897aed3943847c4ca658e9eb023c0c37ef4756ac7216f4fd536e0ff3dbf18c26e5d944c8491227ab18b1e537e4569e70ed3299ac0b0f56d82939a6bc10a83318c6efc19976c93f0c0cf4ee8581d9a67d9002950adf1faaa8f753995f9892adeeaa53ac3dabc7a344ffb38069c2bf8bd2af2fd578f2fd6bb0ba61;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3aecf05b8d8bc6fbe0172b94949535c63c62f510a282da98087efdf560c9143af9ae14b66df6b63b81bbe846d28a5bd331d7c5235548d3edef4d7db5d853326c712adbafaa30fc82ebf04972525b352cb042a0c7445fc7be70fd57dc2f300db43d82cbe6b662b20c8c109e163c86dc3f3c0ee5256ecf89c00d7345e1b5677013;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2259dc7a169fa6936ffb71ca710a6ab1f2c903e12cfd421396bcb3f280b8cee29e56892df721e750b0bc4c9ae7e18ac8758c207143e8edd9e052adb03d094b0a8f9642e3e98fd637ae1f5f390662d87bbc1e2b96bc5e379a61104341635f20811fe775ffebd5dc8be4c2c383e25b7969edea19995cdbabf142050459f4ce64a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89b706421b75a80d28ee85a164b9d43104a640f78508c1523ba854e5f145de7504be48fda2d022d7c30513805ef5aa814d85d5a58a06f9e36837b4ebf16408c757d3adfe54566365d9a327d90e08b278653fe977df45c1d7d1449bd565c4e63e5c7785d586392190d6a75dd0a18fff8454e7efb30b04d65120ce47aa9bf164cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31fb9f9eead5e245bfcbfd40754189cf33afe90a1d27b1f65efb2e7cf5865e3cd178e1b2f4bb1e88173ce01e20b86ec6ff3c05c10bf26bed8020a71c5213643beaaaf811051d00ec0702da2f9f39ecb63f05d0cf64d5e306e227ed4f52dffbd89301d1b09eb6ff8668ae334b56a439f667508c22f871a752c6e93e67e9e40a52;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c579304e84ea7892f056a4b17cccbbefd0fc474ea5bfa68c00e06f4b1775c59d60f00fc78902103ac27333fac3cc7f4f73fd6e831f815025ab533318d3a10f83134cf16eed38cbe1fe63179e06cd3b8f8b7598efddbad63b0bdefbcffd2f4020853340c886810576c0ff97a900611fd99ca05201feff3575ee6bacb8e30269c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcca7c302a87a26d28b42b3cf8ea6d778e47c53b771a070f37b21f6f2ee1bae7a93a9a618ffe1a7637871ada8e9180fecf2a78d69ef1440d6eb98f9587ff6382b855b14c741f680ac47de35b53893838c975dcc1af12c91cbe980c73262ffeef63cef45a895d491c3e792e36e64e6e3ee65adac8ddb34971da118ee43bcb6424c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdcfaa9e4b0eee00ba9246e01bf52a8285eda29653841d49ec4727a8a7f0c455222f9c0d0f538d6dda0ba3efee8b2dade4f84156ca5092bb8c5f751623cbe861fcd0f65f5e32ec536b98e5e26da5fe17c566e68eef0a8bc2a901d5d41fa85d1b46f6c68dfbeb4cd859c118e1730b7565488b85a8feea0bc9ad4b5748cde611a9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h175e8eb4a29ad923c53550606e94559b45f33b528ab850dd17c997162af7ff20721807ef0da086a08347b106845f42d44144a7f6f1cca2560e00c11ad89798061ce59d834afd8bcc307f60f332631e7323c98467f22d961958c8a919c18feb3db7aa932d690d20cf50ad744e7795fb0425d7176345da4fc5fbb1f217e2d4a75a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h655407d6c795582c6864dc0b896400bb62202278884110f01359b04d9453a69af5453c97ecfded8ffe3eecb393d85f3c852c5c7b4e5a8965936cf25d910f5ee9959c7299b99766d423cfcc32bac4085f0bdf36242cf59b555102f0b9d7cd4ef03c2d51617e0e069c7a1b54e6e2aec3239524f095f2bc2b60af58fca20ac706ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f5be150a07641cd5865be37db724efe230f31ec074e7db1eb009d429b55c99afacc6c3d0fde043e4403ea7f964e1f656b9cdb15ab9e30c8f010bf5e85fa11b5e2be9d3fa0b242817d20365b8a8e632e46a1055c3ce4c48fbfbb70f8fd406067878c171fce31187fb164237a2e38d9d617534f7293cbbdf1c8164d93cf55e7ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37249841ae638ceef4107629d4f8758e9f6a160b3cf44c69a9a749fedd7db3db2b1d566a2e7f32f26ee6bbd2265cb1170cabb538eb34f9dacedc9e973013dbed8ada696bd15722ac583718237c3d4b49577b8dd36d5dee46946485bdeed4a8b3fb09428e8651d1d0d89a70f6e5da7da06e8ed3aaeae767f5b598250baed109aa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf824ec7984554079322aa1bd5f3747953f33104a664d0d14dacaabc483917903084c221f483754c96a866831d3616e6caebb39f8e1e644ff5e662974404c440084a449881cdc7180aee7f608e99734b1f0555e56c187d233a898f40347356a18edcda41ddeb71c72c3529ab792827c27ae9a83c9d5020a4bd00d293805631f2d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haab730336b35dbdbe2a977aed2effc73e6bd20f5cdc37479049aad8339bed0e095707276804d277c9ea36770889151bde1f7f6738fb8a105edb793e71e9c2f9c77501b5872aa39594a60bff853a5f1bfcce99332c89cc1d33eee3b1030bae298f02fe3357c0d83cc1cc4452b9f1be3a4d3351c80e934ff42415cbf721923cca6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h748bcbe08ea37a8d2e162c99669438071abd233082531e86a7dc63ffa8b561caa4d5a034272b933cf5789740900396c4243d6c13915e556b74e80930e34ef4be26835bfd2b43d985804faa1ede63beb1ab39ec6604b46a92ca23a4a85fc9cfb59f4a7ccbe0cc278d07e4905b0c032084131d91bca9209ee142f84a91db3a401b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10fb15dac8e4288c6ff6301a2d60074421dd15726a56ae290f8c7955cf0144837e459deeec8c880572a18f4986a4195887b060043a6c49204533fec6157e50ed275560c78a34818639020b793f05ee2cee0a07cabb1b54254ec876d864c3faf714a352a808cfdbb031515dd112cc9c537448ce81f00b7548c46e0840a08c0346;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4917dddbcbc9fadee07330fe6392878ba90c4b6e91caad60c483b2e37577fa79bc46dd04b448d8a61d360658daadd7260aa34ed0fc1e04b5a5ec8bf7de3621475b56141c0ce1e702c2de318f6a5f8aa848ea3b061b9591449014e5df7854103d15fb8561895aa833ac116707deffa1158e351c06729a61c2d3e3550cc5cfa86;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3114847ec3c0e47ae0e1ac01eb52ca1c8adc52f5df2f44a15a1b95f09b14dc885cfc63a8c78f632291a3996a3dae7545c7b7298f4c078696018c0b93edfd25b2c66a0f7343c79e6583da4c19e1fd9b89f83de51b88580dd45c4e771048ab8b473e9551fb2c9fbfeb7d5f483db38d7f25c22b47dfcfaceedd634f0d6b227e4a50;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h768b2de00c8260308942dfc8ba2d4670804bf951f2c4547927c79c2d255e0104fc933bc3c643aef25fa35624c745da71330e74a1c0596db83ada8036d31a1e2e6422dbc5bbb50e68a81774cc202b51b2febfeec449a1bc6cf4af904f0578a280d3ada9a3b47143dee73ec1d362f2c8f3a09911c3381478f4d9eccfa054de2b77;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7dc15f00bfe92c933ae686eef2aa3d20eb97f3c294e6aa2dd8a7c059090b3acfdf81dfb2ab23b8c5bcc3b38e9d57033813428e68bb5c1b1c264f1a0db3e3e1bba3ada033ac7848721257fe326cf4936351019ed32e4941c66ccc6e439cfba755edf86505efb99c1fdc556d3d83b3543939c7aac6642edcf82126e3d4dee4d275;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcff7918eea17cd6005c7248da951e4d75384a79561f7f38d220c4cdb9a613b366d1668b6a2e419cb7366d0ee1ef0968cf7ee04851577aab9445001f0ac017c11281bf948b3a11e51011ac0fe0c72cdc48c672f9b5c5e7b213962bd9591ea5ada81179ad9bc3bf0bc882207470911a3ec865fd7f9e713a909e4b7e3cc93efd67a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58f2079d7a3f5203ec225486556769d4563ae88ddd6cdf2e92038be2dc5d7bf3e2bea6ae97f7085d4e9183e94d30c97b384cbecbd4a220c217d370f7fdae10561e2783405c80483d2f1c06010a9712a1309ddb97ea4b57d46637d7fa4b89037ec15f6aa23b67c4b25b29309bb19188ea3710c5ad0ab4a307f193d3b687a88ae6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29d9cf5d967f792729a593b2b07d0e7e67bb2a864e6d770875bf49b6a4366f572a97d027b5fe61f823175d095f7ac5fa1fcbe5a6696642f0283eac4a7016d9c8b0c2e10a73ef7586aa537bf45cd697aab10bfbd27615a867c42c71dbf22be184f9f37437ac336cda4a564d40d5776ae563315f4b36e533aeaba315fd3825cd7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c201f37190723867d7272d23d304e091ac160322bbec9f352c3675f5500b8bcc9914c8253e3acea4e4e287fd45e4b85d2d6dfc4af6e69906bc788e8f88d6d11dcd469834ce2dc565a644496af4cf3f7ebc9df862b11a1ac05d212158ec3da070f52e79c1a94bfe6e360fdb07f8ff2a35050b31d83d476b872f4ccee8d343b3a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he955e8f473ec4ffcb4aa481fae08c60786de17efd348856373741a987701a2a231601b41996eb5f61408386fc6db4b969004867db00492eadd24669b208bef72535a7abdacfcc19aec4bc4410da7368e4a23a0b9ac0e9f86e934f42465e28639bacc90a98666a62f05757ab10a8be1458f355f9758b2c16157b6456cbe6e423d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5abbac72ca3901f85178fac95354fdd2ed47bd7776a69482c0c69e20161db0740dc23d59feea7b4ee833c6048208c68a92b11f2c0a326bc54afa88136ed158eaca9321e55632c9c704c75fd9e8121abd619fa26bb8584591bcc69c2cb7468a373fd68aafcc8040b939c50944963831c86dd7e8221e432188105529eacdc866cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4b2234713e07400509655ca12239836e5fcede9b802fb25bedfdbf7e5225eeebdcc5bed078e26b4978de3669b3e2ccb868248497cb796603f4b5a702265103b1d6e39570d9534083ec449a2f131d4874c7185bc37094822b06cddd42acb4e76e0718263452c8a03f00b666941529933a6fcd1128e2177a0d2413d9933882f15;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23c18b5ec220247789c1c641def15a106cf53438b08d9813cf828b30e6546f943fb0978b24a01c3094b2d145da87c969b8277f60e53c56223ed5df9237ffab2c8c8b74cea70ce7b6ebdb7a1afb9107641d00c62548758498ed3212c72ad0a30f6242f00deea6b70d97324c2a1b2899ab43ce2593244e7236aed25ea06d362985;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a6dd180392eb8c3851c137ac4bc9e063b472cf1e8c58f7368ba01a61c931f96e33ff19f20c4306af2fe0c7f17db396258c4a43b0281e33915efd5c7ea7d907523521ae1d0ea897cf24a7f6113566e789ad39ee2bf5a98d18317d0b43a273c64dcc3b1a99e76685ef31825e22b149965a39337e320873361edd12f3d4eaa1aa7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd2418ac2270b075e58fcd2ad6884c810d252c065ccc05d30180747190841b061293ae1f34194bd8c19df4d9809cf48ebc4a4b322486f5882cd54dd300f8fac900b801bdcb1d95e64573b6b568034569f17cf70d3c85f29ceb3510735470515b533ea5c6a10929836a3a1ec0caed8ac60339801f87bafc5c41a8b384add1177a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h358dcb0588569bc00f9b36871e3b4c57e034a981a0c5ae938f58fe887df12275f43655feee8739e7ea9b65c89f7467c6b78cb28e57c5c7ad4b1ab8490ab8b641d1ce8bb9f0a4fed737efdcad9b8a9606e7b675edf3ba00972a0f9ba40f83cd0576688333cfba6d034f9f37bf04049dbbacdd44d06273323eb3b9facc8385e469;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95d6e9274d498f4515cbfa2af2a88d9b5ea40d6c34e324cd08faef2ae43aac466be5f51309ceccf9d10074de98e3d54f6ae8bf203cc23243897615fecf009c9e359b1285ddfe115cdad6e0a8102d42ac5bbaf10b101cef1f396c27597702456b41b0f8d22e1c51103611d7ebbc0ed6601675d55d092625f731708f51788176dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hecf245387599b5a827471b9b9317e4019a5a0d529d314d3ef220c05082126e571d965e847bd22c21e094a154a00d714aa09f003a425a8d4e89aed89691d9bd84c76c3d537d588d0ceb193a66aebfc96cdff1450cd8e83841554152fe2d5de1a7fde92a4417463da5c5fecdd969a06326a7436b9c69f790cb870e15b468c058ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b2fe648b2d8ce8551261ff4f0487cff5175b921fb7ecd4d3f9595e7402e67faa82525f2d59154817bc9d2e3478058d8e5ae44c55aa25fdf627dc10c55a70e8ffae57ac9385a5a6688d3e7b28530a1ffa728050569ab26a5ed4c3b27052801d2f17228f4108a30a829700aae452db0c68287d85354d2ebf1cac70b784d096e4b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b9b29b0063a4ef1f9fcac73520693bf4d1687592383b31db31d09578968fd1fe851863e245a1d536e5b4e1f2369717fa2edce0c46ef595c5228e23723c2e401d05bce37560a66d715a13a801dbbebf90820eaed131a1ff7492894b244b1d3bd13f6c72b20642c1801a1544b1d0015ece585c9cdc7d733999183263ff471f288;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbc4d627eee1baa4fe9f2d9cd80edef68d4e18d2a1da32587861b698e7886ddf420a244af6239728d4b5acd8356b7e87d6c6fd18fe93d4161505734e4302c57a76ee0e6523f423dbac0b1476309e2d920ca7c01f8fdb9564c71b33aa3a360d5071caf9446ec7858100351aba808152d91c02f409632f07ca7b390065b0f57dba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55eae0ff2009ed0007bbb702da9b3c962debddcce030924435b4d9cd7ea217fd2b772598fd14aed63f9afd6ec4bfc5ea98ae7449fb0c763c75ca5ea6afba26b23c443e6e0a13b1431cde615ffba964c8fa7adec218357d4c488ed234ebe8e4cb8c2cd39d7db0d3405633dccd5a1214b2ca431f589c5a66abb5ac91cd4c6d70a4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5cb0a1fed1ca7cd8ee58e8b201d30cae95a5dc55d33300d52059f8dac0971f8794a8cc624d948b44169c2674d896f31a0665d2f535ee089fedeaa62ca14e93f0c0f1ff7e72454eaedf7aa499571f94d7d93b935df3cb96a99f98da05e67f63668c139d7c3b6a3052de8b2b49a4b118c36d48a27a93156f34ffa18ddaafd5d85;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h659c9dd1bfea273062cec7c027b33c320f1003679cee6c38bb4ec5e84dc077912cadd0fc35b4600bd35d2e2eab877abee8d299d1bcdf8850e68c8e2856eabd543d8950285107e940fb6d0a370c1d9e6e4767f5fe8e46677b49872a409fe6fa82ea0831379a2932025bd86c600f7d522c0b26f4a9d547d9bda36ee90df8c5c4a7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74d2806f21faf7532d85e1fe5f237552235b5504da74c4208f774b69b55f2df89915d3787152600407e3bd304e8810b739dc54c14e40cc8fdefc520a4e7e68be82a27777fc99392f2fc189f7cf162c792f3f3d0fc3bad953b492d23a3953a8b6f04410f6c199546c3c624e4352ced29f639a997e5878b560fa41baa278b42beb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa9e030a919b711a5ed6a4c7a846ae76ac70513a6136f24a3d8b20dc470e74031e3d792ed555403c4f76db6c8370e066b13d894e4104c1f9879d07e287a4dc74d7162902671934a4d6de510a993b617113ee822284d880cf5e390c3f72ff40bbc40e9223aca3d9bafc1647318b6c862c1365290d9a9bafd1ed3924391a67365f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2cbaa5e4684672155b83d55c146579f5e7ca510bb8306077a8a2a9c64f766b89976336201daef52b06c5a11cf910218a84e00021ad96ec7c9231feb496ac61ef4d94b0b94fbdb670ed63c6c235e37d2a0ed53fa79658f5d0a7063ab817c83871947eb1563b661a6a4de0f5bf4f312b4e1d6d0ba8594cce0715cbd264a576911;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9966e25150ba6affe9c75d34794cb12ed8a12561cca5dcc6f141b975cd948494827815b63a55cb627122b69ff1b8374ad970b9dcf094c3a6b2037b8ca559b82a0f66cace59b14d331e1567279df7cd49c2bdc1b11836b27f47759db80de3f4e047579bc60fa45abd056d06e130c5f6d1145ab03abbd4290be9d0158ce0895be8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8c52dd7d2794f47ed67674ff2024c03d15828c6baa52888505cfe61c7182af3f267125b5bbdfcdb81fe0fe1f1566101e3db79ab07e9272ec89a4d2c5fa20b52bd7d30bad60c727b39efc93587e40331611905de9e568163d3f42003bbe092a71f6836056be4cf8ee274fe68339bb2a063a701fdaab889099586f9b1972d618a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12b43dee8ab2bce31eea5e01e9b0a0ff91f6eefb8cc36bac85194e7b8e02fc6e7ffe1ee639fb221d28cffd8f3bdcf9bb0962826b5f2959c613f8e27874bd7189c482c7b6e34c2706f3e27a2be1c8e6defabc662d32bc62449eeaa7abe05a3906de53a16762cc0d0566d6938df4ecaf78fe7d915d6cd3f880a16be53d4b13a351;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec6c1bc06748ce225c703a47e04288d57815232c38ad507014fba05937baf8cfbca1f2578add05ea185d619ad57c15c8fb9a0da00be7b14d5377192371694d7a5bcf7b9f44bb2e2fab4c2d6c958ec18fc575e9b9b865073a3217c395998c86b3507eb217976bf18d6c7bbd152b8fe57e429fad69d118f777b9dd843056260794;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h77aa67a0a21670b9d8ec8dc560794f4145d2f89aac0561d5e2f284b72554df818ec4c6b5f11b35051cf141875ea05b085ab17f06f0ddb70c5469e3e03f6933cb9de5f86a5837d0134c1c1914f5163a49a3447ff9529b957b1a478e51e0e15b541587399494d573caa9dc1dc2c5086ce02fc1dff6ae4d569ce1df0ec6de56cdf0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e9f2089275d01e1c6a162781cdbdd01ea861ec3c0a6277f3da0a854175885eef015131637398b740a98ffdb39afe73f70cafcc93c8e4ef78c61f928871d03edd7d19bfefb6024e4ee45307441ca046d980b14a1401ec6365d0d286c9fe2c9150d526a32509dd5c46b1230d3d3f6c1253983dffd62369ce79a93275bbee8bc77;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bda1586cf9ebbe377e5f3b033af5e155ff0cbd9a99ffd1b6cd7f4c2bea4ab510f56a17d064429eb925f961ac5d0f7159664cce5047cbc8107e18a2475984c864fb99bba7df56b86cdffef245819fc1f4e77b13490cc240a96b4f78286681ae029719115721365e3fc0a01093b4e3ba4050e0ba973458ecabf42560995c6f5ba;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h577ec8a8074fbd5d1f62224312e49eb88136ed4a7762bb85498e6b7fd5779db5f80dfb40139b354ce86b2dc3f492ec484a6f7042eff358cdc938e11779e0cb032d849042d85257673af112c06a7f6679c22e3b9ac8a02c5976e15a33f35ac3c0b867c43e196cc13f1d51a5af9f9cdb479a4d2ee6118ffe7f4916caad77f75066;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40276a801ee9f7ae09f2197894568549610f0383fd00349b8f277ce2e997c71ec2fb121dcff921b817bcc29aabf16dbfc24ebef4d6a34981a2c55c5642f71dc0e6825f9c935693f06e68e7f8b36c474cf7b66fc2f4f849da1a2eb5faf8c0d60ccac0aed9db695883e6b830ebc6afa3efdacd8eaaf55f05d1582b2140fd05785c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb239eb1d8d66da214e1d1dc2ce829c4872f2f66ff4d863f468ee5be0ce08ee9b7d261e0c8298d85c4d120bccf5fb0c56a6ddb696861310b7c7051778a673ab4aedcd0fcf08d50259e0177a6d4f27d2c5ea79b7ba29eb39f5f6e982d14abec1dacf6918da67a747ebaf255f22971deef83e1b0fdb8abc211f44af3f7d8fdf826;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6919a7814ec0feaa3f7f6f2f2d5c4f52984f53cbc5fce8d34cdf5682f22e97efb83e583607b715193f1eb7b11c3e492f74b6069fe47947859074c3aed9ba998acaa1e3fbb4fc96d6a696ae67a321e7ba344506944dd81bea6d4453ec60804f95ab1cec30ee0bb72ba822670e8f26a77df1cc6c78e02f51879aa9f0e714ff261;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd37a7e54cf407ba3c4df18fb02235e5a3e4284e8caff7650bdcbce430e88a53bad341c644e474f726f51a31cec2781d0be4d424bb468db4d08f343fc79ea3562765038bac5e6a07d181fdee6fffe9eb5bef194ca7733c049cdc84651028644de4b31ece4db08cf8c92087fcacfed571f83bbe00810a67512a98ac7ad1d51eef8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98918e0d4177285ec376fcbc6ddfc37d7c75fa61d266689fa4284fb7f7964fa469c3a8d9f36b059caf89bf446af9430084ad628c2adfb2b9f92e581520e1b410e5347a7cbf6cf92e38551c9d0bcbcff9719ffd5d5312ea498b46217135af48eb4750850281dac3affa9cdbd0e3a77cdca45617d9d89882b034cfbd58c7642d73;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91a0794f9f700a7797b9b42915671c2246e2a3def74b81f6f361e022195a86ebd0ff677916dad133acd76188012ff8b8fdf8ee9c9d188fc44acad0ae805d949e3d7fbed201ef8a38f78bbbdfc3d774ec665362ba7f00684b7e47e6b925f4eab135d400dea3f360d776ee49b12b78735e69cab229718086d8555ccdcc0e032135;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91f14bdc8132e756f60bf3dbd3d9188cf07400827fcfae612721795cc0e4d496471b7481cb0db2c184a6ea8e73d793b29f5e12a3adffff2f9c7b88448dae13ec8d0dbfc14c9d213ea6cccc89b9bb311e891d478da264163373f097c7737f3455ce98a239d953157c3546d73e5f7ec21391daf113b4a39a48a48fa7f96f2e6d89;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h349f4ac1ef678ce5bcbf970846e84c33b31f4ef9449ea0bff29df867d8c2fba8cefedc721ff805d3d7d54dd6d589de76fb977f050134039f1ae291e0bc0e025ed18bce31a7a21145bc20a84eef271e7496b6b11994dbf3dd255cc76dbcf3cdf8a3725877982e4a978e93d6536cc530872622f06dc0cc6bdb00c2d58c7ed8556f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc576b9978bd174710848d69661ba9f0623a3946a7f01173a528eb4e695c1371885cd37160a869c2d91b798897ebc5c91a629d635f3d6cd06ee30e42daed17de9b5274387160658bd18f01c02095263118d29f7899bbf293de308d80825c32b2caa6da82ef15a8a372547e2ea2e2e5cdbd9cd9e389aff9f1ceff288cd75af08fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf67ead076179aa7d2e40b459fbdccfd6c67800c2b9b0dc3897b30dd74b8bc5cf69a88839b4ffc9916a675940aecbb3bad063f2f9a70d70549d9522e46d7d8f036e4ac3e866d54c1ebe5304017c1a7040fcf972f890ae47870fc093c1e94110663da0210d44671e28ed8ecd277a6c42ed99b32573ce3a8e8c7957d1b6eb4347d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h906e58ce4ed35263dd278441b87b8efb574174b2f00545f99d204c28a565b552bb390a35d9ec53a9d3433bc9ef9fe82f23b346a24d59c0e7b0b17dee5c00f7a6e37504824e9fbd6770a5cdcb508bbdf9f34cf04063198b5d9c0e967ad754b0914c41dc769434366b83b508c5783d505248de31e2e4f2ca5e48e6ae22a6c3d380;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0b22ac26e113c46ec7900afae34949000be5869dfa0acddf303d8ebad4537d000248537f8185802e6cf052ecb897786c5d0818cf15714689a92a36d67b646b672bef4b5ef8784f956e11af96aaa1d7bcbd9d266f9c3bf8760f2237bfeda8b9fe53e6db73d227a516ba4a87282dac85c6d58bbbe163a4b816ac659e798f9fa1c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d6050e009dd6426ccc6b348d8444da7e360df8cbd2a101c1d4b11bf3728b23d8f37c90aac2d26205f8c28af4532669a095baee8cbef0d1c028cf151444ee9cddfae9b034bda6e90b612903576985bb206269c5ac69e87e677cec5fa29e0a4092873d004549be5eb0d180255d0dc5182b39acb298213164d58e769b10324d454;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b65d79bf2dd5ed53360200dfdbbd4ede75e8dc89869c8b3e5aebd8aecf78b4b5cb936cdc9fcc61e6be08962feedb81f98965e2423d4b16cc4efce93098b28471bef4dfa9aca84ef2cd13da62992318a111b51f83ffca2403514d8740e3b2938e870c18b0514c0f6d875c30f7d741193ade00ec63563f59795ef1afd5a97eb92;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c4491edb9f395703cb999b7c0e4004ec5f4da6061a4c1e7341161c64738068fd08319773acf663a2dddb8124573947509174fa9415f99f897b22fc0f7344bdecc236d42c5142e96463c8ef3eed0699087bdc89442ad5bb546623dcd3311d0de42a17cd12e04499d29c368aec700250dbda5b176e3fa2fb39496bd60ee96aa8f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h531d47fd5f063043031c5720db893664a8f52abe4326bef15ee1bc3521e2e1de32b6de41d2acc8c2e43b896304ae43318034b7b1626d257a0c05890868d3bfd228665c83610a212ebb537f5271823d3f234cf300a2ef0dd1c09a89add8db3f1e87487672c4308c4d7b4f49f59a7e3812301ed287f38a2af85281d924492a6519;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ce4306a57363e16435550ed3fb48843e84187342518af1f27436d548896bbe2d2dcda7821f2556485233b2dffb6af89294324a65eaa6d770b5841f9ff82b8995cd9b0c2c5b9337244accac2072c5249e1cc518bd40a7756774bdbebece93600f77a83aa0b9ae676a951df312518e76fe57e9896f5f567bfc86b9ab8ae6668c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7093bbf256d3d6d6a5592872d3f5f1b9860756c400b5263e484d8e8d2f875acd353221728008664ee52ec711bdfeb96fa2d20393bbf39f7e412b33c24b017f9f655fa2b417c0347a3274f97b8000103f0dc867b13f7468453409b0901efabbd2b76d7660d864c6341920585f97e7a7f554a2e0156073091e9c3c966e77b64148;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha279dbab75996db54533687014b576d98000c7bdbcf4a4686a06950e2d71c462347043c2fc77a8e4de0264715da64865477c707b84ac1006ce42b397e010aec46c14e3aee05a6b48c8e0246dff518cbb9ebfe7053038388a8531020a1e9065e1738baa853fbc8b294f1e44274b38cc1fb63eea5a176fbbead5c499603e1c58f9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f1cebe89c67cdd885fdc259457e90c0203adda68271f9ca42e547cc3df02d5bb0ba7ce461131b53b6115b5c22805ebac4540803d86c80f62d55eca0c7e8457458359f13cdc2e4e13aed7815b71f408faf33ea1aadebcd78f807f05c1ef115132d64c54eeaa464bd64e7ab78372b3227218deea77f388293c9ab9a188b08bd52;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3fbf408f01b735fb9fba9ca9f2d539637af1e7bc1b81d5d97d8a6635b5ec313d6326b87b74003015f056d1fd2727afbc4e6b39a6d6c39b311698f4a4e9071e504b94fc82321349f85e7b4945be2bea0e513a0e61a1c24f27a8a54791c9d5926a3caa33954c9a5472e3144421f4017e9d1868f99ee5d5a26bd4b19058840bfd9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bdf240f67c01e4a53600e0e9767035139983c07c967326c48d7dd20a1f17454a0f832423eaf77b80bcf11ca127491af0a89e3ff82cd0474724098381548533b4ebd174d1bd7f8cdccb27697c7b844865bd643dbb237aed94c6d49627f4773f14efe178a4dbad4a79c59cf25f17f2eb6692cd80c8a447f17655768ffcc10f2f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef9731fd97765918a5ead6c349b7ca6c106a13e205db50b66f68652d6f9724c6219f87a1019e6b69a3deb6a54f9fe85f175554b0403647e27b7f78698dc291d6a17f8e0c13c3120882852be56b8f5a7fa72a138dac5e206fd8d9dfe42d2618f1c7ea7d79c8f5e89480fec94878d7d83475296d4aa1fb5e8d0c9cda50a5e9b6e4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3754ea6ecd5be646dcaba8af7c4dbd0454248154733010e79ba45cff3b2d1d77ed5aa3242cda7f774159c5e9f678e2526a4c9c7c5fa1c2614aa66c1587c1d42e95b55889384027b12920c8d2ad4601c3fdf6d75f7c82281016f4ac21df63e0c08d40f1ecc4811ebbd200c457827afa00beeca1d71c6aafc530c73091c2660de6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c409204e56fa7f16de8d4c470c9528932b8e9bfa3548ca48a53e03f25198f0577805f155e8c16b9d8ff6f7c8ebbeb47b24ad6827cebee013ced2d97381e02e2f7ced3fd9080db81e98390c1fa1b9e69e69c468adb1729d0e4bb2cb3af196af1b834f4b0775d299363e35f1ed90160f5c325367abbb50f463eb2e54cf8a1729;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9347473cad80a8ad8797cb65fa8fb26fc5a1b8f4170d1478e0b5df2f253e6c71f839e9f15b71ffc2e87580c1bc3fc33ac42fa0a953b3632c5fbce59096dcc76eabbbdfd018042a6856015ba97042d733dc9cb68807b46caba2add6d7beeef75837549fd1a5a308e4e3ab6d38233f3428d40abab4fee9398a48a66933ea2ae3c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h413d167c62ca40e7b233942101df020ef0cbb9385828c817d9bf2d204c69459ad9b4315d721fa04836159a2caee8d6e348bdb1337083d82c30c1ee2d4bd186c8c115db0c9495bdad3ed121a44fea2f6539b6783f641355bcc3550d7d8c578b987d2097f62c6a5263c1330cdc2e993291784237a1e669edbdb4c58199bcccc987;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb94609529c5e7a1e1322efa3b543bade34c281c1286eb149fadd1b080dbca114fb485da229c7b9c7953c7d08264a431d0f82d17446cca23378b09da4ff36588940a1dba2492c6a53e0ed971451b30f03bd67efaf89c6a0bfe7a72c445803ad5b29f5ae0662a230047ff55caa738b61bd994457c41b060b6fa74618406fa2816;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33d88f7118d8a4253a4d28b9d59cc66969a873615a25a89c416e3adb910bfb3d406b745e633cdf8b2687ee1d4705fe0f85beb52bed3f643077f6a5d411806ea80e4e5e188488721cb27b6992b40de7ef66571c2d599cea186395ce59de8225869367f84548e7d22a357cd0dc39803c87479c3148592d8933fd6d3bdb37044d1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53be3626324eca665eacecb2801fe10da3043bc644929d300dbb2118eb1edb428aea2f3a857585eafb0e4038eb675586183ded7959b716cbad8ec0d4822c571583a7c2a0deba68a65036f7a1e01310001c6a29beb49a24e2e05f29fecc6f6ff3dc0789bd06022e732e5752a55e61b651b0616759d3e8ba385cd17e5181f4c9cc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h854a113525f69841c7a6be005350d029114b9ba9e73bf177fdf538d08d62e96aa74c2d8fcd0dc9defeb6a135107694773a8ad31cf7582014621e5d673684848f307c1ee0bfcaea52c80b0f2bcc913ae19a8ad248c8ed1b6cd25415370682a0fef257eb4eeceb79bd78cf6110fd965995888ed7e5a30ccfc76afe1ba749f35127;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h227cea9962ddc30531d1e7607a7c5c6dda5c54fbef0bce2232e591103a02117b0a2a0a3d2e607aac2f0c34a96a2cbaeb3f4ddd2eb0d6d2215906366cadd08a27bfab7550b61b5ef5298b73beb3b5b52eee1539afbb42d77322641c4d0d82334e426c2051815c8c0818cb9fdea97255bbbc9b0eb1763f73ca8a0aaaf1eafd9417;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6e6238d59977f9b9f1d50cb2cd02a0556980315065ed97fc54e31a603c4d3fc2330c3adf65231b37b47c1f3ff1f7cf6dcdee3077714f558a8d607b04964491aa984815b5b223d2765e019cc1d72f3a5449ebff905bd159af9de01047297387d8571767fc2a921d84527fef694ec15847559e9514fa81cc1eaaf2df9c27b9be1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h813194d2183e5a4acf78060edaa49d699a3ea29ff6a4d8d412939817a37285280206a551ac9182c7b8874e3bffa045dfd089d114960b44bfade68258a434291da8c2ab52e99fcaf4e57dafc814ecd08b4c229535ded1cbd8501c512701ecea67da0560c53c249241d85e121ee57d46d269e280c2f3ace6938a95e772b115cd02;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87628c4ee5ed9a15ab96da1709ea575db229dbf3fd81ace23f5aea3249ab99d4f4a4e75cfdb81e3d8249893645471af184102dd242b25ff9bc7abe3eab73192f20e27188aa15e1868ba915814b94fa0ccdef2a118ceb86859060f00c5ad4e5b80703e2efddbbead65041b54a972cdb8bd151ebb2951045d7801c9f61960835ff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3438f9857e3ed9e096281514ae6b42923f29975c26a81e3b0ad4e9fee00fc78d6b462ff1d1388be077e97c34881eb6bcc3f477d2bc3b44d4040ebdfde1e147bdb33e6abc19261b5bca4bc6f1a5829a64ee0be4dcef43a4e729e5e0addeafb5e7e71a144589e55186946b12534222f5a0aca3723dc17019b661ec3bdf9769ab66;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d29d171b7e88a27eee4135cede171cffd16968ed0c28725f9da7017ff3e2d97377829cf6f505c500a8f0a0d05b7b9a221a4fd9bc9357c9468ff6fd8bb2889cafa82b57d76b5cdab6e2cb2a22d1efc4852b4832357cfdb390b4a426d940db36486c9e02befd9bef0254a8a0745cf64378a2e166b88e1ab303b79ac3bebf81564;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb6911efa2325db7ee58dd444c89effc1593b75dc81f6f7feef6c5ff1dcae57e6d55e8e6f03c7d7b42778fd7bd8fd3acf442c14cd838b7c4a76e79a9a436ef84ee509f8307130e3af572cfbe9f9752cf0e5e5e8b4d531d77a4e71d88898a80f0f6ce4ced15eb18f078edf79dd69745f2972dd495c366b865f458bfe783924d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1287b0b81924f92b0a54a6f6030721283ed7702cc62f16ba859c3f8b3909ec9acd9f5c25033973f104eed63af3617c19d47403a62bdfede93cda63ad32e760242c05cf51a9ae5b6086561d7715d934a54b2decd91d6b448e687e0bfada0349786309cd078f302f33fe3ae0c2a5e476ac62249c2cbdf76e0191ae91dc20d42c1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf40780e4dbc7ee48b21c0bbcc12fc5d1e816bccfdd7137710c9b5abde7fc2285eff0366569c7793a53f648a43744025a7085c7c9cf7f257a53f15a306b3cf40138692ad7b89db40d6609ad9f3b63ad32c287669a0cfe75337b15cd30b715b240f961c24e1809b4d832923a395806d227720053d1c26c1eb71d0c4d018a3316e6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebf15d95aedb72e53a40f007531b219b08aacb76844b8fa0a54f0d735b00a64b104d38693eb0a21e3896b90ddaa0f7d36a3d72b030574879569236d88e4424b030f6f2dc71d3007d042351488831e0b15c7410f0e9828b641fc70a26c45abfcbb89c3832394d024136020b4a6f2461ce36808b2668f9650e97fd3f6cd9f9ce82;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d587592bbaf584a6ee6ef835fe61788a9f94d8f8c57d0d8593b8e210fbb54a02ebe5f1bbb50ca7881a2e89da24ebcbf1f15ff06ace2cc6fc4d4abe7b589dd9d9c80f3a51de933a9b07ab5e6dbb4b584a5b9236ee7e3f9ce5c4e77d47011a263e3fe26e437b4f736d34d4b069b0da133638ff19f409f2387f92bdda0e0852b56;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h827e672a521ba8d48c43eb4c3344a2a87bc5e0a6d1e275e947ae2adf031cf0044323f7c1eac920ea0f000e9a1e6233e66d51c557731fa1b19a98512522a65a56feccc10227b4512e212153c7db8fc1c17293685f68f7eaba67ef6d6a43a34813c19fd1cdd614aff66df73a35077d648b45336b2724765e89230e47e21f087db9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5abf45721c324389a387e6d3aa3343ad50dd7e5e8a41115ce9fa4136c9317df2c882bc67f0866be6dffd33b02c700bef6b7b872b465df5cb50c27d67f00278e23f16374adf2f26414db16a1ddc0c95f7f350146d2fc4676906119dc2a5bcd72e67c17359b7263d322966056d9d8542d6826d2ad2c27dd4fc1b675751ac2e2516;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h728ec7e67deab2c2ce8d9f75ba43344887d2555f3918afc35c96a63ca4a72ca8b33f524685a67d40a52fe38c6598157c9dcfde2e652a1e7127b4ad00e996a5fff330c8a018256e7c2b491af16803ce4ccc2dbe74f7bf73e49575a29de34c2eb2ec33279e6c86e6d0daed856477e5592230e9bcd86637f3cf6bc412d675cbef21;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2792a247180b64d06c904dbc432948294ca35ec73a4748a03fc09f8fce5323298411ae50f5a3496d855712a5d5b97b56584dd9c8e52dcd81fa013d25be37fe2d380cd9277e40536b404cdaf69b5225fd64e02aa1cac8d2328f476853734bd8b74147acab06d95784c6d156f3499becb54e8fbf9472eadb4544bd25a164a19da9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfcc2b5ac24e49201d7b9198e614fa4ff7384f5890d8a8400c593a5534caf68596d182fd52135e45ec87adb79752fa78659ed14347112667c9be987e9983e5561f31ff6c898a908317ed7f164d258fa25d619a3a5114cf85dbf35cd5343eaf54fcb5609c09c6252f8f14fa6e1c21f8cfb1cffba1a8ce8fb724edd252dc69d0720;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdbdf6a98d53988bc508dfdf2855273af9a143ac462cee1acc4102db86249ec67a53aa774ed27870c43ac58a8d27ffd965802c56de99fe89ccd373adfb285fe1098ae94bf521132be1704fcecf24a22cfe44c27268b23895b13b75fe4a3dcb31c12d461d35922a16c202c7defd5e75b38d50ea8103fa4c444ece8af0b01acbd0f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3163d8e8e5a2ba13e85396d0e89f68e46b30f560709738e0bd9e6698c86f1deb322518b87bbc46e6c148ed09cc4c188354d73a3dc0b482e5e85319388d5c2f734f81bb6455ab99bca319e91e36ecb06bb61ba87e70a08131f31f967bd9a2c6718cbe9e64097588d9b7e0c4d074949021fb11945f69a69dae0f459ff436e98790;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he932faef50d9ed04e1968823b69c96c0e09a0365cfcc0ddcae34f8c6b96f70db56294b40a3da741d5f2fc484145c589a6daea4b21ea4b9e816aa3201d824c32a6f372f5ae93a133e5b737b7fb290345b022760f20d9abf2def09821a7dd06bfd5b3b82a1ca9aca1a45c747ce8d683c0d94a19b0d584a3761afba7188e75cf5ed;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b842d5a7970010c7b413687534ad49174d9c5ab6c6813004916d56adb9e12e822b9943d02a6a2919b8d0b87e46f272ef6bc874ffeb41c71513a3a2c9add6fa7caa138799a41ec239da74465193660c2792061e740571b48b8ea74cb155b54883c6ecf41a7b6d86508ed3e12f473e4c5142e247250062c98c3bb6b79b7f0308;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b8e4a85908bb37eb1f238b9199fbb896bfb9878580511ea59089c7834e115a391d037c509e6711c159ba84e0851cb7726f7719e84fa4ac4e9834721e94185ca40278ef1785c31af7bb3911ede9f6b0acac9a96f2fcbedce21fb4416e70fe30326b63949208b3d4b86e0835c5efc0edb7089624fc8524fd348f46d72edcf065e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hacecb40cdafdc80f860b2073542aef02017c86149fd7449221960eb5185b1fd1bd74665d893eafdce3ba4c5542df6e7a27fb5f43af97b2899fa23596f68c51360197ba995e3df21ca31748c63f814523aa03d46bf418a10ca5b7c2b24c850784fb03e9ac04d97360e5882764cab4997ff971789cecb2890cb30cdbe58b6ec44c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb38e5e3dae19d8a9a54be68f97ff16f07795ea5e0ba5f32628f28f3c4fe8b538c49027a6f4aefdc79d4f0d0b93f3cd124b11625144e7fb42686435a862b2b32d9c9dd6203bda8f67795ac26df801fc11a2ef8130ceb60c27d0f5285393d9feca1b79e4db875a3838aa5a9d30047846a1de4f56e578d3457521d7447b5ef145a0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha75d454bc35b15bb49b5652dc2681f498c8b190f96f05cc054f7b74b9fbb89f3115a59ebcb809c97ddc5daa2fc010582367af8b54f0b1d07593ba5a96ca1aed3599123a45ed8f7d321727f58c1b675b06c8fcfebc3ec46a416ed495d08a3110b6878a348492083efd58857cf2fa6cc12c0d054a241179f0735fc9cfd9e4e06c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ca333c9cf033c5155f2f476b0285f31c940ae1e7376886f47dcf07129eb0e2e33432fca20381d0b3234c1bcb7c49f31d6715d46750d37a5d781b2bbbaf26e2d75cb3e672c62d71d1c7b7c7cb52d6332b976c7a910f971f2711ef1ef536bf8d68119902c67435277b1dbf0a83da3e8a8a93167dd9881c572df776b2941475a3b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57c12690dcb4581a06aabe6836248bb04b2c1905d320e123b650f1183adaf644f4a2b4eed248f8483fa7a1b49aaa2cf591186ad6ac320aa147e1e7cd42598b58f4f6bdc986b61101854013d7e1af8b02191d71ae8211e9cb8924f223f4f613a0aa1c680d1bf09b565d211593b2d806625dc22563a06976d2381957f844ae9845;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h263fae989e5118329cc47ca4fd163356dacaa754aa572498c1bb8a1df58b6c46f92f5bf8195389d71d77d44945f521599bab1b79aec4ec7d8d7536562647a23e64dec10a6d8dd5d026013a92803400abdbafd139a86845d2f586a52bcf5f16372e95d4c9552c1f009a5ecab9f2943a7ae6b2244519d20f23b735c583e39cc950;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9ed748bb95ed3b8cff3497797fcc75389bc6f8279b9bf66f00ba9fc420abbe629ee7b5e7835cb3551c632d6ef9de24e2d7cfe3d7c21d079c587a9a8d4204c147e8563aae0c863caca3ee9644026d5a25b5b3d9704026126e60eb1e8165f576ed0c44b4d4ea75736e9e91c04b052d49456e03eef986e1beddf37b391a3e97b97;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d34f3a701c42fe4d78f6bdd5294d6aa9d232f9d3c5b8cbcde6eea02175324896f49bdc8237627907d3d3d3fafaa693423f2559fbf421463797f729210e60fe3c5ad764ae95398b9ed31bcf264d1b67f29a5aca57ddd62387a83076a1da3f1bd0f36ec1bebf51879f566ba5cb994ab8e05f6bc39af1c4a504ebc67489a8df5c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff1efeaa3eb98e95cd0497415d163a1cf5841d5341df93a7caae97a92eb82db9856c92fc56d090921e4ae5884851e5120434e3f1199ef25612e75da7137412fedbd22ada7802556f16bf80ac54b8ae1c242e1159011f1be3f0bced16b3bc7fb11a0c2c5d794b44076dc95039bdf8f98098e70fc0ef3fb164f715449e847d3206;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7d8968f4c42bb8ae945d50015babcf4eb7748501c862e1a26f8f5f7e8174450e7cd3f347a61b560526a35d09286e8de9d4802aeabd76d46de3f68b8f3702624abe0f76288c3f976a667c1a04acec75f446c3af8b9ce20b34f1de5bc3ecdf47b8c78901970efd8a2bc156beacd00283ccc06bc37e8bd481ecfa7fa2a6f790d27;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f61fbf12ca1f81645f1e39ce7f1f52d5679420ef892e3f8351aa56ae6b422a72e599611150fea142ada62b8532b1c5d0101cf6d040be63fd586b6cb3b68137dd608dd50250872eb758af4ae8035da2049670d42d051fccca7d4557f9a53ab1e14246f4630496846f94ae524371f5a9af0d1555b121f10841a96feeae4fc44;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a293e2fe8267a409976ed770f82c6b09b25d691426c957e458704211bbc4d68c73570f4d472c7d9698a72eb47a43a3e56f0d65bf3a48e1a8eef9b43b68589442fcb40f79866e5c9bdd6f29dc1865ff59aacd3b9729a3451229e6333efd06f086e28414d93e63b27856120ca959d80397dbd66535e258afd879430b70631b73b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81ffc9ece228f0f7a46e7d7716719da980ace945bbf342241c6aa2b40b2dc131192f39a954ce0b2f8233c45dcac2bb8a433db01664c2b2375f0468ab922e8df4bb30917075db2719e2b997c7694e59c2150c748e74ef287547a8efed822a7f8d87c91663cf96d3b426f5182e66c80894ade6b1ca7d63a9cfbc4b59e35c08ace3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e4c378f82cb39fa7e054d7a7290c1f7d7a81b357412800d99b1660b5d8b27dc0c5ed563a8be3dcf1b69b36a8cc269a0e6866a4cd58c9ad7a6824d102d497d9ab9c478848080836a6497225848338cb0a99f4fe54c5d0b1edcf2a6b75034e00513177d436057457f4d66fae8bd3da3b53081e16fc9a7ce9d58faced679addd30;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e4086efbc67554ee163a8810c6a4f44dcbbde62723166e70ed21037a4b9a5aaad06f288ed7c57329bf0924edd89307566c10ac52b5c9f2e1a80659812ac1bbcee90bf637925d32531c83c1833245a61efebf2c95766e15fafcd2fdac5cb31bfb5c360a527aafb7ad555487a269ae68f308ce22bee95a6c0b295c0c5c1529d47;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc16a8790745015008c8887c8286a9516303c90d58a288f8d13aaa7c3dc90a11c87d5d4724a705519126778071a04d988d28b354cec024e3315c8533d4abf02751b209f3a88bfb645038f02f3471963b6b4cbca21de614809dc42f72e90bdb4736d1fd5726581480b3d23a5dfa0853f8ab226dd600d99e484e2f849b503c3847b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2029c1534cf82e703744b7c1c12b218085ed625251555534a830ac80d3182cd405c7e2511476586ec3c64357dfded2033b38245dc492f851ceb73ced3b2da288ca3bb16264a9aa56150616c2e64777e68759cc4165d65464537db84df1bd6551a2163509fa14577daa49157912daf3bd41baaba6fd7fb27f538c7bb6b057e751;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25c091101f892d212ca6a2ae5d2bccf41bfccf5baed115c21a5cade3028c17e75ac9bc36fd3f5b891646072dfde19d45b917d35be528abd444f2a19dfcb93163de01436a5a507f236b67e5a9954b294b6306a6534c6a33cba769bc997f253cdd280c69c9c403de0fad11bb015a5ffe59d3373943684e44a76fc6615b907dc043;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c09a117ce07985883619a4f27a5ea3654cc4f203f42490bb4f5b8f64777aad5cd6fbfd347df3351ff381782e86aa1b0603d4aa8e084397b5562a4aa9ea505bd445adbb2ff751a19b5fa23a169cbb494f527be7ae895346a769d60d9306b3323ce97a1989724d6b018a3f4e109af3186f4529f42baeac3059c31230331aae709;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7fcd755b69e24f1ed65e7f5a8e9026207a3573b6fe84e9969c982521b7c2bd90e17c9dfc09c67eac706d76e201e7193f1ee85bae5160f7d72eb65d9c55af37b3fb5fe3c334ef872153fcb53b7333b71d41158ec9c1d27b9f6dc73ab02139d27a4f45fbb813e78bacfb4c92bc860ece52b3a7c1f9e7e733288e2c8cd8d5f42a49;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2183e9213bfd97e77dc7cbc39e207902710195015e7165e2f55d3987be86f37528885c92c1e8cbb02ef9c5ddc62391f7efaaa9ff80791ac0ee56639928cf9392bdff8f4d1cb115be0a4e54aaadf0bc661c40cb9a3a02585123f21a161668a45744294b722d94c97fb1f9f061cc12274384870fb2b76d479cb49efd7c2ef436e3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f2359925fe4f9914a7299fc345b5b2ca252fd3ed73b71989237179dd342665e0a57676a70e2cdb8fe06dc3755818176273ca4939801e651f88d0dfe2fd5c4dc069e1edf39c40fbdff4dca8be17f3bca11b343996bdc4af5c98625d3dfe10844e9131b9939f54c5f680cd93c0dbd118fcb32b9fd2e12fef71d4f21c4dcd10a1a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha488153086f932f5a85ea4b0f184ecb262b87bb3d445c6f8a79192e0c7b336bfb9ebf8f00fa2307102e07c95e5b3efa91fbc6603ee9f4dd2fd39ae7609c252539fc590ae9602f91d303ec53f09769005eeba5507482d14f0f756cae51b7322dab5132b17e229f01ddd14ad56e29b0bb733189d0b8644d23f6afa0e2784aacde6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h569b34f8ff042692b6f273cdaa413b09b6039f139b10d4516eebf8007f228b6901f6f31ecdf287f7687dbb2dcc37dcc914e209a9e2070d437e5b2d5c53d0d2d8065d52d5e3e8f59e4136bc3e36dfb459b842091f3e310a35125411c6db0dc1925ebd1f4feda17b6b60707394641ce766442a8eca8b17be0a050b6aa2dbe51052;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82cfc9ec5365a37a36b2a924631fa3ac050a6474dc89263401d673f98ea93d2bd8c133920d2e9b50d5d42cf2393740f409419f24398fc1d6acbdcf7be0c80bc65f94155107af451ea833c4bf93d81a2a7696857db651f0af95e2c1675a973ea24062a177214e5b4600646d0cebc9e06f6a94060733585bcdf716e4e14aa98885;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc930bb4667f7eb3c35bfce117a4300d74a84c2b710b63f0ae45e5b100f3ca0c87b9937dd021ca45c4c0cc12136f23f7ce6b2f180c8f06e0d2a6aef7b6d7c6d00f48c0cd995e923cca82fd19e385a478c31d6790d438f3ec7a9a30ffcd917cc94eb9825c517319c66afa2d67be2c381fc122e83277359bf18d45c887b66323a20;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a5c8b0411b382c7abbd75ee272bd766f1a271170ec669b95e5570bca868cf8c14f90543a0c357781509d56c5c48b51da36014bdffc3898b31df69904d4562f2341fd6d414fb4d42efdc2a98bace266765cc577de749f2c472a5cbe702eadfa5ea91c740329afac8772e55195a6092ab1773fcc7f5d7d0ea6fec8955314894d6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3c8218ad842b74bc5865c9fe8e763eab93fe485bf8e0f2098b421c765e8aa4b75b21160e098ee170ada267c27afe50907a343d9e22996b07fc6f1d9bf86722e6129824a0fe00ecdf57469fc34a18e0d49bf679fa2e03069fed27bdd18dc8a5731810e3c0bddf706026f43a66190df43df7493af0e5e24177bda7db7b79e34de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91fa062730f9c2d768deec6e6779aaceafa8f2fe111649f3fa05b87b9fc6924720b4663ee5da29076046b4c7273300e9de4cf7fd63e414a1eb7d4b82e04727c9a38d84e1fc095eedf2362a3e538746c7cb6cf882796330de932c9a1779769c099dba78714328a39466da3a930131d18801d43982ee88ab14efb9b942126a3a4d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heaa504061631d4e0236b47498597187fd3c6e852cd2749045890138377310c4e5f3e7339c6447b4057c4c19e58f8ee53556eee71e83d46f8e885e2bb6a8110d6a94d5b7cb02c0d9c9adaee519f99d529cb080ae8355273626d84e7a865598a885123f2bc92323580f5aa290b0bb52cd36b0d6195138ff8c44fa6f0fcb4847ac7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4ab940cfab02294e7ec5bb9ea238c16218cef14397be7c1f52e7ffa824d8ceb11434b7a7986c3c27acaa4135228f9dbdbb80ce52e3a7c063d58166a32e5613def46d1535770a286bbbc87a6c7121afa64414436e420009248d978bc514b0d45c1a080dca9681c84db0d539d7db2e7e4edb5032793afae5d4fd28230f911de4e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb34e3e7732b13268ea05b2879ed45fa6e45309357cb19b7604bfc5110a86aaaa9cd691bbb52532b739980d38997890cc40833e078d0b697a4adb033a25b5936930a721a2768aa85de9733fb94603d6dce50788fe68b51c98fbaa1279a3b8ab13160196e7f8b3f16b9166ed27015bb780aaef078d97d89e967a397ba6a9b009c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91e3a499e7f76014d2b44d1cceda0fcee3de4bf3bb269cb0354bb710d844f6c7fdbb2a247118fe4a219c02823bab07b445ae280e06bec7cea0fbbd4992e1db5d8b261f9a1e67a803bc391d962e44012bfe10f52311f6ad2c543a9090ad891aea02c61e2918aa4e9aed2f410ca30fa1c37c83c094307e8633fdc662bb62a1b825;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf3e16c1f539f3a5ba3215c7741af9fab667c000cedd043bf83286c656efda021d665fcaf1bb05253c71c02de85cad812d81aeb69ba76b1417a26b21df7bc4d94f244f18bfb17087b4cdd8f2246e16121c1205694908cdeae208d3e0710fc6008a140281831191fff9ac62669699e138737021638dfca4e34c2e59e7a477d058;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6ecd34613ba93ba9db15c894c064ea7e138f2472cedd7a6b7f1b562b9f9da3c550a2908a2186339ef8fec4731822f3bbd43f3dfc3ae4eb7f60e73957697d33c00ecd5e3954d691b0361aa6aef43c059dbf7ce6510c674c712f76982502bf51ca6cd13e825c9994c3b89ceaccf816e58b5905cf379eadfd42beb49a3ab7bd5d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7daaaa32808c6381b39e78014de93d9a8a32a5a2238381b93159a4b511ac461ddee2823d6a7aee6e743df952a197aafb5e1f1f1bde8d3404c9937aae66cf6f9155b2785a6c6d62235e5f082635bd1dc21acb0bfaee74c7e5027497cbee49a03f7ed4232df1833a72e5ba311378d25cde7ad35d0ed66a241a3a18276624332bff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f06fd5c9f04eccb2a7c60b3b4756ab105bc156aa0f75fb8e0c08681737e5e9b2d88fde9165675da2cfa7220ffb1137c4cde512e28f4f80e865cf4f20f072e4a8ddf239d04bc96a49a781663f61df378c3eb4a4abfa7b304befa4119924b4cd92fa032b488bf84d8bfc4d3517e0ee91d820c89c5a78c5c9f0f93c3fed039d403;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb714e5147989a455c3582d4487fc31245837caa8fa35e28d0ca58c3ac749fcd56332d7ba0be38a1c09b07d064ab8da17520a7f139166101c0a3b1ca19daced356983303508897fcb914f72933d54c81604c96091c640a6d268aa6cdd32c9f5cd502b81cf3b717cefd5041bac84fe23a810434ef12b3021f73c098a3f767745c5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab11656d3f51f96dc1683e08178ba1b0f52954620f548b66c26cacdd666758104a3f800d06d4fb328678c192fa06ab71d776871f30d25db2b0f0ae0e0beeeb38160633eddf6005f610c18dd30b2295358f448613f3d3dca5139ddff61522e5663ac774b0cad1ba08271cb56a90974ba59fdc2684f43bc0ff6d06c1cff56211c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6aa3ebf7711d9265d971c9ea9e1f19144e522692e798b246e34528cffbda8814a838f49a660b05a770071e5c994cee7f3bc5c064d6f34d3dc261bf964515376d13924ac049fb5bcf6feec10341ff3c1d2406336bed09eafb9fc3edd73c92e84da049b75078fd6c3a856bd03545c54ac983069a17fde9b7af96b1bc4f76d7183;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8e07a0527c4527a1c725e4387e01bd1d3d7e443fb8f3f2079950bd5a68d6b9d1dba9dfe6bed05c42920fc16aced4db7a4ad312b87780bebf335d6641b8a5cc927e24f22874ab1d23d9612aac2a066f115502c1e70a7c5ea861d3560caf486b20e205cf17cc5d179fd76e633105de8c8c981b30f1c38a7f1cb873de85b178ab0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e02ca6ed3c9c9f79ae3cc1e695b58f4067fc666c3ada47e1296e4679ed1ea58af4161a79a1f7f8231179ea210f3c74d14e78ac3cdac17693cd8e55ad817cae5466f2ef4091e5c31a0594451c4b937d0d796a94d35d992f42bd3252465b46313359021384806a85fd6b9f47234d2a98165dda9f5ad18d7651792df57a15f2ecc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h764823a157b320c7f389caa54a26e9d70550d92f01bf0f25c4a27764577e9aad41dec491144c934781bb4a4c387ebcabd04cca30bebd65d63b517b9a981fd82d8231866ac6f98fa5c6a0f79a13d50bfadf5ddbb7ad6b1b555dfbcf413b9ae0513ef007aa5aba18b29abafc47bc3c1785ea30c3c107787b555067167a2ddc81df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28f25962df8ad3ff3ad1c5d6d7fd3fc095b58af6495dce8a97024a5a92b7e299674954bc1129414680e3414ff1e73b63c2e69a3daac073a02387136c71d960efb337fc73d067848bbd6827fb4fd19d5399aae03f67a5f5c8f2654fef183ebfbe11c94d04734ad6f202e77f06cd2f556684e1200523443ba1a83a0d22a1eee38e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8a5a63f5f8c8fe7e00fda9d443d5d1a06e4c92ed9883fd3e71876b19eb067326496731726152d25d9d91b1529b6926abc54bf4779aa376947654a455f7ed0c814a3ef20adc4814ad05069036074424fa3227dce53642cab5bee12b9e87ac07415522026710b76610a84df77f0d76bc60fdad1afc7fd83f9b0e56106b960db24;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb45e84b24f2808ee6c61c45f57791b173eefe31d9813d329f1dfbb229d42d43a62c275cd943debf7b27c653a1b9ba217018dc02c949cf59c3a88c43640334b583d96980562d472751165398888e77b38002d018d65922e0ec40656637537a4ee93e3cae51d477e390e6ecc87aa6a991799e7c9eee011a67749a619e63f5cf479;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2db5c492ec314707d9a6e10464bb3a0e51b9dcae753d89e1785cf263e2f166ee44b38baef43d043f7e8a65f5ead16622eff04e700d7d98ce63e949b0417c251f753ccf2f01d1b89f8d255cf4ca5fe23a2497d275ec5103adbd9334503a97e7dec850cc8c0df56252b0932bb2bc943c95b771897174893e0a1687f855b0a0d961;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cf1f2f9b23d34e7bf5fbcb054f473a2bb3fe78e529e815638ba0035dd2b9de39ad6648a111a7944c637db087ede496720c802a4fff9b269a188e7236b5766e36ec69e35c096ffa3b091378c19fce24098269b24e7d80cf86627a3625574d832e3f98d21c060b458d0c51d2c92d260c511f09d574dd58d4b45522f7a83dff69b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h450df8c138ee4973f4cc219c530a60f9c7ae189cae3743521c425a8e7738983f14f3fff0483720f5033cecf1a0e03aac966fa0db12e0082397ccbaec746b38484278240de2803ac104abfc6172407e6123fd429df12da58d855fe72093b66dde27a171b6f0bbca34ef4e192a2feea5a785c69fa1a6f7d647c9ba34c749d29445;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11ee6d0df35714d52291ca34d97ca0547d7b8c26b10b15339593e98adc50ff74c6f6f4c61ff7ba49488acad4645edfb0ec926ad18d0c913844eefcd1679b5ea629eea3d5be14b67dc8036044331673b0361498d3eab295b2724fbd73b2f3630326d72a525adfe5b57feef151205fc8237a9db8b386a764d67c7c525cca8b56ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7969e8e128e830f826bf4cae8f1a45797730c3b2b718af411c0cb03358948e4b9dd875aa9748e3c4096f87c3e3e5cbbba826d13e7d20cba2c92ab9eeada54357f8b8a3a655cf7c78dc2ffce8279877e2301ace83126dc12a6acd9908288d6abe73422faca86882e53ac2fbea3549dc96c7b30c7f52d7209e01f99c899349ec15;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h803be8e1f7dab708290b8eea29b384d08973696063792ef016c0317c42fe09f86c29fc72e2421ee98891c1dc459402c4aa2c1cbb9683d8e42e3aec2bb82f964a57df98d145aef0ff04768b3d53c990e5939abebc8d2aec83a3b4edb5a17f5d1cbb77c74528e700caa91b94de3e4c720e499f43037841fb94e33304eaf2b209d5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1898298e974bbdb17c78ab1283dbf4c942a60f52c86d60f8977abf23f0b1d362bc0b8cb6e44563ea8eaeb81892d7c4a33aae0126a89e9ae7c37d0ae9da03fda8bdf24bde52678b8f7fd7bc8207debbb1c4bd8795e25110e019694f58de4ab81b667fc2e6e6f976b82aef86f10a6e3a0241a173d05b1b0f60680373bafaa1f08a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf487efd992617cf1456a32a2c27957c7d6ddf5a73ba8a4ed94835a815f4afc4f3670d8a0cabaf0f170f4839ec0be165559012c0c607a462c683e0f82d4f6e1deffe5cf07797ac4ad5c11e321c141cd1c4827ab315bf373cdd3956ab197b5940b58fb004b874a509c96bfb53dbcf5a5538164fa8562c086a201621ced60de971c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc27adf06739781240922aeda5b5d678c07c4973de9d676b982de79b585eeac37694afc898599cc4bac37018d49a7bd58a099d513aa548aa472211c99b46392e9ccd59f6f0f5f6e81f4995deb9a3875ae58ed5c4d8d5bbe60cf88721634c894fe6afb20e85f9fc69ee7cae94765cb9fd679a2faa912b858d809cba646466ba312;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32b75b9dcfb7bdb06f776859c44ff654b61a7108e803cbdd6a4a53968f9fbdd991715f0ec4f0d3dd2725c99918fa0414b3ca10627cf5b2d4f2d4d7042155eb50a2baf5aff3ca286e7afe5f29a5ef99d0f503d227477019022dc64a3df2ecdd379f5395f07a4b524b716248978ddc60f1c5c67d68d276d40bc26d7fa0922b5370;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f1b33aaaba15d443bb3323997c3c936c1d3588825a1ee99a9158063eb1f2dca6fffbb9e47b5083db51e8b8d03783a0dd5931d0768557598871dddd7462b205df078e85875df8b7a2ec9f2dc9a4c72277d7cc4258522d28e112559964c939bc7577bd43be481c0573c0d4222b49719d3b2db9f40d32a592266d4004510612a6d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha177be8e143767dde945241d4ccffed5b4321466023100a4fe2d8a01b5ca7a07578b6b922d18c4741bb1c66a021b3f4ea801656416e0305ae98f9ae8c4ffbceac77fb7b23f91cb656f7f3c6e9051e977d18e708ca3641b5bcc270e7c3bba8d01a3f5f54459a53ea415c18b9a6885f01da68d69aa47bec33883e2b7d9f76e2732;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h955397d518fa1add1520d7c6ded9b8630f9ddc0a84510f97477d64d95809c06c46b90e522fcb416d4d3444a6467e1201cadb02cba794919cb1fd68c661c9d6d3725a1ab18d1f6683740f7545c06d7075f0fe739cd61ad5328f21cde06256560b22073450ac5ac17cc112d106e5e37803ae3dfc9d8225fe8b331e8be0f2e12f05;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27dbce2e2f970c6a49a988b1a7579512719da1e93a3bc8226b8ffea418a4b8e0f10b2832e9f0a6e5ee922f3f676449edc3f308012635ce039c7eb0579a265e7195d044fe00cad7880a053a60bfdf64fdda4bb75c79d00032cf23e03a8860eb0b5845c3c823f5fdd0544c5e94ff10065f5e428fe02ff9a3e7869c82376b1c2038;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3fb0af77c0f46af23e2587da57cee67f2dca4334ab69f709c206f6fe0fd340015230a15c14746f893022db6b4d1e72ed963233f5526dc84883a8c8b54535baff9e945f110e576c2c128dc251fdc88672d4af95aa1b4993281d87fe9d516b51fdbbb324f6ec4a6c3f4fbd7d6b630f6a4fd18751536b8a8ced4fed00b28ef5274;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d9c9384f697a1908733547d7b553abcdce8b23b19b082141647cbec187a3f733f81606c6fcbad6393c1ee9a12715acba126e9f98cb5d226917ca8566b555caeb54b63e1c950491e8c0f9dbc1bdc893b1c4b37cd33b88f065f52d041784a23bc78cc8766ba3eabd91e470d03eec20095f3f8a0eccb9041d2a08223b84ce627ac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h324d4fd59f512727aba5b3c87a69171e9bb38fcdc47f32cd4402ccb06112ff6313a5c5f28427edefa741511b45a64dbb5e64a262520b64f3fcf61a3d25e2715a209200f1df63012af89746f7091829112b849037e56372d59c8bfa683da15e4082afb5463a196094565f2d746a7da1f1ae5a7e63a04d9c1da5d60086eddb3a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fe69e30950c4a83187669566c18bfb5bf73f46679db96957cf3ddb3661ffd973213939c3d42c12bc3779a2c7d1bb518c92633c8b038000220be0e3f5f17ab819227614e1bf90e335cdf88b2ec9c0626f5e1d3416d036e780e97d3c1ab61284c4699412e373b2a3c9796633d0bd0a6756c1a3aad565a93b4ddb85cb00cee7a13;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6b2074fc467990c988c41050410f47455aa1f9d77a2e9f2dc605880613a352892f254a61edccdb41071671d87c685e4900384e125fa50ab08d953f5a33ba344c1793221974396f6f3bea8f88cf681e6e2edcc23e1208a3011b9a511e24550cad0f64ad173244f7baa3643bea4616323071140e0f651195ffae82f1e1621a52e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9628cf69858c582e918df58dae789c340f29d699b91317d61fb2e90bb46fa9dcde4e54b9bcca48bbbd8f04b8f75cc881b860e88df1f04dd3d706c2aba1974dd132c1136d1b8f4c03a59979985d8108be0cffc49f9080d4f3a7ad7282c1a1fc82052a866407de7d1b4d7c610eb137af2141fd11836c7b83c6c0c0b05bb516648;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h365cc03c5ea67f6db3ecafcfdc5bb622f63537b78fb7ac01f130ca655555f32f340d4c98c2f104e2342a74137e0955572b0f9c73017d18412117781515e7669921e40330d4a4c76aac5febfd5f1a06a361f4b255eee31fe43c73a92091f38dc762f938c7e06c4ad8e54cb8271f83928426ede305e09506842b834d17dbaa166c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f9cc2960b3b9e678027098207bffb5825b69c91eaa11455dd7f35e828206957efb6d1166b7ce6ffe59fd931b52df9d5748170ef3b6541041f4faa335f80b203d93a6ea085d32ee1a4006496962b3e36bf90afdcbe9a56d2d069ad84ae07b92684c38adcec7690fd05d5be722b757c73b671cb6e2fd8906a35827238cac94a84;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32e3e89107bfdcf53f6a13cee4cc1a898f747a33f5c85f995cb0f7eebcc8b852a30037f490e081f00ecc28bd2c775b9f0819f96da3899e74098f25a7a521ea8e8d592baeb04153327552a879d37f0fa875f7dae4d089012e99e3e686bf803ad10f880b7ce9f85d55f3156ce58a9dbe5e579b44494f05fcdc60a0e6a538419c7d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f38a88baee5c4a55f9b4ead9e05171f7a289d491fb495527eb9db7db21a54038f51795b2bccb80ba371c508c06155a510a7cff739885beaff15b8860ddcbb7cdea4bdaf7a9c2a0e15c86b6e35ee2870b3ba32da2fa81d6a6947610044c03f973869e66e4558ccfe53a8a73a69391e44d2314a47140bce8843477a2e3d31caeb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3479e8b35bf502a39f6afd19806193b731fd7ee22c1155aa4022356716df30a3602b32b14caa22c801ce146e4de7ea4b9bb75a2edf8281cc4332fe173b152a08d3d7d80476a90579d34f57de553db0d0eaba3205f47a35d6cbbf2e00ee1ec53e3d6c3e04d931519b27abd04437c64a56ee62fb9115ad3d5d9d80fc64160cfe69;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce1ad12a7b65511d517324cdc7f0076c38865b4c1e1b1f4a02bde0f0aad9f3d9489ef3c21583a16c89ebdf4b6576f0ab0306ed1b1664c60c1015a3793469bc1598792e065a1640fc2c86afaedff65fa6c9d7c78854d01ae245a5ebb34618dc70547d7ecb9ab1eb86ef70912d1be74765f6f5bf33e8f45f2fe37570c09f284bee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7baa8536a96d5ad4968f04b66720719faac5d83ae88ed8c9b5966abb7b0de85f503cfefc2ee0222c0b694f84b237f7555588a50dbc0321ac30beddb348c6212cc3b454a1b456cdad64e1b3b89b00b7b1cf9c6dd34c34d54dc7c9a75385b3eae732913d9f8b1c125e76e8056dc0adc962b4b1db4ab5e1ac56e2bf0961473e55ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83e2b570f46fe0b7a31e401c860099fa4759912bf2a2395b9bc804d3f568807ad9b89644cb44bac2290f78a6797505b265eb34bf2aa873691b85528d3b960e232ec9b7c0c7d3bd1a7bf63c783311c8624a8e04e61097e75c10621ab625acabddb047a06c05136ebddccc9a755bc25d50c6ae5c2833393374ab5da1af9de88d7e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hecb9b15d88f5432d7da908e9fa6a4da8f9d77e18c4e552ebd1e1142116b74828fc142f39f7668044225b169a22c76f0bd8a6602e55644add6c53b3e11473c442f124be481e8efba16514b36055462c7de1ca49c955183774118eeda860aa698511781676587164afb33dc66807710ac4e8fc72bbe122f068f0ee4fe64d7678c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea6ee6c146f95efa5a56c888d660779e0906b742d6793033ed7f1ea8ecdfdd5a2f71ed6be624e50b9bd254dd1d49455e20360bf290fcd26605e344039dedf55a3d07069c15e030493b9a818142bdb5cdbe92dd0fe03af411c7147159026c6a88e1558af1edc609ab0563cfc5b833917a9922a66bfc4596d21dd3f31dbaa09ba2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h769a53e1372e7778ec0defe21ffbcc7560c7186536834d343723459219039068a9c7649ab7ca3ec4ea2ddb9b53cdf2ad3cba5635948988972d8bf4b36f4e65f6277216b3cee077c9be865f2e43b741223d4903766b2443720cfbbd2f6b4ac295b01f025ae6e9ca1d17fc60fd231400ef0f181a3e8833bb169d6a1969c7bc130e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94f16eec765c015651003827513c0b1b3103e8ec87d50a036bce70d1e9840c0d818b09489286c1a4ecb6a54ad8c27176ac7877f6d95c3ef2f0290d48eec2ec13ad1806a9370c005171830271ddd8750e48597a2f0423b0eae232426f039daec43ee2a7df5f08d4ddd5259e7c20a4dfd3f99b4121129c903f462b7e7ad5f4813f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdaaf5715bea9bb7d0bfbe0dd414a6591d80571bcb2570d2a4fb285e3dc9ebcc8390fa57df7826ef5e493c4a0661a8af014277fb734383fac99313a437f8559c5cd80782122a43fa9f43c323f3076e48115497d9e7f16e3a8da77743c7b97abd6925489b66d4ec1e78041b01d948a3badc526500fa083c05ecf74cc232a0e6a90;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1911b0457b63b7d45dbbc0d54f8ec9704801e44229e38cf48f279bca67b62a6ec6ef2c09ef6222ef6e1e7843cb5fd9868f94f6ecbc724620c62c5378a2a9547bf1073eeb774ea263f7c2c2f888ffb0b2ddcc4960a007a62830f2e22487be1a054c0cf061069eaa4d41c5a27186d3e0068c48a4fd88f97066cfa982305328c06;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19ce0fd58bbdedcd0fc194c46b86b1defc437877a92734a723239e14150ff1bbe300b34590e36ab27f32da6278432701d6d9c80059fd74587bc48a3ff6237424e72cd0af622cd394c6900f5b0340d10d615b540ca619e4eb43c684d10cfc3a45aa00c636eb645535a21a468ff441a414aab88fb51e31a2911c17f2c78817fad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd13fa2ad1a5fc5917b4ceba6424e2aea78db1a46b50afc2854f0871ee34ee1eea6fe450a349cc04745e2f744de9aa5e81008e60e5be71f4e1354bcf8f9d6fcc112aa17e923e8da6aa97ff90a0de0e754ab5ede50b8e9e2b088d7141675ea4dd62cfc12b5bd6f7018ffd9032643bdd2a737f65a1a59593016b13a313613cc74c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42a9d72dc03abe068821702a405d034a611f15c4ba40e4d0bccd70786ddf47dbd1f16b7b45ed7110f32a32aeab52a2f8e77f4fb1cb49a6133acb60066fb1dabf84623c054413494487ae99254d9167b22ae5f5addc00ee83aece31c407ad21e4267b496d2673c42a605b38f64aaa69be89585a0ee7dbb2124a2ddae33032edcb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he95271a891c1915f2b368c8158bd3b90746ee3a1663a0b84b592fa5189bf9cde09d6e433d852a127ecc1098c1c69982d4fa690bf564e562b32241743080a2677ac7c47b226e013f8334a16cc074a57e1b2d1a7573851d7b4949bfad45e99e9333a9d6a1337df45a2d70c26ab8aa917d5232aa6a8075eb99062336c0697226be3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9302f7f8fa7748c39b55de863e4915a54254c81b95e71b69dbfa1ff1a637fa89a6c2f9ae87e0c679b549d2d4bb63d87ac3a0b8bc1ced07e9a4518774a20924929b982ab54b9b73fb8d5ea1672d77196c99a9234417a3c3408d50266dd1d93b051c2efc6a50383db375f880947de60f2ea240d6b189fff4b16983f92012c677fe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf55775ca105e1f82dee3fc1e66c78ecb83d2b60566cc9fc67129257daed3691dd167f17ed7cd1c68a23b1c6cd133f9f155f70ce094fd19a11495f4b917f140f2d4316cb06a6ed427512fdaf52fb8f1643941e372f3cdc7a3141dd385a8d2f4283d5b5038fa87a4fc43769adce607d2269a87d7c4f43ed0fa42044433823fed1d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd77abec4859b1aa257e86f4e5ef5eb3ff20df7f7c8526a3947a9a1e728d773e669c992b1122dc6bc619a5eaaa893ed69043024319487365d57f6d6ddf1419bbd8574c93ed263366d41a84a80327b9c13a08ef782ebb2513688d4397436fb5797fc4b87362be44860ae22972879fd8d43c06621bd15fc0e63d1116f18c28ca6b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he78eadf3ecf20d11d8804800310b592f907767f750d87eb262234715b677bf4a3c591f326d6b01066f2d737020ac7fe4c4299a1aa98924d2710bb13c8789aaee4e52001da8b58d0d7cefab36a4d1a753f3be05a218b247ec51c590bebe61fdacd6c9e67e16799b48548fb6883239910bf752b278af60f69e0015fa2bee98d517;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1ad1a8d4d99dee3626fa78b248163bab7253b7c962a70b3f50642e7db6a983b2a4189f4501a988d560cef93d7c121deaac0e0052e5a0bfe615fe0d29d4576bcedd1dd29cba670e264e8e4e5635694dd5b7384d2d3296781a86f036d3a05e5cd2e65f7f61dac91881194e63303d4f6f9359755c8280f5a48394f62fc358d2878;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h831eecfa3ac4a8fd2a6ceb6beeabdd0d4abe8204fe56ce2c2cbd134e9c986f19d451367d128eb2a56e94ad05744b6f16b9b67e0a627c6a99b0b0ab6dbb2604012e4b373a0197120802b110709c2e4971435badc63320830cfea82dbf0c56df2e4244b82f4dde0513810f77f823afd18308bcb57cdf04c6f3464fe28a853f1e1c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a4bd8f9046c7c31c7e456189383e72b0163fc362e8100dced35550651d5a042cbc28cf9238aa824d846b59da43195d2d0bcdbaeac82f69786d268feb973cc01f5141c0ce03fc37b9066856f95052098ec62370b8c10b8f0a49ecfb95de94ff55b49557284e71e9d22db6d483424c1382eb785e4ce1fa0ab8defdd3fd09d42b0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21de6ede13572b2e07305b3d8ddf7dba4bfbfa47c085f63f23974c036d0debe08da5407531a60cc20d35974c488cab31575418dd82c4bccdf366b05a7e1bb72b56aaf3cbb875cc8058fce5090c3349c7fb8e04708bef0fccb1f8330dea1c8a110843161affb24cf956bd705cfa1ba54ea2018edce70663be815865b23edb9b97;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ae2fb318f2ecab093588ce781b3e5a93074bbd8785dbf9edf14a4606d1b47ffc2af73755aca1502921c9c69dc78504074ab2c75defcf353a25e6d2b49db8f1a754f9d12c7ea4fe866bc1e882c35e66b226a47870f3f07673873f65acb330ef20ccd24ad02dbdbabdf3c3d03983c560a68178789c4dad1ce383954a6bc103f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haff81bf6408fe1972bc2984ad0888293facb176536d323e547068c44afb8447df8adfea2db0806f43862835371fc60c366ac59d4a49e9ff676377f70509663abe6daae7b42d36b1c305b5c9d5d0754d9eb6627eb41712327f78db4b34ea74fbd979060e161276a6840fb1a44970d22a1c403626e4fa08fa31a77e1adec7c0df0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a68eb9b7dbe10abcd1c1cdbd907d5927f945247159bc17076fbde3d5c84bbcede247806c118faafecaf9c2ed4bc40d413f23e5c63bbf6b5686329ce915bc2c3a5ea13638ce6ba433ef915ddbc4f945c7b02a16609b0c04355ad5c975340a383ae7a7091885ec92a416648e039ec7b3527be7ffcc2c2b96174dde820b561b230;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf2c5557c08f7b65c240410f8b3bf293bf269b0488c241e2f0086547a9bce8b35727b044afc2e764b89e34bbc2511a2698a9db26a43a1a2051ca66481501b897b9b87842cffdc3ba2402dc35c3077096f2bd414980d58ddd27443476cf547d7785fb6fd7e26e7508591236fbeab48c6ecdeeb973cc521ab28b9cc6e172e52c12;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h418c818adb6c3703c9b4d4f01b2534eee89b39a296506140c26a9214d55417275ed1dcfd0de1e70c4c8fa63a8d5dbc42256be87fa908c7967a004edc4248db978381b423e29e1437320d43819b53da2e52d7e632a31a3136c39c0480c9a6d649da0575b73c41a954d5e204d1d35ea683cbe7c87eae92c9b1c6fbf10d823e0c5a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h407340f463f214f6806b717a2cefe9979fdf259c969fd12c5da4ddd05b7b15fc686859e3ee7751adb7908fb2b147e73d085656ba358f3e5d09cf3b4f4c5b4f1a78fc16afac6d1d8afb9cdc195c3902c22717ff1a20ee8529a2a32c46a89b6bb9ef6e34f04d04872aabd37c1f4076b5ba84a66d2011b811e18b0cdb71c376e3ac;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67a768cce6c97d98e3f6e317d9cb5f0e7f9314a0db83a7917a6689ba8cff76f11ff9f00cd1f0556cc048e126a67b34d7d02944f1d0d366c6f459b5921cbe768b932a13bc5aed7a1cfb2f19a01a08c415a3ceca1e0ea9accce9f7425e43eccb75dbb3750a4235e2dac03b7d56859e1494dc79e897f8893b4497ca2a621aadf040;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h800c9f194d4fe0b09f421dcf739471b3b161c24731405a948ef4265797b7498f1c262c140a26c8fbecfcf1b362f4ef8ed029004a880984acd8a987c07874ba71acdbc3bc7f34cc70f20f985c888c50c9fc04758a04acbca444ef307de067485c8b4eba77286e82cc228b823c75106efb708989480b91426a989c82676c0d3e3b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe025b8a4ac049213ae01d17eadd469dae038889d65e080582d1ed71c094d549894fb684584b130f9dc2db3474e5b834ac9630f1a922788fead0f065a09b37faa25756f4a0496d110c966e850a23b5d21bfca02b37940f0fdc3fd62a0fc39305a74efb9313de4371cf917cf6f4d2bb34b817edecf6a2f93793e1e5546b6c355e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h569455ad5a8fc7a83040a5ebbb55754b13e9f244511d20a6e08dd17d9240079104e7cc97747d1f20b779709daaaf21fdccf88e64c09643b618cd79f2c2fe8f4795fbab6a3e6cd05a045fdf6dea7d0190679cee58f1023bceca281d6c7393ab8b69a7c39c7d6c97239bcf6b1186ea0709c2399d0672de5f1536e8d8f54e5d05d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b52b28b22ce7fef9f3eb580071a8b888d40b7d6ed13a46090dae4d612280c4118bb6183e8d7cc4f58f33b6cbf9d30f14d32b444e3789a95a6cccdc4548b3127e2cb41d9d08099bb83ecc3b367079070939f5a42ff8dfacda1bef09f7ea8a6af0ffb5f14c3f17727da889c2c4f54d5e475f1331ce4f91e057ad4244d993e4263;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h330448c855ad3ae54c57821bc0ef5b772829f7a620ef4b9dd19e09a66e172ec579cf75bf7096b09a00fb29e10cd47fbf9c3e8ab772459402e45c1d0bcd7d1440dce08704c483a80ddab08e78a09ce6c55f51935f32b288197aacb4e8e7926f68f08678eed718555b18ce4ba572fb817f795b76c6f5e5862e4797be7256329234;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdbb43830ba20316e5225ef55117cc13b6d5a77e0a3a4056d90bd89798ec4eebe2e414f2e5786258421094262b30b3e758c8b1df821c8b9c5d578e9dc32aa4248944ddc0ee22b9c1fc16b8eaeff8fe451025acb5a5a7e266f8fdf9625fe8d5e55848470758a8310b0fc225dabb14411233eca1422438174fdad19ab2b3eeec3e3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82f979380f1e75ad522ffa634d19b8d905fd621b0d29a2cada0f8fb0c2ddee079162ed11317e14fb07bec9e54cf76f506c559fe52848abb9bc3f2742f1f1db5075e09ce8e39ab6d296b19a801d72d2867fff2da048d1c245ff01d84a406c74b69c9e5de9cd89d249f0cd365e24b7b62a8e787e5e99e3f3d1a1226fb5950e7339;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h895b7b8824c4591853f6a72feb342d1bf687c0da7400fb6e1891889e8c089daa7c4e2a27f49bbc26e5fad0e4d7a608b36be25c4110ce7ca240088ab42572a781525bdf3a12feec38089373414baa1c96640aaa9fca732d1d30e44f45dcfce93ec4e6b40a7a9abbf1def518f23fc3972e6b580d27675dbdab4f27877ec3920f7b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f5d15d19d723d51979242c0577c24804f3972dcd19303ab8903d5d2b352f18215c250dd9b73cfd93f4d15f8d6159b0e22f58f14891ec1a686afefd720d3d135deb65813e6b3d4cf1d624f112cb6a02642b8a62a77dcb0f1b4a6b3ad11bf9d5b50ea2886e8691a49ccc9ae23b7fbeab84eadd9ca947526df203b3b3d6d9a0666;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haee848fae05632e9127293cd5269ad12c17a2e373fa264e27ce292eaeb289a34d1396d7332a936447e59c2074bbd0710539410f6efd431e3d76d147e3d0d6277b69f8aaf5443a74df565dcf58a32bde5cbc5114d4bda842b54a89996da7ffa994a77f49b36454d9997df669fc1ee2b9d98db9b797a1d3bfcc5ecd605f9d18a65;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdee3de1f5e6cc059a08934dc9dcaffaac85c97958c87bade64b3225dd2193db9d476d68ed2c53cf5d892065c875a6c86d7587db32556a8fb4c9cd34dddb3ac1a51b19c170fd30f26435f88c138aeb481ac65d42d65273b3cf5c5a3d72c4462d8ae2c7384821cf15b2552c411cc11bfb6d39fdd091ab890d4d922db286a74122;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ea1c679528620817d90297ed4fbf0be15b24628436647296a1485e9c43b958015c3cdc6840cc8394744e8651e18d6b89a1e25a49ec2b181b230fa3508ba12b387862fdf626b6f856f39d5cb43738b5d29cd6f7133678124beb43dbc7cc8a955145610b67c3d3edc84c7c3fe7cd0a40caaaca85e13dd1cc3dc457f41b6e8fc8c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e492446561acc3b879ae3ce98a25e16c6c079faac34e31ccefaa27453bef81ecaba6c3743f20b05675a0154865d76169aeda1d701614d5c14beaecaea48d9e742afddf3ffa25556c15ae9b45e5ccbd3ad09b2f7485ce01881869e7cc5dc4019083cfc28d5418587ce4a41fe3363feae7247201717ade31482ebf923a5ed29ee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1d93914bba1a702442974ca3411ff150ca2457c0d2c6e3b26694537bca9cd97b2cd1a6daa0070ed70646abd2a82896dc8ccaa2a3ccbfdf749334a863b551440a1eb75ce6bc1c270e9334d6e038c3128e8050b70b654de83a2c6e41ad7020ba6e5539da4d920acf86938cb2602448c026796d579b06285778eb8f17bccc0c1cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0235be165692fb4e4b3dfa7bd015f9dc40d6d3fc5d23c60141278d950a922d1352e7f720fbde7c5406e111108fa40a15b2a6acac06ccc783da5bdfc9da8ed4087914ca9fc4b6d9e641d86e0942df2855b33398d3d83048a1d1c709fdace9746985a5774090f6eed1340e431803e50049174e01776d20b3be63d8cd07ae23170;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d3abcc38e42e18896a2e135060971ea27a95d42191c76a27571020e2df29402d3628685920483d6b0bb2a83c8ffeba9b30aacc3f08526c7060707b9a25da9964121d68cd9d4ed00ef4c4c6e36094e9ee7573e3eab7a7c2f9197926abc2d2b85afd7b58f37d1e9e12a06a86845ed7bcebf0e6d24bd48110b42fdbe568ddfc88e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f4e181371ddb15ae756f062f754ddbc5dc8605dee79c46eba39ce70d861a2b6d4a2d7ae0f3103dc38d3df7883f766cc415399b8a6aec63ff2ae2c6baea755c5455f39ea9c095070dbbb9685b66d7826dcd37d188586fdee2d66b45a31d3a56408165fad7bd837dcb6594954eacaff2112b6b7686f0c967bfbc7148af140c362;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ff49e0115039af47149831f2728e0049985e98178dd550c491c0649441379c5d0b11473c61a10ba209409042c27b83b2f372549efb85d4701a5abb903a073f719ef9d4c182e0cc32caec697cc6913e56235cb4e8b7363ef8b8655112a483be524fe49d9c906c5c9c642617fc57bf6607775f4a088129cee09960e4bc10b5b14;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10de01bccf5e201c51d479ccc47fbc8ad0cc0c425c5f32d72b6f40003cb13e8178348c18f678c350f67e669bd5963cf3d32f7af31bb4f8cc9ce95dbe6593a999bfb40deee42a85d91bdf93ea52344c6c5d309e38bd8c2fee862f1abebed52cec166a04793a3837d1e4d6e52e0638fdc37ed10c80bff6067401d083e047b95fc7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8027f6116622da1bffa78698675def8d968af912d8051635b58d4b5e5eb112a928c90994f01bb71371928c5dfcbeed3057994180659b111ea35ca8f590f3ec28a949521b4a68e6d5ec71b5091d0b72c60691d229f8c52db5af6556590be111269a9bc3bc80513e3b4c1f06f3e3b175b0858119f1761efdc05c3f797cb9a197c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1f30b8c6da2a76e009d9b23df4450e6e046ec0dde98958e9f9c4f6d6ca663ec002d0ac2266de7f3d597754af6c0e13f804aa6e19fa1c380a56f56f2eba9fd2eca848e1d8f0722c3f9c4e2ecad1c41eab169cabbe0f7646ad3326bf17014db2e08327eb3014e6c2a4017c8e550e6817996a79229e96a0d28c103a34aebaa7109;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fabda5d0891fd9acc1acddb7ca50df5afb94dcf77e541533e2787b033395c2fe28795698784a7b0125bd15fed32fb66d90f71169a9e090008104e4a6cf4c5860b54630696ab33403c2ff8f0cc537712b7220ca7dabbb0d672d74bd2b7b753fed4e995272b5987bbb66378b14b026e6572d3141f041118df6b6c01406dc75671;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1342069e80da3bce538c7a40c188d4fce2e5304a6cdcb4896b7760cd3cc48aa50c080d5916489fa3ec68ded7edf8f6cde7270533fb73d464976d6c8d395617651ee0f485efd7f8bf769afbc77c1627f2a0791c8eb8578bcf139e62ebe7922920b4b195e97544f49e449644856a00ca232457e68e41be4868eb72d6734154ae91;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h959fe4289de3fb811e5daf489da096c861cf1d7e186f18ea7b1c764644f1db256dc8b9394ff6f25fcbbde482d596ca1d7ca9d5f639c31a8df9f7eb1e19d72b3c8eda4e0cc362470826b8aa0d0b907dfc7d4f6409a083a1644f168c2239dc3bd47d6a1e5b00c4a113c50ff4db00611fc05c50ded38c2ad0a425306cd536a65565;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d5468abe54fee5dc17179c86bbf9208525e065f3ad8a50b1b480f7f119c40cd48864dcfa363a654ac818a19d0d2a39ff4045f3402a069bb259c66bc01df91c6068d88505b4a489954e2d372db488f2288e6d62f938d221a479e54515607c9f887ad1b07cfc974596b33534e156263123cbc6457a08916a7471d0d53d2c15c09;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7282c4beaff071295dff116493f9f33df907224a13e14f0e72fe8e5e4342fcc243971278d3e19efa83c06f2b9f73c9f61fe512d8a48379c602c8d15b78d9dc2f9c30954f28154fec8781343a676efeffd4ab772b7bd605258d13124c6fdc939a777179f034faa29a74db837acf31810d76f3d1164c9ae3dc7b9e0a8a486906ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31087ad1e6a2f4e95cbbbe7381e4fe7cec105ce0b80d1c9c966b9c27af1c16d7d80614abdcac72040c511f7d3ac1c146c5dde844ff7a321718079a3dfcf011d377cdee7ba794c70a771cacaed334367ad5ffd83e4c64a441479943a61be6d06d04ad55296c1dcf06c78e69da2582edbc68ef2e1043fe1d78e9a4c93705600dfe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c1f7b248521e7e537280fe6eeba2192f823743681167c0cdd189014de1eac827f0fb6b181086dde0526f47e2e4f00450ad7f71a159275c22ac94bb8113045e42273fbe4f41a8e888a95c2e45f8ff4ab9514012eccaec1ecdd03bb817948d65c09ce03177c25e32e802c85da39debfec43727273258dc33355f8a894c0c224b7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h77ea1dbe86cead7a994691dc3410e157c9a321b14f59a5fcf2bc7f040ea1f8285dc0c083e2300bde19705f09317eaf5d48ff042000652ecc7e59d265c4370da59bc21f90f8f01a404b400d30bd6b8a4fe332882ffb456c240308659c0a29953e70c3ce71db858dd7ebef608ddcdf6a77feb97a5dcc5707f2aefb98fe87ad53f7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37b203b597d9ded2ebdb3de979b90f0c1bf7b580b0e645cdc398736352f2483f1104fb1c5fabca63af462b64d26b2e40165414d2b821df36f7ebd77cbb6bcb3565b862a064d218e87be673ee56dd7bc01398e3b002108a07266e26cb0547d7144bf741f4369b1c9354cf7575080138bf376141b1a3ecd9dd3afac11ed0dab07b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he41627636b540efa4991dcee68119688192c32248e492c069548f003a2a4810d8eaca42f4204a6cb566bad5df8992acf12c8a19785b05000a23189cd29cf42a597b3869303e512228e7a995ce6455f346248c70c25d42b7272f33f368733ded587753f1b94bbb19b4bbb3a94d2834c8f19bb8cb384102aeeec01869e39905b3c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24d1ff7c59c29e1bea219d4771b543dfb6ae1da6d54601c07949ddd122e5f71c7e5db66f8187ef109033621740d79f355a93de33dd3362810446f31989a5df4af88c1be238413cc13fdadc8d96de57b265676535210ff4252189f1329cce6abe486ddf5d4bdba0da7cd4508e3051434285eb40debdb81e113cb8f97a6b4785ef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f7c93299e48e4a857ccf759690db58917d6679bb18aaacc6d322286e3202143a6884838385518bae17259660cb9b2d9cac8e01f01ed2816ea572896155d4d34bc4caa5023fa1f8fec46353e0978c1b262f3f353b2ac5baa6f0e24764f882f8648954b611fa11c1d8db8374b5ea29431b12f1bbde9018cd40b4b42abdffe32c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3007772e8574bd7e66754ed34dd6e220d0536ee9855135aa1a3051690d2a44c912b693d705cd1dd484fc466e5484b6280f28e1630584c6e799a8578a30f525fee197d4fa61c26abf7022b4bee7ca92d27f5df3817719cd8d8126f81d51f74eca5c3a433026252c632f9cd910883d92c0bcbda68d2e9c1d6416e22c19d872e4ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h576aa30416aae083652e9a98063f5d7b3a14af64aad9d518f0fa89b8f38fd2099ea5a255dfcf12238fd22f953ba993d0fe469274f511a047d8ed307f0e4fa9adf0e045d9fbb8da964fd0ec1fa97a7d7064127ca177eea7c3bc4362bc5ce415743c32ff15e15e4252da14d201f4cae161abdf1f04ecac8925f7f6108307209899;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd67ecf0db43ad4c2955ae1bb8b4682b3e5d0430a0cad5a617559d378345af0661929748f4ff884b129405bf445eb3f8ff5ae844991344214099732aa34a0091406b36396f686c97180c2a17a45bc5d7f167f4ad980f24612b98e179b1ba7508c386b1c8f2fcb0f1d5d72969fe65f08c3de52093327724e84340ae1d39fa29e1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd65deadd6810d0454ec62dffe19797d5867cf68923688acf829d637f01a6b671c83933cbfa6ad6741c6d586cd786419e73885d847512f759ef4808efe87c7bc1d428e459f4b1124deff83d86e6a49ab658a738db50b506bfbf4cb9559a2146caf88c72e87ddf367af82c9004cce3a07d8d77c9e8005094d9372cf16dfdb7e8ea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bbbd3a6e6267eb94b198e61f770f7e5ac32da4a132b0bf57fb394290f7a8a7dec45e726f1d0ddbe7a12ac2b383bcc26795bc6dabf6c49c5c833fc7f7ee6a7a13963c5e34da64af0904e171b9f60107b7cfa162a06fb08c86525f38bf405cb8b16579f8c5060c68335d743b0a63b4e44ffcb4310c72f9c1d6f06f9edbc7e3a08;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94bf7ad593166a5d31f0538e71326babc6cbdf7fc940548b3877426369059bced897a2d8239e3ce079b6b91719b3e96841a1a0fcb8b47a5aeeaa1d21a881ae9ddaa59616ce7c73aae41f68bb295bbc447f6d865cb7df0490d388af81a8ccdf407260584541b08c0c304938cc47ca48f0b3703ceff90afa09e3e0d2613bc688ab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fa1b7e07a299f0b6b3d437a73dda120afe152b76e9baa3753ff86116c47ce31e8be2f631eafa666435c116b6c15ccad501e720f477f3cc9f9b3c988a41b82bb7e205c02248b3f036906e7a5cd500d5ef8393f880edf121e0561bba755069cec161775bdfa6ec75d390e63e68a01db601defa888f44463e949ab6b8a98d12354;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7822f7b0397349b5186baf3184c7f2c9341a6c10c96db8b7298b11d1d762ed1aff4ec87a2e63e161cdc5cd42399751216566e5ec04845473442c76dd636d03fc4b69e70ca1429e9ccf2fd5ef73c40b26bc5f0dffff145ed66ee79b35886d4156435ba354785f409815c73c1a7bfcc5df8407ae7c417ecf70ba9763939db51786;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87badcf0e6bb0fb9eba551decfd5d45f960239308de3caeeae44d21a858c699572243d213becbb6d221d55b76ae79173c2e9c6f49900850bf29bae7270e2fa7386d55b01c6dbba1de0ff7eab5aeb13c68093884183b047691380ba30f428f14e615be9a29b060490afcd4c302116f3cbcbda1597e70fd7d461a0eb937d6119ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a668601ba5590083b0d9784ecfc867e547ce63aaaa2c424cb482c5269cc1313816b3d138eb3e7d28fd0dc79a21317b58ae2833a89bd585d9b50c6ff28f24f942952e61a7e4c822bfa375cb3c65e1fdeb205a59aab352b35a64f0fe61d8628808bd28cd63e103408bc40b8334dd9827a1c1a2a3c14b3d2e8fecb1a6a9544b0b0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31f06152a23a5e3aae0283e0ffcecaad9dcf7444a451b1f210f399f51f64a0cbe917778b29e363681d1d54a5a45c251248b2d8cfec44a08e8effb3ab0e1eef9e30135c455c8c5dff2ef16cb5c1d3c1c7cbe4cc8684f50b9f54a3fe7d6e27b07f6b74b62f4afcd11f1558f6c739ba4cc52459bd759f67399df8c9a3078dc01b08;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda792592b93405fa68dda1bbc02b02cd8094f85bcc6c386fdded44a65027424ec119f1a36d463722dc53b9a2fe35f46e0cd8984c6130b72c884f50d49caec8777a7c04d559fe6f4797b0de7de6b5e958ad8ee69d28016e064dcd897884b5b5cb46734309e0e382192fa6763e8aed805702b4ddc7675adb38830d3db012930d09;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1469bbc724ae5a7e1d1c8dacc0d6da2411952c25fee715212b321c9f120a8f79b5e92d047adbe35ef5544bd062709777bccd17aaaab683f102e0b4c02e9fc8c1593d04b58f2a880b0b7aac33bd2a7e1e0a325c90ef0538ade67974b7bff8f491e95a72422ca46b633e9ee98532ca382dcf2f1e9196172d9950489be18f21e11e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbff5bd4e26c2abcc592a9fa5004297cdc8c55de0ce9d6597928989c08d20330cbbd93a9b9d19e2b1a08a7a47bfcaeb9ea9e430435c0369803355c66e224c5e8e81b1b45f81afd230131a8687204616e54691b03f8f43100e2d2e3699e7020f153325cd04adced6c48ac15dfd192432d5bb9f81ef06f6ec3bd0c2c2e9ed67ce36;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefd4b8e186b9fc403e81b9f86ed50fccaa476ce478556843ca0d65f05795f1907883d00e70f4e784e198ddc5a8ede6cdbe62136255b6b7c84683ffa840d58b39640bebe0b92e6db234d72f41b0574135194bed70b365a542af12e3e144bae85a9658795c1c50e56e2f5ff5a08f0d2f8a72e0cd7d9d4b4a9df4391f722fcee5d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafd2fad0721108fa2bf492897d2dd910b234a2b89420f193ffd4cd0cb1a7102a8f3a991cc19323b11c3338f9e2124045b6da2f2491f38e919e20b5d7f424531ee9456941d8c386887d0e72b38b1fa65573264c287908ae8d754344223565b5d5c4656e975081288c859d85275dc5abdfbc21c0fa261287d9c3c5229c0821e806;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c554ab0bf98ec58ce3ea09aeca8454c847d6126cad4215905424b362ec1aebc0c31426767c7311ca788156bce2c821252ceba013bebaaa74b94d8e527c2ad9fc4a15492214898a543c0b5249d87f088b976e850265b4aacfcd824fca2948c1ab7ebcbf69bb286e83a6c3ee502c68a022f05640f9e956317c1a55287447af3d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f208da8c73395e153a7012924c8758f6e13636d65e7ed404de49e7baa077db3be7b65f361add1ad869bdb8fa86c7b27955a84ece632616efd50701eccecd1f2e6cec9c29b84790229956e30ff58a78a7def2d174cd3a093f9447a6ff70fb64127cf6be564cd01393935b16f1a95d6c06e06ebcb6be28230b766d1fb17b95706;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f3d215703c1c87bf7d5482f8db5df6816172a7ee3b46d66f406b071e933134b91495c83d989be1f61e027b69d374302c0b90ce64cbe4950ea613790071ce49c4cbae217c334357b323387876e46dd8f69d2c1af63833c30ec489e0a65b457cb678fd6510207092a38c4aab94ae6a05382fbb05d7f87cd277ecce87b29c7017f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c55dee31914f2c4511439b2478ea43270d7a2f41d375910995936b7d2e19be786b840a4e171e70877ceee7c78829c287dd263ad866a4771896d58065f6129671abd2f985272ac14d42a75934a6d06e9d72e2bae9f998a3ae5264c3321eed18d2c6e2bf2ff2a947b494474d74847e52af7684919ab0bf0efea6fdbcff4a2bf36;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h793731646a70d34c45d888f9aea3e6c8e9d4472a0b96ab3d97596998d605e5a2d32cb905ce31d21182c1d0d1103f87e8c0dc875342a21a2a4780951db67e23029d850914a0285df1432532a1d95a0f1310345873323f4b3b18a172fc255ce3f44681f74fad4e300b3baef893e6a446f28be5a8aebfda93eb18793ae94bc120c3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a037ec794963faa56f3e3a5bb4e11dffb49bffbde81c247ff1598f26c0abf5ec37cfd87987539addb97f13d728420407f63259672a919ec10e2e9caf61efc031200237a4c1b51f86a9f1336213eea6c0c26b5f080fd75baa67fb0f112fbcdbaed1ad8df4cab6606b203c6ec1b4427a43cbac2e9db5a3f97fd81ec43404c724b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49a416493bd3d4d0e33546d2b075e0fac0a75f7edfb35154c124ac16cec5f626ed8f481f09490be64ab7f2a72269b85349b3419f2ee72b70e72fdab7f68d93c4ead00c0730f2babce34c9f40063a767a8d6037c9242c5d620cc2f90245f9cef09bcb3ef02001bd58657d9b40e8f8f599716e15bc955317f5d4f565a2c2e0862d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7dd7e2e67721de4e6ca1b9ac142fcf7ef6bfb7ed62336fa4227fe2cde26444a9131e204e06c061aeb1a0b99099f8c4f770412fb0ac3b9471d00d88b927c17360898b2fe7cec874e5239469e104e4f56c75d764967b7a82f5b66fb7f74772dedca294b21c055e40183896a5c4294654336ac35db7b48af9e02bb09f9119f6cb04;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2b6d6b473eca7dec9a0890c3e91bab989bd287e49fb9586ff97fd2ee161d5f69ca144f392ed401347d0f138c67179e89071e888da40567bfcb504a4bbf2568580192e0694c329b2d4329ec89e30dc2dc9af5495620e643824e7954cdd63bcd153a6c33ddba26ec79419488b722d6b0c944e55a296ce2eb42791e955c94ff451;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7da56246c8d11bc4407239b57d2896e080ab71268e47335c6af56294dbdc546d3ebfd2ac0bc4b8ca2675a79d501e94a7bd0b2d985624e2a76046c93a2c9fcca6c3881d2b28fdb6d4e4c49caf02217555bc3dc39e467c7247d2c7631f8afc1493397353f54284cba64934947543ebe7e79811a12aad7d93cfb3c92c4bdd83f49f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h317671b2fcf9dcd2279580a14844bbd2d6456ee8d1f26d15794a258f5ea40f8ccc3bb34f320b28a5bfbccd0065f6b1755f4e06c84b138ceb3ce00fc680752e0101b19230be73270dfa4a27c31397b281dbb6abbc6471e7674e12a15b3cb4939d3f7658ac90369be15351d9c6002ff450123969e38319c8ce9f76e116ac6018db;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc5b31bb68fff16aa867281c280753fc47fa6414a596c4fc00558d381e7cfef43f93f4db5e6cb6efb0e7c06a44bb8a077e37723bd85dc36aec477bbd9344768fd1383bb3d6c89e3c42ffdb20ed38f5b3fb48772f51eff154dac40596616fb520e73615518b45fba0300f6cb94e2779c8c639caf5267ac45432f9e507c3b26ab5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c2b51ad18112f285645ce614e5d683dd21e75d2e6566635862e5482266863c58dc737145a51fb6953ad19d1fc2327e5c333fb3f341690d3ebcc6111e2bc2675241f6bf7e5d04960fd8fc26e3687a6fca57fe6cabebb993eedd935f715714d3b05905eb73fe4006315785aeeedd2be2e86a77d2453d4558600631fd1178e1391;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35b5932c75aa68269ec0b24109e6949feda92b9b63318eac0b3ce611742be8c6b9722bd36e6d80330942c56fa1dac380e3a6f5033a1b5ea6569f77c06ecf1630d1748e6cd925f61d2e9acd426ac7cf1c5ea899783d462e7364f308dfb85d9e172241d22b294b71b3ef63a5b8ab6af78c35c1bc57497e68e9505f68e987564009;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4e84839a13a91570b06b518b929c5f39fcfc28a7e7ccf9eb22f785dc6bdb03288ca4c92eb0ceabc9d57d5f71816dc20f8e7b18025de617b7ebff2e804afcb85fc5c3143bc6ce4466bba8a08814dbe4f410344f012419be1e2c2f80003ca6547c598e9f7b66117efc8d6bfe2fc2a74a6e72fdfee48b905da1bf71b36a12b3e3a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha811c5700d389f3ce83a99a5b551c8e5e50dac97c1cfec894fc813a63f1cad77eaf64d4083f2f153e1a3efeb6c1f9de38a2c127b4c45e4e4553eba2ee93b5c620d0697918ba88465cefd8847ed8171d5724a9fa5492c89410d50acd22a3c0765bd9265737359c6cff8aeb90fa8acbd2ac700385caf85fb828855053f77533840;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5def268a06000fe5df386c5a293d99b4f2abab968b8f6a390e2f2cf182916593d24d03ad0034b4c47d1d35a629567625f0234c2125c5ce496e5e8f3cdf5b3a32eeb17b204b5b93a5509119ebc2c33df2ec2c33a10b812071e1d73be912e37bd48ad3b483e96a2a65f33436e5f8d2215e5818c04d6cd6385981b1e8aabc6e4c6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b694c2cfc9d68450a6c6d4c3fe34cd5ea79e26e74f00cdb1054a24212871731e5903390cc33b41c297481381009e7bd1257fce83c152f0703dfb1108166c8be8b222f82d5566b6183c32a0beb950141a9f123a5075b746ebad7d33c029629e7e16d3209c9bad98ec6f9edc2aea38689328fe81e3668550754745556c6adbe46;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f9a5293db92124900543e976562074cb41d01485c684f98746a7b38b1cbad4cdb0772f0711d73bac13c953c32d9c735e1eeb3f6be5265bfebbe892b36396e911d4f9ee921119db48558c4dca14f37c881c57c6c0d60bb8d7038a80addd849b319a6096f102f7cae9091c2a7c9f1d24d3b591de44b7b2d7e1676aa85284dbbbc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf08fd0ce91d418a1a9b4dd2e3aff0459db58ab48fc559c2e64b1a380c312f3b870fc8c7cd5e95f4c3a03d24fbe57a88f65381ef6840e11339101bb4b838a58ae89eca5024f28631078097bb9cf1d6423fef352c3ad86e748fd46daaf67da42470438e705ce223a71a90a01167efdaca4df3567779aadfa4cf794a67decbf45a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf43ea74ecd5caf2e633fc4f9cf25fb2ccf5a83f379e910fd31b00d80408fa70d6039b1fc892a39ff4f718a94d47cfe663fa3543b3ad811a44b39097effea22c36f612a3092b4c37164944a5166dbb7b977c8512c5c98a8ae7680aec63f631c583a58dad053bb7e4630ce735d70e4a673d53349945dcbdecf8e2a001247307c26;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b5dae5fc4b5f9114d45b83d5fe0aa72cee9cc660c3804a0cb76a1f60b38a77f6201a00e8c7564c102ffc01e88006ad414110e192098f785def00d2e8609be5922f89975669bb392f984c9adab3322304ee08093f1586d4e824e7761fc6f083468c9999e202c20ce48062e20b832dae8f5853efde3202c559dcab717b84d028c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbaccefa0c1ef4a21bb1386f572026e532750151a938b474d929c1cdf9d8a943f06e3fca0130c8d2cca5ebc72df3096e3b73599ff68ef3747e30f79cb6553a3273ca17b065f39d7489564d8fbc3f5b6d4595ebd6204c33b3e9acae47bba900fedaf36e2ed2eabbd6f6d62350992882052825d272bb66e0c0e794e5328818897ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb35c4c32833f7b11f29fd18b430c06dc7d361afa7d8149181d0d00cfa9bb3a331b37a3ecdece226c039be834ac19f027ff97c1d5a91ec3bb9ee4ce470661811f586cae85933282ff848bae6a1535e5aa47d2cf9734c8966828b933973c9d5f311f6c80eca1793b3ee150d71672e24d24613c21941a7f53a8b93ff5f83bb026a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70219c7537614470805f9e79587f05b22602c980377fa96ad238e7144338b4fe2611375dc7f7773ad9dd7d3953d42655c76152331e5e9c94dc127f9dc8dcbd1c225ed8d863ac32ff02859c72fc76eef3094821909b3204b7710feb8d755a7957eb722513d419ec3f176dfae5faa487fae5155042a54b3648ba6a42df6a52ec08;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2988dd5852aec1e91f098bbabbb96c4547d09350988f52e279bb6e542b236eda98db961edd288b0f8377e94f0665a6937025ae0fdb35ea948ba9822a26fcda3adcd95f0e52f3e10dea5179fdb693a9855240178781dc852b6043ef02bf14377d2a3602371350e22a692d9677c23908d29079b5c7dfd20a4c434b1ce72493a29;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf2ead5f26831742730850a95c74f74a5c84335201a33b65bc04e646a3985dba9c4cddfe60be9bfb9429d0ca8950bf64cdfeb38b8cc0e36416e12ca22f59ff1d6402062a73d273d6c6415f78d469c772313c1ee88aa7aa87f4835351a2c2d49e703e5f884f59941224bfe0592771af9b0039120be5731c69e74df6cc00d94a02;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61c2096a055e70998cae7783bad7331d3df61fb3410942fcf09068c2bf4136777b5f7930f6be40925e4a2ad0d6a7c9cf20816de866d16084a0a89854fde2a8d994154268b9226dd7e6c38c82141a8b2b33b0a9b773a7554cff69b14c8b3f382cb63a504b58857d704532bd804a8d5880fdfdb3fa2c22b26a977d2960d2705197;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76f43988bea5ab6ab150b185b2d7b8514bbd2a8e17a37959b0927caec1e329eff60c586a200c94830faf688481ffa286accd3bbe99f8abc9a55eadda9f718d6600336cb3e9e5cc5bac6681f9956ccdf3e6fd635aa5f040ded7e1254939f355b179c6125c2cdc67a8f7455eb1c414491f20a9121ff374dcdc66efaef0b6982c5c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6d3a6e5a4f0c3e4630d46104399304ac51bd22afd267af74628326948173316fac0cf9101f4ef497cc4a63297ca9f8a7d480cbe61cbabf7ee19847ba6dd6c19a3e473753179e44642d6d29a739572b1032beedb59466ed901cf0f3e7f8f25df5418b704f40d225988f42eef414cd6f6d933c16eddccc47fe887c1cf642eb011;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cf0f22738c731b21634d64d12d813a0e852b5ee12a21d064f371dd8eb5593cb91fd89fb87280297d0eeedde80f5fcf19b752272b52e215a4b32ac39a6a863c28ad7c286a3f47a504318d871ab8b45b6a3beffaef4b52338cd86b7cb8efd3d606d668bf78a653b1ec59d47d7d2ce5dd6adb323464b1c5c3a0c5af2ac9677595d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda817bd716bd5abad812836f341d90c0fb742be709a925673b4d6f4be86017985bcf65653698723be2d908a4acd7e5b29fefbdddf146315d4dca9154b9a62d219ebe90ef2d1d031b0aca8819c056e01cfb37b1552b87964c766ad9d683fba2e0e82ca00705a389a786b9887938b2721f6e205c7616524896b5fa9a12372a2655;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h319cef8e1ac46e513359f92efc7b54d98f89862a902fccff68cefc6bcace48beef7877630dcf697136b066c778f2268919b28807deb26a0d6bcb1f55ce5bc2bd557c677244258cdf2806fdd2500028ae54fafb3330ce988e6822420fabbe9849523ea0cf861ff55fd0c6777ff61f7b3c56d3b8fc8a7fd18e06d0299674b494c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3f967a7b6f612c80c9d8c45c72f937f20f7648452ac2d6954c869b09d27b47ed551bc83578180d7c20ee06eb69ea7e557c2c9cfbe434de32a5929cb5276a50aeafc9ce12ac62a7bf7575e356b8acee78ee5af7d445ebeba38fbfbefa1b997a9807054f749b35c120ce35a79a7aafa7d12a61115cd4526859819fce2a0bb2ed1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bda338e1d61e45851db4bcc74d53ce9ff831ea28556f7803067c25b82d613c027e6820afb55fee444c09f713f3296543ad5b7d5460bf38567b70792e578a1f5655663ad14532e3aa816a6f4e9c0ac7709ee030e08bf54a61c0ca28c9fdd9b0e32e3506ee062a292525612d9678821d58fedb18553ce7e29f06b74c1312b03f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85cbcdaabcea346399ae9c308a9930c6fe1999f26f1fd2b876f398164698daf1897967b2c7401b9914e5c23f5e7db39137cad50fc3892be107e05ce7c4010c13b8f15fa04b218b71238a5cb5e486addf790b7f3cf2711250391d0707f69b02116eb88ddd0f2bfe5fcd45a5a9a72189758ac58df671d46fda63333c8a78a834a2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef53544fcc48d95d06f89458f2baf492f5c0bdedaafa0182976573bd3661b2358c8be0b4991635d74cb645c52e64716ca44218d2e793c7c8c87f0873523c873b5125a573497676865d939dcd2cc413db4d21da4acba76ad3321ce75d727f4733b01ee5a59aa8fbe70c0fd6c1912d72def383110a82fab7e555785d24053bb171;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0946903e7f7360666f35d6948e18051e6f6b0e5463bc15fb18b1fa8539e9caf3711f0e8fbe59bb846d76ff0a37f97596db9e7fcd9f89400fb009ef54f582ef08f79b3da72e75e5b858418c708e292bb462d46d6d0feadb1918605079a8b44ec69e1d0d14f278a9adabe45bc22fd8f379a655db6d26a073541a83fef00b6e45f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha754134f73e4ff476f8cbd696e0c658ffd9ac0d1cbd9c10bb10a0a104ab304d9ff9e6199dcecdd4709b0a5c87add201864c55ec7225b20a74ab773babc45aa2b726bca1a2a72cb06894bd607c01e8f0de26f888ccc4d146c184c85a9c1cc0404210cf005c66d03685212ced115068baa41712dcbbe86886377aa72dc8b85c784;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdca74d0d95b93e0cac58bde116f1fc8239b5244f5b73277de0757d0f202fdaa5584f9321bba69f6d1151179a83c0da8e3cd0ee733f49a1a3f6dc7f814fde821a5205f1ae69b8f372090e8a739c01933f532f00e557461827c220044000eb1f2064a3ac6f9fb2f87d4f4fe70db9976e3a2704af08eb7b93db347337a9e24bed61;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1d8963f601fa802162ac44a85431a386b2840ca3ceb94e785fbbd49361758a657d3a8375d3010f6997f16f6e733ce1259256dc99aa0e86869f20f3fbf50d6cba053351912ef7b29d75a4ef7441cca6eed7bb0cafdc2a33f94507463aa6331e15f126984a53417a8a6e51d7361b369ad8729d1248a26161e3599926e63fb39f4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20f19bb3be0e5adc216212cb2ff4cb715cc32d041bbc1fd6ec856d516435d9a0b7037fcfe45d161d77164ba6505719f5b7b8f7988a4a7a7455a9f909ccd65beeede27d94aa94e2fcb73f219345a61a156066fbd6e37c653222d11490205dc3bb30eee714ca62fbaf70e92ec9c1c097621120778efa6c69201c1c2eaa0be9a4b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2bf49c5441238099aa55c489c8790aa48f7d4e9e89366c2d6ad6e7ab062650358099bbdd8978bd723518e3b81b209748e9787ae8d67bfbb38e72e69ca3fdab98ce22c0997412da725636370a6a4a366f55ab2de1f327bacc77038e9afa9d95627f051ebe59bfa2ef6535fb7dd05b09198d913784e3740e8a0628e9e2914083f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbb5bff547e7539336e0cb4f09f9fb50994a7fdc6605e33d0805bdb3ff003fe9dd8a9e712679edd43e43711d3b9f3d2907da1bed6e2da2c02a2296a2f495e6398d74fab1283056f55721b88b33c5f20f4e8aefb12c88b10d4e450ac315728d991aa66c64251b86ff99da40942c860dfb091e1d9bb876dac26cc2e64eec74df58;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e2919d787bb62d40c904e1d04a6af82e87205e65afc36fd7ca0eeafc2596adebf970261d1a695cf81acfa0dae8491cf6ce069a363aa6051b134acd2d5bd0082ed2a87020a669a7b16d8f11ad74dd3a3406bdec2b3981e75ec4897703ea6b8bdc836ad429c5a1e78d888aac38315b12911e6ccd551ed1215d355c3b6fa1e79d4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7274caa6050a240f38bb62edf26f2a9f2d66fac59c1ea04186233e2045a175bf526e96e3f0102e763bad915d7e766f87139a82227cdf826c336e0f074cf020bf2bbe1852d41470042dc6c99819daf7bf1a75379cf7aceb1ae19e65882c8e369578c8241be98f8530fb512053050d8d0bde226c12f7ef01c80b256e5c73e6f3b5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cefb76f7d5c72339f12a0f15dfbcc8ed42f1f8326640f8cc306e8e01a57fe3f4704c9ea5a40bdbbdaa49051971707f7bbda9f40873fbf798682e00f05d280f02303e626c1d2c7b0edb48009dbed2c4726e5971dc3563936c89aad3ec56418014e285cbd1bff6aa885a7e8f3746a84123d5f73b4f9fc1835654e34603abee9c2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h729d88fcd50e3b62293efa7615080d0733e2fcbb98e6642bd616708028f6420c754d0c05dd8bc80725fc858d5741006778deec747ea41768dd9ab18c78084d73f9db250e9820a172a88e4fdb87643e3aa488bed05a44aeaf6f9f2bf58827fe6165d466f1954b314fc2fad6c127c14a38309118c375c36c08a8b8832390176279;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a2512988e6d573a992c395df972a9fda127f6842ac4e6908c3c211fa98e371aaaf9da738c51d81c612f31f672eba33e072493f7473130dd50a4fcbeea46980aedec15a409764f61b4aaeafe9451681d4d431082c1e9bb045a5fd2b3e7461b297b255430650970e962887d74fd0a873119b7965dbec930a2df0d3097e7f4bc5e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e133859abb927e87dad3a2b353518fd8bd81eb55a44b57ea1fa166978666a8d4cd3425499245e09577c8247dcc42ac7d76acb65075bbd918caa6c729d1c1e8aa763080fd9d759080369a26468e340c97f3c08fa5150c21aec042d6400b3ee6c163af1d3dc31ca78591c2570c10e8d908176dd10679d02bbd88e3a824568a162;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d3ea8ba74efb0380fb554d12654513beed434fa514c2e347255505cb922c440a9c18ff37f181ee66e7f3e7a81261f33f6b2f5d0007929925718e246a266bd62c2907e6f2c02fc799d76eab1614b33204cbc06c07bad0e4208a02437d10d0803274df5398fe91ea4523361a1bb0126bd721b107c045a6a8cf5e7f8515ac39496;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8905b6b994b78107de3baddd553f2127356276a44f04c324610a3926e1fef463b5a81c4303726871228fc8fe19f57351370ac7e2ec1090cad6b538d8bd4a3f85b4b36cab30ad16095c83283a6322bf2f0a51b48c5157fb14fc1254961d439dbf625f6db653924f358829dec3d678796a518c6573a9cebcf41d882b650e8bdef6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa9aafb6f772dcccd9f62f3160eb69bf794d290322b196bc5ffd32dc2f837b47fc2f1e80a80bb8984117e3f06ba7413fea47dfb42499c09a50d834bc9920fa4be33b54604c1af8d7fd3c33dea9aad2cbe571571943dffb84fb0b59f8cf27483cc270cdeb1bc676d182994ef74333d5e90c3a275247550ccda1ea505473afd03;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8c6371feedd20eae295db716c43446c09d5f0d2fdeaaa1d40bcb5e983df27f15330cf0e57cf9e334eace4ac7e98e8691912a257ca7065b950ba255ccf303cf12cdb2c72e98f452a0dc6ec16ccc80be02b922f8b68fe82b8e8a3a58bc9ac4ee9350bc77a2b36974906d09d5bef964f1b7fb7852f889a96fc69a178ecdac6cbf4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95b045a78c3f75bf1a497583665a644970f304480703c916e3810941bbb0af93b3bbcf1c37010d7b9b56b4e8e3f109fd72931dc4a9a9752b231d769c4a545a9798a6108d7a7c1934bdd9b1dfcca85e3af595bc5d5414e85216699ce11710b595b2f2c06d8d60b8ce6376ab665e79d85314288144c90e3747902cd3332458a746;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae553dbad2d424467d6671b4b4be866d76f6a16ee46fa0e44fb47da648696da1e8d20353852c8cd19ef2cb5550b197da391823b3d4b6dafe1c5402528d78ad43e2832d1630069691ffa9a88d86e138eb2653207c095249b0a750eee3152c56895795b308d26e428b794d6cf25468cd44264067926ef3a10881982063ab6bcca7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4a22e6be06e7b7393ace2de42acf18e25aa11551f76dcd17fd104bcb10815861fcc5eb23682cda911f6df2c6bc6a0df1cba1ef4e31d6df4a02bd6cbaa04cec22b37a05bc5fd58302bdae571d16dca2d369b0c01b3b723e8efbeb4703c9fa2dc787322dd579dd2d9acfec3fdbe0466b407c70041c95a3c6351f005e0b3376820;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90e6fa77d3aa6849d2a68bb6d1400367bcc2d29a82583d29566e10682542b5870b4e6010295021e724102eed976363a8b756cdcc4c101b136357faaf15dc7db21e7c6729ea79c58999b964f6da76bbfe55d3271c13d8230787c852af10d03e821e9e635617c7b76728a3002d1b97627e7c1fd2c340fd1e5fc3f62c6d7018e9d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7fe359c9c88c346652731d6733e80735f093e3e368c0ce7e33dd4bcd5b0b9b15619aa9d858c0d3294f8304ed1631f4a369c480745c16e19d33390ef8bb16dfaf30c85a261fa3c3e7f67c61f920ea5e83093aba2d9f86e5674191dc503060505d2a17a3109b66de2a58767f8883a3068b709071a2d2f47a60b396d5d6f5b3899;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heeec0f4a6a43d86ef4ce2d5d80d439b7fcf2193ed3ab5460e83b5fab199e5fe7e502613e7d0fd775d40fc0e13c2387829808ef70e2c98d0c4b826c2ccb1b2468a802b4019edf7899e7d3540c47fdbc4c16ec435a322dd124062113411406edfce609e7d265a4010a8ef353dfc9de8c45a5e441917a7d1fe024d5faab61a87c22;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f041813d38afe273238c936d2e9c6d9b2cc4b9d744d6ab9ad20dae75210691f5361836401b0128a0ca6686a3138010912200180ed362b532f5debe9bac0c6cd38e76753a7ade7b900cea1b648081cdb9112335d9522d446b3ee783f925c2e49ae0ef70297c1f62b3551f438663b67305daeddf3360f52cf56f3f53faf139363;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec12c8f98514299aa38fc97ddae40663b1f4fe896db024c767614059699efdce8c6c7d9f8232cc89327ebf481bf61a67497137d7f2dc5f948c191a140aa1d2acea2776e758803eb89e440b6254bcae9ec9d1b02e354320f2d616bda25915521f49e47326f82e99ee325a9c4d02c3616fa4e55e74a674502486ac2d314a00cf65;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf09d32a1095a1ad5a44749d8adc101b82f3b1e8e93c53a8feb31e0a0ef914e893f065690197ab357571dfb84f6ecd2a9eb50434db413a12b7da4981bb3a053e68c9c40bcf0d77075a5a2b56c7d07c47ced786d1fe217bbe0fe42d3acec9050d7dca8951ebd617b1e89e858bec63b26f89715e36b2423010fc77eadd4cfb04bb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc457efa37cc615376278b4087fbba958f39bc426164ff3b9ee8b3a10a5f024a95e8678eb04168c944b816abdea95d7bd1bbbeb3be525ddb6c0ebf4aaf2d0cabaeca8d3a2c0f59cfa7c48df6394f8cf0669c6726e6e8380c1a597c29d385c798599dbf40a19e94ea0cea05a63ee01ba7d8a2d6fcf0c9c02bbe728147a98a866a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3bc6d04a042f22dcb4caa5e8a71aadee4a830f7d0e2f368a653b57680c708e01c54f458f5018bff96ec1c022daf1ca3c02b1508cd80d2dace80b5a7469a58521409356d1651002eeb08a63f37d6a103bfd970182fa3501432f2dca20cbb12efdc3b8e5f4006362a9f85683be63c5768c2af6ddb3e94360736e8fbc5514f3c0b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39167ef84e51c5163d2f3f5067692b7b51552f3a4635f628ebd7ee6d7cffb16ee124067c7e2b9f5e1ca8f25365cf405fba72fe2f9cb20a7b4933c81ea4a7c345d176eb853c12c02f7561485f3952a457b75edc8c04bba22f963b97f601e0bca56760f56b27073a224f544d5c987e5f72d0023c7c93cf93af0978140a589c2e84;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48bd7106e5a068b2339a8e4636fdb3b21e8a9e2b76ad14de7e28e6952834f43a90f994b5013c452e7b59e2d4e74643658a83ea9cb5e113252fb305a9a36ea2bd6a1e4173651406975cca492c01c7bc29a3850613f02f68e1306407daeb1995ce2573752bc361922cf363c55d59df7fbc02591895366d8ec092bc0aab836ee076;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39f7caa09ccf4d03b28326dc6bd5186ce8251b5115ef78c1163ce0ad07b6995e5ac1b50924eb2a6269328bb60260c63bda0a35016a599bb1b2a469ec80b90ffca9a982706c0004d2faa0d7a0577c63bcd24d656d335fbf796f2f55a863f440999ed97468a73318f551ec1515e51762b0b9ed711bcf0d7a002eeddd8641e71e6f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cd78605e93403bbc4d6aec2523833690b798c440cae05e9517d482c16fe34f53886c1344c4891ce7ef778cd2caa6f3bce95241e27ee839621bc66eea764dad44dcedb0115b15389e9eab21b8e791df443ba4fc17ae5fd14d2d8b7fe3e6e39745300a5572f71227eeac2738ab9b883d80a9e95973e861d7bd83cf924de3d0af1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ad103b8cbb0120251cc9b6557c756d3234b8df16a092e979f80b760c4a1e72da414ce1d3482ae75ee07c2525c261046d8f7f04b5662d98e130eeaafe1f156e7ba08bab05131ca7f3dac0abf90b9fe62cc511d85179f8dd8ebf79e49d2ed7621c99fa1f97a489458ace85ecc55dd49b3a87db728c8a632e7f09d1cd7c0c449ca;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3c24647fdcfd7de775b375224468872c2ab788ba1261ff50066f055d379ebb7ea4a6d6bfe8a32d99ad70ea589b2c1e01c301fc79ec34816678cba254e487aa47bfa6eb1a411d55ae1bab699b46cbb34c23446f797b79447626c4c1b6c1b5c5431c003e3d1bb54f0b50e62edee3cac0e4be3d34f3e0613fed08285b5c30af0c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31d8ddfbda9d68889901dd4cc269268b0168ecaba3c920510872d8c80f3abe686b28d89c4e90ab41032b7a1574b7ccda877dc6e70914017813909e51f57e5baa35d5d542d240785ba532bbfc99766e4eef3c08f593b58598a348f7251af26d1808dc9f573dcb55d1e8df718325f07577b1b4df9981207497d5905f0a027dbd28;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8aac1edb12e965bbc8749112285b4254dcbf07a50667c498cbe2e3254284e3753432b1ef49a4e3352ea4b2bdf95a7ff0534346645af71b67d686dba55e422061d77d933054b317bf89e9a1fc492dd5e7749398e05b1770b1c0d77697efc4e3cd512e1580a5ec549a12a410b62235714d4ddb096945b952ccb5363d8d9f5d83a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heee36e05b34ffa9224bcf660ef06d8e3feca2983c17d773cce6859c3589865526008d5c200738c73e4bf85b5870ffca465464e8a2870fda84eb6320ca7075db66d81089ac82f9db50e2ee21ccbd23597b4ddaf10070999da4ba4ac94862791dc240c7169f8d21990ec6f980e827b21d2e582c92f7f28d2a2273c4aefa48419d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d364f630a93f5ce3e2b4fa37070f6ae662c43f707ec9b9fa45eb21feb7171b470392d7e6990c335f91e9c1a3fe3a8416f84d8e6e109c4627f206ff6c81221536df5e4cd115b86e3420196e11ecb5207df4232b4ef19425d782f8ed527f424d2f5b1cf48787f42bb29a365a9d529852bd40d2ba213b22bb9d6419eacf47127c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40f51f0531b6ad60cece4fdcb2b5469713f9d93551d669cf57f6727ff81c6bc5f247f0571d74d200600acbf615bc5a2e02415f8fdb47ed35388776ad5d4ada7352e5de732fd0ad463a221ac4c2a200640c3807ff8a4d3090f6ae352b15cf2dee9d2c520f6ac97be60477ed5bd6eeaa49f86b996101f78e7f95a2b9abe7ce5588;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73457013efd521eaf56265f915901c9d27e6ed6aebfdaf11f3ddae7fc56a63126606c44e6bc2a8c1a9153edd9b64ad5e11adf467538f8c2546c4b8db21c33c11360f5b6ba09a48705460a34d4a094d08da7f200dbea36c36bdc37683a2b2c037967f1ac881cfe58fedf921b55e05370b223aef775ba08d7a984f42a3b0d3c080;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a913a82b28fbc056530de8ce900fbea48224b2812645bfc9776668b93d4ecd83b92c118d0348a94cf1b40d052ed35149ba3e6e44772120ad4617703d09c2c530e2f6807dc08bf9150fc83fc6a533250f0217f0806dbd561e29cf3bf9e97eaeab5690484cf69ec7e7ffcf4a32716fb5d4be53c21dd7ffc816e4505061d6ee232;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60d1160945127c26464589c20e5a42a54d1bd66e08d6e6116fb6a63457d5713009f32b7ae8684310fa4bed18ec817fe51747e6fc93e420dd5911391def20a8afa910a89d17266599b44f4ebe347f6affb997a169f839358191f9341c2f23ddd3b3810db181eb1c2a9d362fda1940bca657b52cb7cda19d75a3c746a404ed71a0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8d7589348d681a3d7004fcd697c8f7fa5cf633a8e626dea557a18007d21a5bf743a83de8a6abfea9238859700fbde860aca7b1770f6d589c8cc715a96143ce474699f1ca0547d6665ecefee7930ee728fd8d982de2dce573df468d176354bc9ca01e29b1c67ced5937a2bf11a1d1e9a81b80e25faed438a4383f35f77828872;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h814f9ff61c2d04580a8cc4d910ffa5715226bdcd63e3fe59e9eb60d0e33c1d6ec6bb7f6cea73c571909a0ba74b8c5fa08a38c8cdeda978f8405f79efa33104650abcd9517b49e59fa46f3b0e8f4da43f6f6f0baa5b6cb5548d1437b320f97edb337189463693a7e585a587c05fa87abc7afa58efcc2656598be87f4a925f4e36;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1438d15442693cefc9a6d96c054758a71ff467c6c8a1e17cfe3c28ccb60c39029121d2d6a832386924cc12c0de17b7b932eb38d479e06ac2af0bdb949efbfa213cd7035d91d29c75cb3162e421ba5b056f8afbc2196f2181d226b2cb09e08395bb842bd5f6ff73af97e1a62c847ac25f3f98a2f15ac9c8dfc4e814613c5645c5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50c5d72947ab5295b92a43416efbb60e67a4c86bede41a5f691145f01994ef3a74d6e5bcde4562c7d784e4c5bc70a3b25590efea787c8299059a6797666806a7906f46578404bbbb17bf854723cf929a08e31c84c0aec66ade9772e7400b753b1762c37ecd68c4220c10f49aab8773a9de5c83e9c9293b41f42704a259ca2e10;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h997dbbbdb7035e1f0d56e7c59dc3a406ba18b875637d3189a510c06177bd5d3f6853f173047f5680392281a5e3e10e28769e8a9bbfa34e331ce6349a616518529ca2c71816af9997c91a9f9c13fcc077bdebf516b46f057f187c215a3aae925316c3833f53850cc361cd0183718862ecc73c12f361687eb82d7f84648e4181ce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3fb76584f953377b15a0a8b7951257d7b1493b7c822ea3b29b9c2735c8c8f7cfddfb16bae1d1657b046a29e7b6d5fc019b55e4f8a2ef7d8b91bfb0a76e8c78a7af05e9b839475ad18ac374359e86861fd9fc4ada48968300aa525b71474f980a070d0be2051b6de2bf17c741cc049f6c8ba4648e04be881ce2721ea5b837f59;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a5da9c089deef5f15e06bba1929a5e132a2799443bac004fd5c86da422a1f6c2e8678253ea872ce0295e404e81f8763744332cf49915d13ff8f0129ab0356c5ceaa719caa8268223c2b0936d7269ce0eac19c11a218ade91cb584ce92b3d2f716545102d70a30e284212eeb2c903dc2b0225a9543865ad8ae390097a3b3635b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h262c23045a9815dd171458d511198b1fd69d2f97f14df9418868b109ddbfdc91d9050fe82d7cad6966d2e3320feed5fed02afe1571b9abd5c872c9646c9e9280cd3c2032f7aacd023fc5df3b5504dcb2b6e778f46a664f115299acf6c0e71d6ebcb0167193255619ba699827e8c2ba4ad775a596b637331cef99f3d4339db6b4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdac96de3d6a97b235946e286f3f5413ac326daa5ced5bee07fc80b10b90afc7f3d963eaa6afc1cdb99f1eab82fd09232432928872c4750c2c7fd29e7def80850811b8c63d0dc95c30785484fd0399e8f3e1ed65ad2bd68ac2c9bbbb5eaaf9755fb2413cf9b2a8443cf4b555ece07ee8cdf32555e90ddfb401c4bb0f30ff5017;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had1b03a7313d8f8249db20e4b264a369576f1ba77f940bedd555d521d00ed236100838a9d78c6e6b374064afa8da2a76cc91a7c6e19e8bf26d1669c184ed6c7ec1dd8953476ab0e2d46765982c36154ed244a0700241c0182705f6c113ed0acbf59f272d07ae6a1b744acec962dc734de024f48d4e71fecd75304b6ab950e897;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8bd5e0073a6a8d0d6824c3ce9be4386b6afee79f77c41c2e0ccf0f8bbff879234e2a5d535e1905535d3351e2c5e65ad9b0231b0425496b918ba31e8ac85cd077164e7360fc799da097d8adb6dafdfcba07f74e5dfc475992f060dd62f8a0b97bec950d64513537000dc3e21e27c3180b9223e85c25bf676ba9f18477580a8104;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha86167b0662d8e8d92399439a54e1db7d5ce4e6c91b488b0071be21dbed14d80c0ec31dc409ec97a0cde2de4b3e89058b93dc95f8cb365a908ea201932bb244c1dd4ba11c6195142f3cfe5b3759e535878f20d1027f95180ce2857ff9db570fcad42212af1d98385ecb2c432ebc107d4e4c8821c02a5c42f4cfd44311f3e7243;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3b850d721dc57d422000fc36a6936f1c0b852edd34223fdb324374f564566d4b3768a0fe4bdef136666ef84c9a2dbe69a4ca077e66927f39253121437a5b654e6ca412ffaaadaaee6bd3921155b22ee59544e21c7f25e9d1a37846b7e7023351d0348d4387a01f0aa501d72d4f60492ddf57fe184431c89d0adf60bf6ddaeff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4ddcbff96e4f8aa4ae58ab0cc4e8fbbc8008e1d8745028a4c2631a49110ff73a1b2e2b7a4bbc26590e0e7b7d109852c75b2b3242cde0bb7eba242a71462857c465c9e69d99e91dca56ccf96d9b3f496e5253a4b10baad693e677319feb34ca99cc4c604d30ea405f5f1679e7c3d45238254bf85cddea4c766b3740588de142f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45730b78817864301beba304b943fcd693a68523c0165fbd750392cf1777523d2fbea1767635dd79a5643833b3953b19e37f2f3c50443d8201b68d3cf022f8c0abc11b62596490b7d6af8d91a8be688ac0ab3ac10c1eb7eec38b9acfc50bb90357b1ae7ab2fbc70f8b4fa14b7c69ea3558a237a74222621deb8cfe3c13640be5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec01a8a898e8e3d03e85bd817c4d98de6e1387aaac7c0179e47fdfe56f56657766cd0036c1b11cc2664fd2e4c0d86b6a931c5d9ca5ceca7e09611499081164d32a857488ea97805b634aaef9eb6bd7546e3876839ea28d731d250ff0e4849f204990dc1efe62b074e4b9cbfd5d67fada232cdaa9bfe6f6ca068b7b2ddf6b83ae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5b09b1cb6ef24aa77360600cf7d4443962b46ec9078bce4589e2de457b2721b3497394d004bfa96dd08714c310d56d2b6b352c1762c7b5124419d4079298726dac860269015b764718fb6f722a34c8d4e271b9cccbba52d6efa87035a0d34ad036b37fdbbfba118a3a05c22bdd5575c1c48e8c5ae31c97f2cb84228cdd57ecb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e0a7290b6c6277f87a14e77a1e6d98ab8a389f68eb797db02deddf45565d0d11c1f1f43aae72aaeb1fc1f4d9a36135ab1cc4c033178afd6243f045099589bf35d16f12453e05c9d9eb4903b7f858e421147fddc54ef21a5e96c1f8329f349d55359dbfa9d838ba8f15ce1f6cb5f976dae177cb0093fa61de5eb1e7e38217353;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4174fbeaef3130220c639ca7bfd0983991f005171a28bc12f6fcd4971e20169da943b27f0799b02ee67698bcffa4886727aa04a723d4a2a2ee0dd4f1bf0bc2628daf8b59482e3d215c0d95c90e3f3d944582b873db909c7cde710a9c96f2f19b36a9ccd1146adb3b475f59cd66d155152e7bcee7ad4c778df5450e4d53e39f27;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9e263b09f3d6ef69238cf24f5a7000b287e0e5192140b97a5fe87299722ae9b908a5be90741d5ffadec752c0c6ccc7c9a04f3acbed5bfe43a2f59add8520d108584f8c76470c9aa0b3d34afb3ce94264f85a60ea074b4b931352233a8f4993d949fa47d04dec8c6052a1c88389cc579298bda3ab230f174bbe78293e8c1102d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4162ed93d1e0d74dafc6149f00f40d7fe66390729c578f39636296ba954d8021f84482ede639125edb9ec94a3d0056e6eb64e43f7d78dd202fe931dbe7db47e0d7396661767902da86e419695096ea7f8d9a9813206188ffc14a4742b9254471f8554ec7ffac2708033becfecb10a70c5e89eaa4c68afd50e8f00bc2718132a1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90996600d4d02ea3e79d9ca62a4461ac6eea7bee82f19fac0c8ce4d6e1739fdf99cbcc85d4e7e49a4514bc3cbb8e242d685fb27904f1bd638a7a70fb527ef70bab80269c749f4f7e8628638f3664ae9bbca3166ccca7cc6716e290eacef262369dc18cc347e782f2cb9b793ca6104aae3675ecb8299046efb4954b0c1da5c01c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87c3a7a2c823e8042e3accbc278c0f1f37e29d3c7f724765b6666b0316f2e6efb3e3ba3c807942955076fb090cd36e1e23d6a0698acb9c969ff3e82434af2cb2377697b92753b93503a6a00131ba35d801f449d7beafecb1e5b1308e7d1d08be2f584021ae5fba05b5f0656ebfa6470a528d779cf641340e5492f2ab807fa886;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb14bd672dc9bb09148b5f27599cac9e0cca6c8c20da56f968ba41b7e2421c579f7dc3d3d0210d8ca9915a32e5203cd773324f30f25fa5ea8d9e0c917b7b68f24e79d4ed8b46de5712d9c5f556149b025647588212fc257d8c7bdc7ab6b2edb0ce73fa1e6a174187cf22c2c31e1e8fa499b8f25521a337393b60e07ea9adcee48;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb4aa19d862b894c25e752ae29a2cf0fd21d640618059217f9e0879fc05a8ad8737b9ab0af31874b5760c71c04b1c5e70c4b130c98f890594d4c1e2c8bc8591365288f61733b45c8b9ff57cafb6873ab9dc12acddc74f85baa384ed6d07b66acb17a64b455263b8a5eed6e589cf29489187947c3f33133930a8a44ec9656bc8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h423bb5e3d748e3a2f578d30e6839c6f4717fe1b5a09b3528c3bd3cc7c56ce8a9fe467a0b39720297b79c05d6135fc9741b66110f18a63d5ef2f677779d7b97551c98cb495f8879d1e9542dffd2933bfa0fd761ca32b3a583b33a725a696871724463d8b60abe79e8dafe5bd1afdcf7d56f0c43a5095d6d55404cb2731f219e75;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49b73c884051e10451d0e70f24a5375a6d1e2dfc61ec199971ff682ec0f41cefa3975a6f048cb2802c772315b0ad4930ca8e15d6aa4444e5224be8d935fd7f1f9697c5a67cbfb3b6fa7d22931003413fa7c0b2d8d60b872468752bcdc78dd0ef71b472ef2ba76143b3c1e4f78b1fd544dbe833bdecda4382fb9b9895f471e837;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50ca9ad5d6d163bf08d2b61e9adb72aa02a4c5b4de5a14f721275330459304a736a0f02f350f59fe9969b9a2b05a88ba91fa8b9a529f80fe0c89fdeb624883f1cf63e0da017ad77ad73df52db96d4d318dc7f426fc0b7230dc4a709980ed06f85f91108b7f84f5eb04f99494a614bc89c5b4d6c2fcd50e85a0bd9944897910b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e48c5ce424bbf3d653b8ab259325e5a3d4b51884585de1b01c0ed40b210dde321b5c145e8967695c2859e31d0989c4af47982e80fc84d8532e5c6819f529cf95ac8dcb733d395af4ffaba63ef3ca7ce5530d9c49cd99af796ea46cf3278965f9fedfb3d18a11785cdbf0855f9d740e28e30299156c70e1888cc13c340a28a66;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf16ea94f4dc064d76504a28588cb8f60dbf032c8f06d5339956647a2fb22dbeee832a022653e9fb52c8cd79562bf0dc73b24dec4885d9d142e53aae8f8b55d4a91a9701abe23a52a2f1c1c7fab1b8aeaf5ee26208b5f5b7cc7070d586534358b8eeca2e63945c96a2e29c72370d98dc006883bba1b09924a2b52d3da06b4b4cb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f8ca1f187a38e5c334f49d7504207d10369d9cd1e77d159865d0dc6a0b6278fa80fcfa79e2d9748ca021561f5b4938c5fafed4ff0ea1d217ed6770380d7f9f60512160f1518a1a2d703ee9ef2dea7e521a5be9f4eeb5e7abf9918b1cc8444071a617baac6bb79c3ea8ff3c273fab648d8a0449c8903ec65d749f6bc08e9a6c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22491d50b5e5c4490db4527439ff0872955233aa0db20e0bb1265d2d66d3f82816b65b63b6e65517a7bb612b51668008195a444208cfcc3d20f418e58fb9a9fbb3c87c611746de0799acb850c7f2dd4ca039c5dd8bf5043834b4358dd8cac8c06af7b1dc65d5da9f784ff143881580da6f1b3c709cafde9891b84ce4eb4d6340;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5dd3a306973f2d8a97cc8d2bb3844340176783129db83ad4d6ad64de159dde070f5e1eba586d793b9c411116030c6aeff2c8995d717234ff115d467790e6c320ba712fd8aa77522ed2b9f35b8a1e3dba101bdd212228535ad4a03c0758bc4afd3fa656664f26b3e0f96a30e3271593fce8bf86b0acd3886c94f3bf37aa6e9c66;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha231097761659131200f5e82e830bb240596dcf5ab00e7ab45dab86ff6fd62c38762ba0f6f03b965d3a13a95cc8ece89536c0fa143d482ced139c610266536afed34d0a3202840deec97cefe7d508ea85272e5269e368d4bdeee1ae771838eec14deec3e28415ee2a9b93e4bbf175f0a6c9b4703a25a961f23bff98d519aa58b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ec3e19314d9f45f895046a2c1f16f0eb012578959401bcb4521057c4520e61467c5a15b7016fafdd017a111a176b99eb2d483150ac76d4c49a4a597cec47f63317fc631e46295ed07f4e058a4c08416ccbcca745f29a87572194aad1131ab36018023563f0ab66df373086fc6ebfb02843a0957a4a7151984133e491b82af45;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56ece60e8b2d6735bd7c0f73fe803124381ebaf50b9e941cd6ae5fb66326e03f960185f57370ea040b82297c89232883bf67301f7bfecaf04c8e0648d90f66b77b4c4070ea24cd807136325e622c15c4c60272f9b8a69fb47ad778d697fccff6eca214c26540f19db233e7aa4e2eb31172ba19a7b648c9b6b729c422d444665f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f915bb8421c1da87cfde617d9cafc53b556cd872d6d6c707fdaaac3b64bed9fa84ccc91f0884fb3320cf1a5aded109fe32056e3130ad482fbd6190c2927fa6aa68b65d5a0d7b850d6f8f658c0e2fb0986d47230040a26615a36ae2fdab6e6af9ab19ba85c8e17f28653f3164284df701eda48832c7ff8a56bba042afe85d0a7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5672f0b7b71b2fb6fae260cd049df94621fe04c84de10a8754475fd792ef969d186a73472e7aeb74f6a5c3cf80388e9a8e494b2703d55b1cc0bb339cdd9341a35e6b1d61f2ebf58694c334823a4cf25ee126ddca6eb0340670053f39ec75c5e90dcc70499e42cd2698feb57e2ddd677a0cfb07b6d5a5af755b3c0c6e01a999a8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31f2f45f85bd0492c4da1ac634b83d1dc2186e10cf24a6b7058d790bd7819f1a2e1fd81a9829ce1bf66fac2052a5cd5a620f2f217b90a9289fc668643630a81b09e4eb35262ca7a8e608afc35ef18b864edf09cf097bb519b9552e5d231c943f1e4d1d871ca52d306025ad127f2aaf6fdcd53510d68de01273474be30417cff3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6b5c2dfd961587b5a3c8f078cceeafc2224a9d1a652b13c86d4403e51f5e8f6da715a8c04c674db7e5285c859b316908271d4ba4910e5ad1fa606f9bffbbd390a9116b79ff2623b5f6160c32db533c69943e9b6392ca5fbabc94451e7938ed42b7ef61014629f3d2317b20648ce0ccfb13018bb453375b6116f20626abc6b16;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb6469513a6670c0958c354fd2f3f06ee84c13b8ab352a1bedfb197703267c084b5821252a656c6015bb1c09fdf5e797be45b4ff9fd595487602ed997c0fe54257ed526643208c23eaa337a735f7174c567e09709d382912b52fc06330d4bb9f9022e33e70a479e332672f4e4008a236f69fd0519b5a3f57520f9d658aaa15d3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0ab587d8c7ed441fab5909fdea4c14b3d239c030c28c94b120bcd5afe032f1f06dbb364516650025e19fd7dcb6479c0653f6f97fd3b0de93309a56a3ace70f8cb9db37faffa46fb5efff591802ed03b5ccfe76d850ab54a2bd048a3ea5ee78ede9955be1db0e24b35102af9537cbae3b0d8ca525c3597b3e1d3ee64d1f46381;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d2516e357d12508ed6ca2eb806dfa3c1558a2fcfbf3a1db407b0d250ca6bff35a5414019b9e69fbec223441f520f8e329069747027f202f25c6d37a40e253b2875bc226fa39fd0f86dda2b08c893a94da2271e8c62e21938fe1d8df5970934ff7c7143b6f33af22fa5305be7807f0ea782bf607a7739eb32dc82299739701d2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc991bfbcd195ad7a720c972ab939dc51cfe136ebefaded50d275349002a06b21e778ae790b50e50fefd63bccd9115f019ac954453cc9ba465ca3ed1f68b464b970de19528e8432cf43e02d84fd184dcb7f96f2369609ad6796c13176695dadedd29e8c210760fd03e9a1609b60af39abd628b1fc18c805627b86078ada81ecf3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92a8e75dbce38dc61c94953b2c33d343e515cfb1207748dd93f385126ef70b9412c8786951fa7556fb9c1a9532dead63554576d85ca8eeb1c5ecd374894626c15e558c4a909a52d3210ed053bbdea1fbe6c3c6ba8daaf070a68461941abb2ccd84eb9bef6abfd51414153c29c2f888950e676734f9a241571a705b0e531333f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8af13b889256818a097bb207f6cbabd585bb3a15a6419328d7fa1a0e3648c3cd14eaaa4421f736be779916a6ce8b43f29f59b8639948f5c61f455cec3112b9fc09a42111659fa0eeed7ce165a0e9b1c54a1ce40674639fcbaae70825bccd9324137aee7dbce205633189a11cefeddb6555d335d82879686d5fe5698e510617b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf633ab8157e832f3a72790d0e4185a74b5d9cd0f06bd3b65d14c61bc6e1ee7e2a21c3c9d66f0d126b6ab20dffbfac3dfeff6015ab32a2cba17547a52d3ccb1b4e6d98f9a7f6174af93c659c6db5f356eac8fef424f9c1eebf4988de856cc7b627a30d159a2f0252a35427d8667331cd2f3647a668980f3a8aa2e68fbf95b7139;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36d78aaf5d46de850c368470c238e7444d9420725122516a9e64944f62f4622dc07ab55c071e5d1b36013006e6d3d8b6ca07aac399f5202f869836f5b403fa20570d6435f9c72c178ec65a34bb9a04f047aa9a90b143ce170c6dca58b896e1241ab5322d241f9fe260f94bdef9a72e008e2dfeff688645d80123a6f4cb43078;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h255eb6aca1ec1de2bdb9bbb23e8f3ace5b612638a08a4d4b4630f8a135c448e9aa830791e7962ab2a9da27b863ca4e7c766bd597c80d6d0802d16bf7511d1689fd5bb0580153aeb2193119cda54bfbab452deee83c5c49974f1957671438cb44b5f4515c36cc3091f799862f2e793717d506f0f17e9997234135429dd5c8bdfb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93d4b2dc4b73a7d08aa245ef09e024a2c96946baa56faebeb470fafa4c6455141754fd512a3fde06cad1ee3e8af8f25fe29614776f21ce41524c26f66e546ce71140d4251ed92766c77349ae590a565f486fcc27430a23c4365b49ae8b75f914f0c604c40d991bd8141fab43c2db7ddd28701f0a174d8aa0e6f5f96d8b1ceb80;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf19b05a10dc6c35ac864457d69bb6b932b2e39205780b9f713d9dbdcf5f7d593f43672f84814292f56021bbaea298de7e5962fe71537424390894557d7505927af769817fe6559d69220787d399127344e002e97198a2ea48887cceec6035ad45679269db6eb7e1fcc7a13e808e8731fe30fc0f6b69c85a3d7e1b61a050bd728;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha59e133064e0a155f44fc516868be2763d4a60168f3bcc49d17fa8c2cf77909d368512760b65097c9677af21c5e801a036c410c7577c6969d41f666905781939a887934e18d8f616331213715cb1af7eb6277571e80825e1af882e9515cedd5047e9ac4156ebaeb1a671b49121a823e5571e90c359ff8d3fc8578783f8aa3983;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74084c24e0970c841c1dee91d3e78f35ccf7adee890fcd6eb3498d88905cb68770087ae1e1b8ae84ce2dbdf2d75fa4b879d1cffeeaca4d29f42bffae4303bbb34e5f43c6a250b3906a0671e77dee8ae5d0476af4eab174042af98d3b69aa157718808f097f5a38adc96f7c89766280d109b67c6e6ce6bac8a74158a5bfd7a4d4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e49bf81cbf75a6c871fffb099c35b23f88e0832b29da6665dea7c022b295afd38cd27895a88184a36bd54ba52eb61821fc54b25137f7f5e5cf5854a53f484e3fc18f8c25e1692398ad250d68bdbdd783c5ec342bc1cb4ccb1c35e766f1ab6cb1abd1fe0f89e0346781f538d90ebf585173846a590dd2c1524088614f52ed0a7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43fc5fe41fe2850bcee867afdf76286ad65f57a3202a3b7046635f969be932facf9a97096ccf280ada04251f86dca4e279871ee1038b278da8d1ccd966ff0accfe12a2e19b4330f6e5238cb31bcaad52bf234c58e323289399ae4e648a9d80bf0424769e3e81cbb1ee167dd314e2af929a5f8e60b6e99952e113de20d1fd5a1e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d8df443ca58416feddfbb77e1b9728bfc2be4c6095c9158d1fb2ad9261b9d17cae7d4df650f2a844e252f37148ca915605a2b0a95ebee1b580293f6a052876202796d5639146648d668cafddf297af9c1dd142d22e933713bc24c122f9eef588e5c9a3a9ec592a21c1882c8e989baf5d711221dcc1ff2db2ed38377e4265ff7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5930d3cea5ac13aade198108ab4be8d8ae4fa22317b8a7dd02c0de1cd05f905ceb5eea2fa4c966f9362a5fea07f00822f2dde48d4df9f1d0455c884a9ab267cc5f61a859b6a9790a465ef95384632be680908328ec3a263d4272e24413499c2d3b463f02626a8875f6006d325c4da7cee613c4b989f7607cd732ee546859fd2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6609f5d4919b0dcbd34621273a6e0096153721e38ca2910f72a97a2614b699b14a2eda2cf337f47dc81b168d34d52a209b9820d5beb46524cd67209dcab27336653166609dcab7a7bd58288ba57e8744bbbbe579bbd4c89166a46642f75508b62b2f3bc05f3b42ceb7bd6df7b5f2c65fb1118d0074818fe852cfb68d0c9b8934;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bc6dec3d9241165d470a5fc1c4c004388d1114f85d2d1c61f077373b540da1a370e70cad816994a91fca330e7ce4722b9de2e4ec67413b9f1afcf9b5a4484f2f6158ebba0e8a812a5e9132235b6bce30a8a457eb96333b788f421693ab67006ce974ebe445a104690d28b781007d65bf00f6adefc8f73dc99c75867dbba8f84;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6039bcad7232b2c9bd130521e3f50a57f3856cc3965da8009ca88b0d0a2308d1dd6cfe0b1dad7eff2d6af1d783439649843eec501b4671c4cae84177542bf7e49711c6d452be7bc1a7176e3fdec3009fc9809a91063504b3600e720874d18df5bfd08e630d7654cf03ddd01e375af5424351092ba1271c8355cd3bafd7ba5eb2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4350bf3882a57c029bcb556f80e2029b709550035baf1fdd31be725d5c373e053fd7cdb1bf7883191b50550c732f4e07774543e60c4e99089a8d9713e2d0b7263e861f2ed2c7dc9bb664db5c6a976c78765406f7e2a61535a40e86316a6c914ecd7832966a250992be1aed99e06c38ef6c43af9e1bad94eb9f4f39680bf43653;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h776dcdb008d3a6fc1bf07b3aaaff233b545f91636adf278126d01e9e223d65870abf5b134cf5cfc9f38a3036002896dd25d16719b080f5e3839007d6757f1410c3ef210ec16b51bf2235ad094abb0fa8c0f4088ff24cf0f6f607625f18b69b19205dce53aba5492119ec3fcc953e7c54f09084b3487606d16e238d2d9ab1ad07;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd0b87199839df900cae67813caf499f57938cc5b0cf990f32310d2728b374d3e66cd14938f660590d502682fa72a49ecb726464c90d3bb0b9dc52443698c200b27ea4e3f67ab5fe75a4f3821e3b3c94deb618fbc2e3bc1298a6a50be994a4a4be1ade688a19b03d851675daaef437d8a0ed79f48c2b4d275214fd692f133233;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50ff66ea1ca3cbb1c562e634a3537617a16970300d771d10e27bc0003445209b7ac9a491eb86b71f54c3d0abf565679210e3e07c28d34cd44433224bfd35aa01ab64a1a52e4b81073fef88cdd72b4fe279833adbf3bfa9165c39a40c5d726b7da19f06b5dfeefaa988a925eb6defbc7cdbdd6a0717a3348a5c3001a0b46da5d9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d9054712af0cf96b1367f481e4249185d68712afa995fbbae82f2c795e532a7db19fd0c36b72b6d528bf3df9fb30a4ef833632e13254503d5a45f582ddc1870f7cbe2e08bca56b4894a47ff284844456ede1f65cc628db74c899ea5b1657b7c2c1ebaa9c5e433939ddc71e32a8f1f0fc456f7766c357a1d8c14d9bfc49a68f5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h580bb690893c63a147563d4c082a025d520e899e0d019b050048881c2666fc781baae53c12c6a56bb26621793329fca7139e61df90695f34a4849b087d6bac617f7e4075607def890619971baf1be658c4a8190ca9ab9f25a4018dd787f12941237099d8f167689a8101d364aca446a28ee3e050c412e298ca7d4dbf1846acfa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18ff324d09b4d153a301c251a95b84a8839ae2016ccf999dfcdb730f53c069541691cd6464b374908c164f8520e78fc9e2c26574a0e9e62cb36a74a490af15227ba793a16ad7e7b82f9634b1529abdd14c17a6bb6f897cb1f65511d399bd431099ef6a4815dba1b744c226a0ae368d12fc8ec14d6e8d7b4133685adcce463494;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd047b848b4242ed73d706c92b9562bfb4ffd35f172dbbcfb5d34fbfd62bc3f3429187be4ea5efe605f802a15e7289b11e3b0add86456fd47cae2534cd490e04ad218f91643288a17c1d8767e771c7a558f9731daa67745305faed5cda396b59b79da2c18d0919756f7817d833a02b08a6fb71841eb72a65fcd665337085ca2d9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3e2edf8cc0b0b24abae88c1b95178648f09ea87722460e59ab2e489e02b0fb2b7ffe973bda019620d657d54b1c4cff3a6d4ac6cace06ee5e8a64c6d4fdbc7efa5d444f6351b031f2a70d3e91cfb984922ed906aefc2a4230d275745cff9838f73be6bb046a949761f38ad3d406813a489ba192aedf84865476bf035896e40d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8227c55aff3ee18acb32d0f07357ad6909400c205fc1134568711de4a1adf5bacd443dacf2dcb67bf1ee8169d5c303c50b284647f219a671134c3ff4c6238d248ef5d49ea0a8b475e598f3df02514551ca1151234d08ba68cb799535b98077a05ad6977f1f50f81b07016891de2bb0e14b5638fc3a161d68413c2e9eda4c2bf9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bd5e9448768572c2572b777e2a84bd48e4118d36ef42098ee8271600c3c8dcb1e96538303e1ce5738dc498ebf6943e70c68d7d90d855c5451b4505f178a42b9122175eb8864a434f3197d6fc6ee7978bfc37119b3aa43ccf86c5622772b200ffebcb0cdc739258ddc7b325dcdc05e60f6faadc5dfc5c3e45396d5d5bb038435;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61aa167eb35cc05a3feed9820a89dbab00ef964b07c548c005085aa0fc11cc5c78fbedbdbd36129208aacd2bbdaab1c544f94a322bd363768d83bc05125e0230e299a70ef096b746e98670aa8541036fcf6a4faf9a8a5957cf0726bb5acd7da9c6356ce989e7284d0cbe15848903c88ce0a884226e6aa5d94ec34498e7209c5b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h578ef6cc1c20104169810f49a2589e921fea43114f279a61c529ababa0ee0424b0ae0bb1b0eafa4d82232f21108787e9b49cbb23e943718bbe997141c5b69db528b97bb6224d0bded0a63ce624f549c56ac803e5951c45172b64bca1cc0f767ade600181dfdb8792b3b58148b383ab43076a97a475ed385bb8081f343ec15482;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb11464ff6781f8491943817e07a0ace67c1349cc888e479f6462d6a400dcb44ce36fbe449dba04281a1395e729339cbb6b905bee0aaf1f9615a6449a91928cfa5c40914b0470bb842430d51745dbd9a667a461f1e13b19ed80206c3421ac9dae40ce9f7d4128b3f8b06bfbf96d698b4df2e8ce96e3c6d4ca92e041a604b73324;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf73e244109d21edde4d5f0f08dbad9204634007889faf83cebaa02eaf4025bbbc414f2337b84b196020d54fa34b8195b530f11913b4a3eeb2d174622ab9597cc48a8cccc2165a4ecc12a1917b428d93dd71158b49b88144078eca1c5e6f2bc81f67640dce0582dfe5bcb9891df9a5144d23e64bb4dc45f00fba9c502fd3974bd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6e413e812436188ec770065e23f4427f4852f1090072d9a402f8f8df51448e430911ecdfbdd9fbebea87b922bbb5b39ab56817f2a3a82b62a6f307f0bc5b4f00659942c696a3cfdddb35f32641342b9fae33cdec0e1213155217fe03f1905dd6476feb4c22949369fe9d8e71e5b4e38d6ac2955121df0193960b6e1d405a015;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef7380aab20110406438564e123bf009612348127d61026ada13098dd2daa5348acd33f99fc3f8e791d21835af16e2453cce08e56f990a43fb151b2d58b407f7b63a7468d061adfa81ea1ec44b02d146b17428cc622fe71c8125fab2e4b45a79f23270e058445a2b454cacd928723ddc47da9d7251f9f114646ab924a6da4cbc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88d70e3f575e87d6aa443930993deefdeffd303dba73a09a99a1fcddc135dd5a5599f55d1172cf232f595922c8d769dcad41996a2e02f3c5e2fe507d3a54c0dc428981fa493c54e4d0aead5c3fb1ad67aa29022c04d25e49d7b187dfbbb96252ddc3b945cc2868c6c0d78f5cdc50f804d833d42b0b9b771f31cb8e5882754505;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26ee2039b2897a1ce8d1e1e3aaeb837d34413cc991d9f29a28d46ae48dfb31d162f5fac0af39255d350fce79091b9531ffe699fe95ae3d52bd31cf6b0cfb286c1dcf7012446e9756abf15625c529027274d583d096da5f24f2b5bbe48e438b1d0281e6252460be07c654e4a8b80078dc40ff3c988629b0110e1f07c4e0671a4d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbceceed7fd3670be96a95f527d4368620720d036e864e6b81d66a002ee5ee8cbc8a5422242faa1e81e69685a2654b4e25464d4f92060130db336fa4abcd6d4069227c2c8c684832f9383c77863ce1c294f094c3c22e0d16ea3fe7b614f748f97ebaf2634dbedaa34dd1e992a70764a3ef1ed32da33eb997beb44921d4083e596;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d4deb127ca4f7cf9c84480ae52f40cab8a221f94023f92e4472386810689810ba3d17701db4f3949268fe9ba920a8102716ca0ed46ab03eb3b6d36c9f99620e1c05d237cc554f3aca82ac598c84207d30930b826219a06a4dbab53e1751dd26ef63f1648b5a4df11164a95a78c69d34b978153c1bf510a92350475b5becfc19;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he38a9309fe9f636760ad1cc6227833d2716c2040f233a39fed070c4699ac077f4def9c2044baafd51db6362391d2c0eae40f234ed1d104b416319133deec89ebc6734974a11fe8434bee8c5db0f841c0813812c71b4da81b6409ae6cf9b81d9fad164eaa521e4c5239be78422da118e4781afcc59ac5b6bba8128efb9cacf8fb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9649e0a5e36b4e7756efb638c9662113e530e50725d01f10f1eebe398ec0f8260ceea700c74f15404dbbeea47acd2e896b8b3bd93ea91abcc229b8bf68b19c1a3c176ae7467cab415ef3ddb9ecbade30b75f2cb7527d21be6b71a2b68c3c7705abad6c2608fd638462bf34e0798b5297f70440624d133d35a01161c97b492451;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d68e61a7bcfd2cad43423fe726d46ddc83032edc9af53a1e32976f9478491f3a589e03e143f8ea9acccfdb1e8b8a0f024540b3a76e5dc5f99f56ee985139df591af2e25966ad0bd7e301a8e79408aee5c1cea74afad79a5a233618fd0300145ab282bd82bf06214c8868c23baa5d2b5ad99451855c5026b7a34df961ec63e91;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bcabe9c7f2e2152032bb75fb5865e1e1c25af79a7285973dc96210461d7b2d1fd07b6b0ecd750f0732657c2f93dda44db91bec41ef20954ae2e9574d213e68dafc0dce23e902eee6e694cdc144935f0530827d31ec966765ef9bc55505c739b575e2b463b5edf6ec8c77d6d8ef8586a8883ff4493e937b56c3f1df860319a61;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h927415a496f7cf03a9b6e05a8aea430ca06976166f66bc450cec99b9f7fb18a8dde220ac9b702209fa4196353dc7bf0ddbee6d0976e83bac8e2a5d31112945dc27c68bd8273484e1716b18a822550df1b0b16897fc77ee20f8cd3d48697523efe51201ae8fc70254797cdcc6bf92ac18f64c74a3dfaaf6be46d153d13dcfd7c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he83da24ed29412e57aeefe9459bfcab038ffcdf628c0baad5b7eb21725761a23a9073734088e69e7d8889abbab03373ffc3d5a1e60da4a2bb445e7dfe259fe1666cbbdd1048db6c0ec3145b74305f93eff9edf4c4d980fef5f11b508a6e03a5f967c6db665db65f46e90c07a1d5bb5f0bf85e2e3f90bd3db36b1ce303cf8a69a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5bc877d576235f2f9b6703c2f8633dc63fa071616695a1e530388e09e834b876bcdb95c77e740008844e58259f4cb791c5f07db8dc988c78878a53268552f7373953f394dbab86350baf6523110b4e6158f7f5dbd0bca566a59b47356175abd7e52be37fbbb10f2387754fc9636fea4312b37a0590833c0f59ea606e5e87b65;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12274c5af01a4d326edd6085f6ead55501d967b0bf876a5d36b36de3c5227a6f68c952aeda98373d6b9442377c6b36e99810380400e141891bb37b416a9c80b88bec546a30e890119d872a92e20fe99ee7410e77d3e8d0a7554b69f510402c6e280eab90be74ed5d034244a2c5dbc3bc63325ca5b25dde4cf31e0dbd611a8945;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c96d770b37da0fc98a894669d5640c9606728092ae6adf418be934dea5872e93909d6afca13fd421b5ad5ee2ba5613a0b04016317be6706c8c8029e6273fdcca0b542fa12e3fc7587f4b58f895a6c7d1ab9239cf2c2f302743b9f898a1a734ca09e5386df680391dab472fe430c2cc1bcbb0ad31936acf277233c59f2409fae;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14410662c6de02884807d403b06d132bfb6ef95324891f49d4fd0a45960e4100ed2b02694bf1903b2f3bef694d928541744a2b538a4c60c86d83cdd723d660d238963931b9f8a0c43d909b931ea9532e0c986a8fee1e1a0ac9c22e8869a7fc7b3bf134a281c636fcf0918436c60e3378b7e93e4f7ae1f52c75cefee6c83eaeb6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97c6fed5a59da74b10af66bb5efa6de4497cbe35912145ba762f6d9f6f9ac2c1d0b72e39a89404e42feaf3cf97bc858ff9feaa4bb05b817c8eac6f66371962646d9787ef2bbbb81f29de71b189196df10a47d0bd34fbb2a1fe37b65da82fb8917281fe4fe51bfd1f37ba36cfea67a5922a51fa673da2ec88f79dc6da88f0d44c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb49b4c0e00860632656ae11511982cf9630f798a22d491b7ed39c8be8c8377139a28a328a13d5c229554e68e7250257d865d1df3ed848a9cc1f421a5b8892737c8a6eed116424997db4bb5f33eece97b77edef665cd0cc3133d8744c93f9bee5803cc4c83ad95a1ec83c3403f5a79f9b969355664d7c26ffc88d1a02aafd0dcf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h432acedeeb499a463004710dc4bb2dab09d6053db92ef589e95eba475160773d3205e2861e472a8e9b73cd348a80c91a8e35eaba17d356030979cfa3cbb72619893c6f38c9ba6e17dbae5715e887c9819358e446ef54f81edee66543a67d9260229369456e40b8c9dffc45fa1d85bda0b33d47bc8bd1246933338f337b5690e1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d7fec5e401f48d344514f6bdecb16af09bee22b94b773736c4980fe3c500525326db7a7688a960b528ea0ddff65774313e615479c10b80bf4dfde55553f57562342531cec32bb6dd3f0183ab61942565a8dd2640ee0ac6244650469e3a364a9c799a5c53ad552faae3afdd4e6feebcd269221316188e077ca76d693789d6107;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3f87a9b0e477a37a70de6286fbc636d60e0b7c0cdbeb0d550933e6fe16a1f5b195b043ac807653dce9cfb3b9a3dedca16f36142919ec8c559c933552165b84e1678159aa9fd44d7bbd084ed617f67ff6ccceeed259d61495b97d3da99a56725d76b496b286d305ab80d5aae4874a59794f2e326f7cef571a18fa307f6ac4b17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24f12d798eb6d378db6ac7280ab3de94c8b7af6528c40f02d4f494a54c0f157a3b770b794526000c421e81131a62d3dd203c7e57c7d1017b9f89637ce3a90775fbd00111da648b2ab80a3e74dfadfdbe2f3b3dc7a744e6e79dbac29bc4a6ab9f04fa8b3610a10460f7d67060127f1bfeb09711ffab4135f0933b3aadf5d36f55;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h146dc5ead33d94fc527f96b7ecf29f9c3dd833652456c914279e4de70ab6258d0f89ec23f9dab52eed1d6dbbe31a7ba22fa4d3c08f532d3cb8613b68af8202fcd6a4f82e3e34bf42541b4879904cf53ddf81f9db019a562ee5000963574e62fc98194d6e16deaf4093839885ba508abe8d3e5c38325101279c388b2e469bf640;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5aa1b2356ca200facb97662a7c34e64264fe2f52af076de9f098e565cf4f52c0d0114995b06d76b6b35fe8a24db53419c9687dffb9db6ed1ccba88922861379cacd12b7dd5e7adb220cc1bb21904c117b58226136b77ebea21fc0e92ea73727cc346ab372c4b2956165f348da335a704f1b96d376d15b83a4a6b0bda3f5bc38d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c055255a0b277c04c76acf7de2289a35f4f7c0b69b57393bff339d00f9d592151fb4a237c9f315f217a2d1d59f15297620b812e3703be1bf12aee79e7ef72aa52d767edcc2934d821440bfad6dfe1e091176feaaaccb65bf742c0be0b7dc7f949efea728462e4226f6471c43fa456b2dfb6dc3a286f77c1e9bba9b456d7e8f0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha49a70d539b50dd7ffc80acc5e6e0c0289cae4fd1c7d796a709d51dfb219a033c0ea49a8748b41772425b3609ef390755b3f45c4cdf06c58122e4d970edae61e9edf419af1e32af29428d40c77c0eb7ec27a56761f9e0959d93f9fdb8f93df4fdc383053a5a2d7334b096e0fd7cf959301f8a8528904063084bb2c9b275a8b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h366a90d68b00f5193ef485d4e7077691a29745d6d294793644d942091a42934ffbd6a16556c87625b67139a3ec8fb74da031aa4786f84ea3990c13ab82b496557aaaee40b1c772b49aa3aef1b77fa3e16b96c44fc2ee3d61187ad8e63b5d0fa0be644048296e0cb2d9c793ca52438643ab7abcd1c38a6aee1bafe75c341283;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7531585b4ce64b2ffb311f45f12f8c2d5269d8f3601a3403359fb4692bae5c0fff8a3e802b526693f09f57e50f94552e1502cf8b1531c18641bfd630715aed23114ae55e500db4581065d58fb0e0270f2a32d8139ac3e266ebdea30aff31cfa769bf80c42abff34ca9531e43f531f152c998a388b6a5bad87b3d256b3113317;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5e12672c5ef1ef1ce3ad43aea5250c5b5f1ad7385d821fbf0f328f2159fd585952a5d927d6c40435012704d0f616798425230468e92ab60d39a7480c3435f94daadeb5dd114fad7fa4067431e87e574cdc0ddfc94b678debe57a53e8060d81c8a871c8ddfcd5ccb6079ae1b962f55efb9575d04fdfd1e1e26104d4edf6bc21f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6489391f50ee414f8fd21efe6ba02416cc83e6feef3afbd3c0b8682b9d864f6557562015268fb50f2dd84ee4c7a339cfce922038af3ddceaa41a09ef4eeaadab7eddb42e0c0dcbde9932b9076f7be79b2fa3ef237ce2da1ac13726f3d6eb32ed3ccbe5e47eaf060a54876242904ac0ac9347800ec83d6be5d026c76e6c05727a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51ccea13400ed9022a615d185453281855d951ae9e66f772694373fecde229b08240e974a48f394c55f98351271334bbdbe13a70364a450256aba8a902ba04460e56726699203843451b895b0399fff46481329fe73676f19712aa778524de1250bcf6a5a215eeec4914e02b01a8a90ce9b8e85c2e1daeb7067c7d73fb478ee0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e47bb78e0eb350bd6870373f50b7c576bd9cbdc65b5d09450f876acbe54395d741ecc38280d904c9471943e004c16a317ca59eba0d21a741be3f6d2305365bad657b8434c660501106f18bb200baca6a30aea5c3ab44b9e78d804dac5369ea82fd7f06b81515a91691194ccbcb79c8ad98586a5df459c5d5e6e1ff7d3554e28;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa84aa5f8f34fc27945dc5ac65b91b1dfe1420fdc4b81ebe0a718f5415e673e9db00487aaf4cd34a1c68b6315bbab5cc7a912b03abf2937a765b38913c54ffb75cc6b81cca97e4b0c3278bfc4a8c802c3b0f0f7ea25fac188709dc14ea0ddacf89ebc399a1bc1d4219eed6c674a3148a7c8c9317217e1b4e72461982584d5d32;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf473aeefa98f525dd51603048d252271fadaafc963b89966f22c3af68a9888d4d1b4891d33564a31e442c018e8a2ff5523ff4bee53a9ce9831a5230176aefd874290507b10577117eb733ecfd213fd3b50fd371fa871d6c7eb93edcb282737d852d8480a3f3fe1ba413b3fa084bd19b851776399a2cc4531afa33cd1c6b24bf3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b2e91e51c71d8ecd2494ca8d37dbf1f8f3c2a83089b7ec208d223631749417cf7a607b778b99e7340e76a3c735d2f43c917756ce6cc94b3e9e43cdc0abf723a0c6254d09cb9ba36b8b90d360d33399a4f434a03415e912d4bf05ec83fbb07f5100d2b1561b7e66b0178f378978d70e3fa4aecb9b30f7dd958fd862e2c9d6045;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3254135bda436095e0b8153dbe9dca3c8a4bf0d1cc1ead69c1d08d8989d631138972580b08851905a0ba9065b11512d558012fc30d362f0de3cefc2ffaaf68430e74e5c8e4186e28ca53d3bb517e7440f44f64fefb2ce66353342b15934baabdbd36c7aa9ea52126805b7c570c02ea0ef52209ad6922522d381da2f1077ea10;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8fe0015d7cce270d3c82e92627acacbbe7bf5e0654f44be1e012422f0cc4065b22ddf4748b242395b25a4177f206c2b06bf50ca3255a8541f71231921cb8ad68c5c2f43def8b84bbafc93479067777828ad0217e211ae59e7329ddea2fb5e63b9784b8edb24e92df03b4b348daee6ad82d5c0356a88fa90b466e0b030097ee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90455644794072ce2457c5b6dbe0081dd04d6703f30725bf27a8a3c1c5a3afc84a22e7d04308214e00b88846510d4e06d0ccd43996cd02ad9316473fd0dbdd26f9260f9c91e172dd7d134783b8f8358dc9c3b08204f4d4fa9ac5605f4ae8001420e5d10cee3d91c5202a9e3a702c36a82deb5452d706d4732d6a1c44b920baaa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4309834cd95bea0ce7e9df18fbdd9895d2a150b3c6124915c156798daa1f70fda95711273213980daa3fa43a47d2d3595a582d637f00476b897bcdd641e93ee0f788f9046a1b11dc60d404303b4ff189bde23abfe9bbe9b3337d02168315dae3acd55d2379358c6c7c9eecc999a66e9aadfd880a56ba45129ef3095458bf49cd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3435d40f5aaffd24f1f226a40e3ed3fce6c026752d58b7ce8460b2a5f14d24929ed1b33c1ba42c2935c6b86b1c968601ba110327f7506fb01dd36516169ffae5cf7d0b6ae614f54c8bbef3958f6371d555496746b0ac1f88eff11ec6e60da45d8d53e9f1efdcba67a943bfef52412e9e549b44db9057075cf5155fd720c0a5f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h265ca03572d4b993bd11a4efa62a73995527d9d27bec02701b9df5ec90a48b2b5a8b208330a488051c7578042e3f27d3151e32db445d97c452f61b5aa2419e2e78996364773ec95ba4a593107ef430caffe9acab621bf9e5c58eed1271669581d7d837489a17d58ffd084b4ad39854a8cf1eee99080970b3d58981b7b8ddc1bf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83fcf908a4ac73869e43167e9483810bbd4c102248a423e1e2e373b1655708f69702764114ea8e1a93eea048757c836a1f6f3587ad70ed0ab7df3dcc0e9437c856b70e448fb60d0aec3379271a9a9bb9cb09f17597cbdcc190ff5faf992806c1cfac1b0a5c3545733d088d36436ccd3288515d4daa6a5d8eb541ddea07b2af66;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72660754991017cbce479f4065070ef5497fc8acf9aadf152adde72fc481b50edcad13eb32dba3f4f2c0918bbc1d59938f9b819d3d9082f455d0f66f9723bf73395a0bcbfb65a86652a4be49072393b3835c8ab06687250d1d569b400901fb783a14cb525ad660302af18d5b3c69478dbd30cfc530e1abbfc6934e1b248be87d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed2819f2bede39f590768b9ce233792352b6cb729e1f18551b7826b168654ed2d345328b17f6eaa8e41527f673d20279a8e54b62c570347dfe1328221f12d07d6461c986024b3c650056badd38bcdada6714089b06f18b660f0022ff2a9805e20f9d2ec35ced10ee9a55edac2dd381ac807c18fab43ed68ca9f842ab94608885;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5cff790e83f46646ff175e708f456e76f099633ede4e0ffff04465f3d2178607fde7ac5b3afb0b2e770a97da7c77d14f107e2632cc32043f7702320dc471e3944fecf1f65110394ab94268ca36e24762380e18acd87f4f077faa95edf55ed0e84c100ab843007d8582b8cdf608c49bb86e4b5e985fe893251215fd6d65f2830;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c097d42f99a8ec0b5e11af471c7a2dfb6e6d205efafc20ce0d2974ecda5d4c73bab0d168fb2a33edaab7bcf970f61c33745dd051a675b60d5edd8440f9c54eddd80b1eb09c9ea747193d046c8db26a59941e28bd56d1163237fd543015bc1b0b6cf97621ac139d55d522a26d1b04cd8f84617f64c9f0fca1adfbc9b8290f184;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5015a17c75936d55ec6f2de84167ea4ce855e34ba45cfb32d5d1a50a4f15101e74b64a21fb36fa670afb6a1e78eb34e7236c151a512b5051e733a63558988cb94af0a4bee997558e7cec57a3fc862aec67a2bf1e53682b7c7431aed78062ac8bbba1c3c80f9ef607bee500075f514d5bbef7c268d59d185fe960e8da05366dd7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83289fba1b5737a1308e15bcf19b0225064007ad398850fb3678ce9acf4e560c9f12fb1bdef5d0066105a2f7effe789f711d9ab45c84456946aef8dc61a9b6b093a72166066853672e1a2bc59e62f2214b573647c533890503796cbea97f68962a60193d5c281b9c4306221f50d3d625b15eddff6234cdd5e49efad4382c11e3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cf0cbc66983da71802d265a56a5dae86ce049b13067b6f42b088a48e4276be19aac939bc13fefbf24a20d630a6292e0ef7b7040558525b715991cba134acc552986718f217f206a60889eea199c9fc70dc890f8c34f5d5820796c9dde7c7a2b8bb5367e0e332a77a4f90769fd50c558c80b470a8adb148e0892dfe9be6fb6db;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6597430e81c069a61c9a809bacf32a9cd80c420919dd4305fe905a1a149d8db9a833cc0c7d5c91b04bc44958880d04c1ae89896d737990eba1a2af5aa54641f31a5efa76eb0e0aecbe5f2e77c4c621385cbb4b5bca59986ce78b782e1ff9ab8f0a4c177061d0717110d3d60cf77b1114ef7a14d97a9bba219b30393cacc7080a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb1310bea27d82583823149602c31a1a748dafdb3655e5b17141db357062ac07eb5e8677e634740c5f2ef3e83e09dad6a2df72566ad51b0095c4cb701ecc5eaec95f45321eda86be4603c9a35a2902efaacceafd2b86e66cef5ef80495eabd6e3e3080aaa884e1d3649a071476d871c26a268e35bb59cc331b6c9a41dff112a3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9fb11eda6028e1df9375332d2e4939dce0b7cbb007b7c968380735278a953aecac66f02e0bc7853cda383fe8996be092dc589557cb883c55ae78c0344d80225918ca06ac1b404616178262a921428e5a832e706e1a679205ef3eec41ecde624b137ca954108c3b7285f86ece5a22100e997caa0826df2d8b4fe6ea67d8c0b36;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7ac759c40766933019348cc5eeea6c6e36e0fd9d1c5fe4b0a05caa7e2ec243cbecfe9063286fbb13f3338b2787c351addb0c95461d87d607b22ed52d372fc6da9f7d7a2d43ee8b597817d0c80c38bc3080f72de036537fc47d4c0573bf379e5fae09b673fd35f3edef976023adde3622f3090bcd14ca495880cc0a291ff65fd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75f7b8d2e84d81df02ce75ca9b2c9259183e6d5fee3a8307b24a4a5857dd3bcb882be0b1f120c49715fc704c394993948102afc08683a2d77b60dea1181397d5892cd9e391230b9faa91094b9882b8bdf230c09000a1ebfda1117538af74109b1b62f6b652c5fb5bebcd77be0805bef5032fcc51d19fe9ddc072be1ea9df3009;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e3f198435356ffe5db310b71dc28498398378bc559ce6a79d8effd53d6a26638ce4607887f211eea3b6a80d114b7fdaacafe0a24cb3d98ca0af231cd1b5aa3a5c79754bc30313bdd048cf5efd0c728acac0d7125bba8430fd438a03e8db0ee705867895057e5a848bdd5f2755cbe8b3c86f8a1620c12c89653c4807b99be399;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha61a4a2eac3e7b607474a9b5d3e2936a0086e8dc8bfe4a0cdfae9ba5d5b5fe9ae2a6777b19c168887ad2f7ca0cf937cbe1cabef605e35a74f53d802e21375a3754e1467de02eb95027e802f15f5765ab54ff2f0ebdd86f65762334f0cdf1cf7fc456d72cc118c3910cf8a40befae6a72d4f00690e0845996ccbfdf5d9679af1b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f1d4bcaa6805b007f8b83c9debcb293d2ce8c265da3fdf64b2f2344c529e874be943f8d79bf978bf444499dc8125e178b4509f5187848274ca914da6548d8f75b7d73c2bebd387a3e3364266239982cc890b4f0ae67da1a4a4b29340372f4ad59913d33aa00f30d13631d7046bc3aaff17784f95d28890ea9d15185f26a9a17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17ba499d098d9453bf64724cf790e593214def40b77f7bf3f2f7ac5c6215f1f5b37c32e2dd608c79860049f01a07dd2bf17230d1fecca86a707a72decd847387b5b677e3a402b96773369d6b428cef470021e112d4e0d203d1ea242daed150d7a5174f7c92e30cdc50e440b9a280a50e54a49bac69050fe08fc73bef1d410ced;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7aac536c9f772fd418d55de59bbd123433d1e85207a3eb6159278a5f57aa47e032fde92cfec307cfc9308835cf2c68dea6b6b4638d643b3bf81dd7d6d273400d682f39e40e9dc84091bebd95113f8a134930c5f7a014d60c7d877a7a727142ecfb202ca1207f73f4fa89a48eec67f545bd0be063b05136087a30e5ace08994a5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8ca37544fef8bde3c32b46395e127c837fcc36586d65ece409d5925ae090fc0edb2bcd0f2c7f540687910ffa0d869d6f841220874b0684459023809d5f799ac15852ecb28eb1c7f21bff72ec73882557708b0e0f5b36b50177b9a3c82384f288a623fa3e3a7072c2c0042d96150372ce67f018c15886d4f409c0a28011be447;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9205d8340e4a948ac8d4f39ec76c2e9c4a29511b182b16d5af7c06ccc33a70f398bc95af337906968bd4b2fae1d27c2439cb5830accb88db696251555e7aa6e1739b2dd556862b09c8c0e2d1b25631ba639779310b52a82cddec6c8d5249cc538a6589d6b240133999873210765f3060a94b8de1e55d2be32e9ea961b1f460f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19d04184f58976fb0dbe0452d4c581407379ef657c4563520d321e3fc2019b55ecd1692ae0d2cc5a3579a78228106b9c10b7d130faad4b2232f58bb075c5e04bfce70c8b06cf9db873057c49c4c77cd02722a4fbd51e07ad13e7ceb5f0c75eeb8749a6246bceedc3c283f228560e928f8ce1e06110bb9cc5f2498e882c62d4c8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h807dfb4413f26a804c4cdb00979fce1855e6db554fa5c27ff95a72792e7427967b401d40a6b598a04c4f730f056e277d1f04ade915284a21c56fd733c7044a7b2387b29b157593fae6a9f95bd1c7f624ae666bff4f0a2d54e30f9e1bfc004ede706f814f57b241074e558507a35cc7f08cd3e904aaed0a16df575aa1b7a5abd4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d2561f7180f37a3ed4e52884cec0e0ddd6b0e709cd74d0420fbdbf8ab48d1cf3de5378ad7b77e010f53ab8669196b471bbf0ecb4ab9e12c1fe027fc27e109341692d8d8cffd036ba60525f8b076b6c4ecc3d95237ef9e1841c59fdd0b19107ece25d49789e3407fbdf49329237358b424ad239a4ccfb38836118a480907a375;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd9320e4919f77c5a441718f5dc016604912f112b2a551661aaf10e56f5bd56b7be106b6a68b9c16cc54772ab429d47be23eacded166c6c8f12b447556d34b82b1e8eb5c2aae5c136e3ab5cedfa03d42d3405b21331c9a0987b5b8ef4cc40715aa47109d0e1d29e128dee27d8621838c12290d62e9f50dace5d152e952068ad2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had224b18f14e37f1c15dac826554d2f0e184c60f7543c80d5560fc9e390f39318982cb9793bbf5e78ec11370528cfc7586d6bfab6f1ef66e4456a985336d74cd85b498c77fd2ab7978309c718e4e515e114ec4e768fc98fa24126061d02f06063da331e197598dcef4b92713f01e1890cff02ebca641e0a0fcc2223b25147f9c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a104afb652dd68a7e515a2644b6f57ccd364f0a99edd0c302cb02e3284346dd20a9a6497b6603b7ea97ec1a94e3a3d40bd3cd107aaab5df27da5cd505d0f520a3a527cba14c11348ee8d19730d5c0434faac2516f9a8fc8d2d0c4d7733380e793a77286b0f3a08237edbfbc47ac136b7abdb3a45719faf306a6b7bd84605e27;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65d2a6abdb64bd9d879ebd7e899ebb311c5d86aab099f11944f134a5269122adc98d95df9106d4a4026bf7ecf4450c51a327fc7cda73267cd721c70c6085e674de3b9f7e3340a5946aecdfc500ffa96c0b75008f5d4676e8c9234c3f9fa72c70a9cbcb6a0a7a8612f0ef392cdb6ea32844c9d9f275b891103cbe5329f9a2cf0e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19b88bec24695dd86c8a24e573a3f62ae465e70a8df6190df443ce2fbe9d1f451c4cd0416797c09b48b33a1cb6355ec80fd0020b5c66f525efd905c94df622f38f34e79b62a3e3426c2f6670694b810438da6b143c907536d572473fa0bcf779cab9695bc234ef7df27d2eaaa0ba81c3f2ceb9cf7e1fe244f9ff0212aedc10d1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha18818ae2122a2b5ad57d882b655468d51ed5607f01a041d943115e30c8731c662af863b66eab0c6dbe4c8f8a095c68842fff71de097199265fcbc671feacbaa146a663cb15d8a13a625e9ab519610e0fb45e441f42951821d98805582641eab51a154d5bae83ee0d6b890b3120823c043a5e6d68be7c722ab11bb692c8b3c7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9622c573af1db14c78804bd5375c7f87d3a24a0fe6db54d572b4005fce2397ef606d359ce218eb8901da3a6210e9ebe17d68f7374c1a7566655f586f3a14f882f6212e762bb0698c08e3e72219bea70813944ed8f4e471fecbc6cc29e8fb2a63f7eacf38c238eec347d69783d236583f3fbbe61a0bbddf75897a543d03d1fee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62973eb45e4df813d3bb36106be96dd24d5e1be9f7fad984a4ab33ad2dec04d6a8a8d597fc06ecd7475eeced952d8dbf43a3c783a1e4a55940e5abcd6c037ddeb2a4b48d90a110f9509660b086f11a145032cfe755bd04f58929bda7aa2b78ab7334e09c02b4506a757a6102456575737b4cd6f2d0e3d69d69c091a370ad66b9;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1156e3773520c1ab4b21524729742abd464424e9b30ff92fd38ba95cc52963d2ae1487b2d0daee001ca3884faeead5c14b30e5047d1da84ca8c0e10dd501557b1b020b23e8ed1692e3aa39b67046c34fcd4a7ae2fcf1092259f21c5d6d024d90806e0fdce4667f34b5e3a254c9736007c47d5baaded51b8c15ecc9a55506b6dc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h337030bea10870db37989d7895d98c327356adde75d15daeeeddadff95d85e75b619d7be8d40234ef5dd54ef9fa7fd157ff75508f6d8865b6adc3d58d90fc5fe4becb82557d65f888f8b8c0221489b474d2628450dc72a8e6207f79390e992b96444178b03d8d54a8a5d09bc2d48025f4411d6f73fe689f361e06ee8af8b520d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdefeb7af6284c3acad7fff07a684362a96aa7af0e60ca952fe128d965a86ae2a0a6cfe2e8f336ec4789c6494b34782818dfbcec68a438608f032c19fe96debb0aa3e5d70ebe93d2f853adf527f9562c8b9bd3013f206e62bc8f459e186d16005e9b0ddb2892c9993212d8396793b9898f7e806f937660ac450d46b06c03984ab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe1160c8863b73caa28e95f93ae7b96b4967287e58337bbce929d43fd3c4cb46a614a1952d691e623247897485a9e015298f18c948cbf28f114d2b920c0fd415055ac15f544b44a972775d8fa440e3fb54ea3850ac44bb688f3484ab0c9a1c5f9a130f7dcea6d20e8d363952049ef92dc19ad9075ba96b028e3ee7b698c95b72;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4048686d233edd16e245c515abdb102b12bb2d389601c84ef0414a0464e24d6e1c54b8af0c19e7531d2dee05b1858e08b42529fe7854badc8ed1ee288adf3b5b283fe0688dea55e0321629d00a5593fc93d03c1b01fb11c3ca6680a5a1b8f642f97e88d40d526cfc3c000be7759e10840231eab27c4bf04d531eb0fbb793a690;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14f9a7f165f72f69192684e7a5d5ea11bfd80218385e837ed8f7fa9aa081cc29f90e391e63082be4bd5a80b9e57681d6398e1e2fbc76abfc74c0069510cd56b1875ebd073f06aa1bf5c8c4d79041f8ad7fab9d9688cba6d95cc333f3d2ecf4a8163bfa7825915b696429c6165348a026d8b18dc3208d66723ff59b424f1c83e4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58f756176ddc742d2201d1fa3dcf39e78370cdd164b9c16f21f7d7b7f9cbd2f014f068939f24717ae040a66b7a73b9c00e50c434ddc08c7487fcddea5d5ff4c55d36079f5c94105e7fcec9e5f56c970a6789fc79846e08108236cba73a58a4e8e92b331a9079bbd5eea4b373ebe878ef83a06eeae2ca1dd938496675f797acce;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d8e555a272c72c617c3f7bb85ce250ad9dc9b844792a247cc8deeb05d6c63218e6fcf53340b5feeb3614958cfe047b0dd54df8bc242ed7f23c55408bd673797f2389e10ee925dc5706ee178b33eba6540ab2d9933826c780f714a8475985ea153b68ed95d37f9e2c7f6500dc4e87c5bb3a856f566d1d5cdcbab57cd8cbcf3f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca85243ecd2028d59fdf2054d152142b701a2ade1f19b8fa310a71844dfdfa3f24211bb256426603195caecef70fd944bef8ad8e2e59968c489ddf2cd9eeb76f25ddc622e7732404eee87994fa409d617670061bf2f5da2704c996a8181ca82aefe77e87be2bb86c7656e9d26cee239d6b4e50f45c89837f16a0e38babefd18f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45c704486a06fc012e39df9e7e6bba0519fb90b1d2e5084cc7e7d5f4f6aed9364a50e18e107ce2fd224b0d283f63f1f091c8bea82a70eb3b0a6668333c3f32c1b317c237fb9a7e6c607034ff20fe3db1b3dec3f2b5490c3d55b460ed41d296dfaa23c8cf39d513e55e2fd40f583eae55281ec37c7df37032c911ee58b2010300;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17649106ebf35d6a7ac5a176a68578f6a4c5902ac33a9a70944157161a0ae19ef908ad32fe7c7f993863344610da9b000aa58129c410881621718392d122df8d03606d4d77c12a6990111936e982a6b88d5798ce59af2a35468714303170a20f7d935789e11c0d573f15d23906803549d1c910caf71c199ddc4b3d1b93fbd7ee;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbf1c54b7759c9a621103165037dbb268d4d70ad4ee1a8b138fea1fc756cfe0bf58d3b86f4bec119e70c8121532a84bbe1c5e4665fe90b0c4ff4a63e4986ada116026553d313a8b291462dffeb3771853ceced090b87ed7216f3d61615d6cca5c7cb6cd3e96e9d9aef2d59238b1569059e2e1ea6b0eeee436fd68cb39384596a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0fe8d390906f54b9ddf45caaefc85ff08840e23288cb40ddb8061edc5442254c4608026a00dd8ee08f213627f92cda879cc5383c5d4aa1d95ad3a2a800a279070f3fd14bec488fc3557a2ca423374b255dabec977926a9b517bd656076409d015e65e40aa69fed79d923995fd6586bc9efc1c4af1ccba85323e83474fda79de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f01c0f9a0de4c3986a07ddd20a1f0bddc03cc6141535d2c0ad8772169e19797b64a28a81b747c979efd60ed6989a6fad125bc883de6890087e19a3156677d052dc74f0642119f2f04b6b610b16c5801ffe35a7202c6de2fbc285647f12a33ebd842448468e370915048998b85686dd008ffa65b8d67349ff675708fb14b09e5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbae0565b38b06093ad510c12950113cf075cce060704133f4c82265630dc422e82486c2ca270a91b5ce3ada04f78fb0ceb62496c7516d43306c516656745452058f546448cc41d5c58a4ca277e00c4677aa30763c9cefa693bbf72dfa56399aa83e48bb4991fbf487737c44e1a87234ba42f53085a34e9db451203a587a89e0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4acd0b6d88fdf219f113151d8822e7f18cadf3cc4c91136d88832145f2f3d18f71cef2bb653e2aaaab16a3a1f25d20d793a836679738848b84af1d7f44f94883c4993ba8f5fc0e42ecf0ccbe8d6c668e9ec4a0da7e51f5f7bbc2a8ca1c77af32f23520b1ed734089b37292a582aed04656fc90dfb7d754769fa075dc256cf3b6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb103a4800fa0c6d7efa8c95efbce0fd04304b330eff2dd5602534e8ff70417c93f86f0496fe69a1b460e153af102e8f2330e104d3038f2489f5d3c4e086ffcba996d9c135bddcd649f0e648030fc9554fdd0c07a5a8b0bdc0ada1dc43b622fa28ede3a6b2ef1f4dde986f9e74ce4a41c2b63d2bc9c4d89965862bd081f91e08;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9599f4b61114d49347233613bc809f7eb475f145a8dd46652926ec0cbfd23b640fba318a4b5e73065f4d726aa6d9f8fd9e3eb42bad91c4876b31ecd5500ccc44996d8ed09a861200a1705a3fbc743ed6970f0554f25591b7353e35a1a34d1e2e6253b49307999a09b600f4197b05a4ed00fb40ea21e496aba861603fae37c981;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec99446dc73756d57fa86913a065eaf3b1a8a8c57301d00184d18e9629391ef66ebc5e813fa5d3239a998028b10d2e7d1f8f0f1f6e46b96e9f26500d71d80949c2c16b989e906e8af6355a07ca835728660ab11e14875a7c29b668474cd6e9c48a4cef6990bb4097a33d6613279dcbadacb124a08e34db54469af98cdcde6de0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe0a8b7747c6d54e1b77446b224b725156bbaeda12dac67489d23e84436e4963d6ab9b3a508deb5499c2eb74107268df769fcf72b33575c4fce22516e471abbc74e952f489f339be6d075a9657cc9bdfe928fff31c1f8944c2bcccf086f38156101c1cdad5bb58b4b3e4f74d0ba822aaf11dfe829e7b54d4bbf731435d3c2dd6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6d7854257db2ef361eddd26f18f9c7e60be47703d3c425e57b32c6f81f4bddc61533e29f1e117fd94408c36fb168ef5b4496fe2e21cf1161aed330ed28f166badf9208b88db47d8b8155e59b3c924761d33e864fb1625c169ca95cfdbcfffc9cb5c5e43956b5fb5d40ea2a0e670713787e2a7899cc2dbe58ec2b1cabd1e75f1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2686836b4070a4144f9e0a576c1b4fabebf7d33a51ec2e3b0049399d97305d38b35773a718a3a2b80ed45ecfd9576b1ff4bc834b2d5c7edd9d7affd156ea8afbe45fd417ee1b786af4405343d77d8fc2e710ad452525f847c57cc336bb94450d58c0bd9f3b5505250b06c23bae3c73f1c8b90078b42a866e7e9c309aa0c5946;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h354a29f7f1feb1aa6a5054957ffcdce7f9446b6c2268a5163bed4fcecb063a7dfb5f77d0779700c4d97ede5f187df585fcac5285f095b6a79dc2457eec078a2231ac9c01c8ccae30178d9a9447cbd209ff09a4627541037f5236801e35020c0b462f97e239a7353ee4d16f5c0206184128b9c4217d3a01dda4f724276d3f04c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b384cad46faaa7c71d68257e275a788b3de0149f71dc9c16e36037c0172dbb2bf9c61e6a77f98d5205caebf8b220ab5a7d7d0ff93b043d51b86dff1e4ae920744e2055c58fe1bfb06095e35587f5cebf8885a57709848eef9bf7454506eeee925e7c28eede07d7783102a559b6fe0688958d04ce6ebd559021990bf48de8bad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63d13040a86ed4abfbfde91e945d2aefcb4afb07cc30490f8b46a21cebfb72bb9ed4dd2e134d6f90e68257333c7e59a30033d9ead62df26db89e1678e6f50a2f8c3fad3fac6e70fa13604d721eb2f8957000d67a4f19ec9b8aae86c183cd387153598834cf105bf038693483c296cb43c5dfcbbc45a366aac88f187c630395f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f69f74790be3e8207c0ed45fd094ba5339f48f7222aa872a23ee82f48d1f8e01eafe19ede00d1403d9f9a659f804afece37636fba583b3b1569860c722060b40f42295728970a45ed66f3239aded85b9661e763e6b1eff171f3b521ad4c9ce05d5efd5d0129d1872e9ef1c4530102d21fd22532861559e6128e1a19c81a0c09;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfcc9852b69a06911b6a01dd0a0b08dc74256f24ce5554109550c7f113b3dac61435ee705ec29def4a3756c5a7a6506d5b907b8451fd476f68565382bf0f4b9f4a9f8f5c58fc40e01e8c775f25152dda3f506882365d40795a56bc9acf011bbb40432732a411e1362df9d0429b4083a84b2230df494b0fc20914a047ac023a320;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4603d375895a0041f47b8e42948acd5d86c51897fc5f0c311f137c9f33e45819f807207eccb2d11c0892cbcca821c64cbb9b66ad0bd330b6ccdcbb26eda7026fca37ff17d1dfd41b0ba5836cb34024c1f291ce999d1bec5125796c0a3e9e81405cddbf1183266f5fe3919b27a355377b1a402a99196f73217359e5a4f2430617;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd7c9c6d608bbe08e4afeef60de9a2964ebff152bc89efc6daaa5439d231f5541f4b5b0bc7e4d7333fb6002be2b5b55febb06d6d62e8bf54f679fb158dbcb1c2f0feb1a1456929feee54afcde5e9b68af160adcceb9b460aa3d2f991bf0ce01c7d74fb85d3b2a6dec421dfde649b75e534155b5aada24e7ee2d36ce8f84875cf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb735487a551d05b07a6eba9c95e94cf4dadc8df85623a55151174d792bba2b20213bb390df595358f4106c9a82fa8f5eedb93b8769e309ab28e17cddae88e204b463396fe188e8cdf0835cdfe24b43e86bd61826ecdbcf59794e5fa280e69f17e1a188e76f6b64b2002695a545a21407b7826c1b0f246e3a6986346850a2b6ad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2db4ed65989c3f42b8b3e200bc252ce06c8fe5132999b0873ef79fc05ac80b8fe67c4e3d3306db9b7f4d358cb09f3c4fca3c75ed321ea2213a61640d9f25437db8f08c0c6468c50e3125d1d18d3723b7c4fc2f60b09312ca4136a5353eee463baa8aa11c78ca7875b03ed91acc0d1dc6f0d4c4fa9aa0b27d5558b3b335462700;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b9938617d558546c33355fe854542520b5cd1054b52e0701fe47a6183c8d399953857ff9bc544018e2dd0050b02dca4191aec48e2ac196d9f9cf92e84cdf0d80f63f979a755f0dffe42d38bbc1deb02fc9d6d7c90f7462177d32936fbda5c47c9c9a2ded993d13d9765b543a25351533b5630519f87af586ed1692d4a1a08e3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ce6f76878660bc754ff778eac7ecba451a2b6abd8b3682eccaea3673273d2f386386d651a763dfa0988a58054d415d3168f5e3a162cae0da7885d7063bbbc62d7a9de6eaca30653359b362c6cd74047b09967c3793a8441f2b89fa469e6d8ba25be42c8e0688bdb4cc34b88b96a753517585935a00bb8f7e8180091006f5608;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4de0035cc9e9b742999032f2b855bb93e7936e2b6630854f28bfe1b79347f04153a0217f8dad9e8bc9603283b70eb341a09a5b50a2970f2ac4dd8a99d98c84c8fb60d759b61c987e3302e0917c70488fc1ec4844bd9ee5d4ebf7136c4b5e284902ddac48fd3465f3541a3f2c3c8ef6b13e9af0958abb97b6568d8641361b1e77;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed5ad8ffd79ce14905df895927e240726c17040379f7d647264cbea580d0806ee4d4610dd58f36b790f7295957301dd248116eb5a69168d74062b046bb9798cb5a58144c768425d8722f377cc2b5b24e36babb1dfbab7ace8e6886bf2d4c9896e8070caaa4791cd7b1efeda43b9385344fdfedcc9547fab0f5938d80a1c1893c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdceef8edd5587de41cb2f685d2cc7d1120b54bbcef364785a1cae4d620f3f62d199d8c974ed43a65cacd1b482a71e4056853647f8dabd8bfa266652fe8487a2ed4b75757b3f2360fc80dcec32455ebb75871450d21eae3833793c3f69293bbb275712af4a4774aaeb0b7982d9b2bccd4666eeaa98b3070f060c310835a7b9abf;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70aee4c88695e877c01ad813250fa2c324317a1b49f7251661c29211d47e322b27de7a94f10ff0f04455af9b1d653a60ade51c7b8231d8470ea9684e28fdb205f5f7d79e0650025373625f859d9b8c51372151a32533da32fe20e895cb3f761e78089ab07453caeead4877f1660182882b8dded22e1650e2819501c6e6eb8ba4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f4c7984c2d85e5a0ddbdb4095b99404d3965e20c106c0436d926e835b967dd8d3f94e920b718cc28cfe5362ce0a635547559239cc29b8fbbf43e97d3b4055f2111e2e06fe5ee52d5563a9d94827d06c20ac75817a318e8f3ed7ebe7b677c13697cf3334380d09e07c7acd91ab8d31d4b9d9ec3def50ae2f6ed11d1ed5322bf6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ef31bf6ad1eca316a5634631790d7b46c60e228becc29ef2d8ed7f7b481ea7533ededac28efdc31d03791bc402832a5700ff072f6a75167a3c0f1fe88400540f1eeb934b2f0f50c8ad27745918a822dc85b7b6a4452d1702f4aac8b6945a47ae489c36c0c9f45d425e8751d45f2d285e0afcba8305574334674de735d5b5bb;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98bc63b6659458f994bbf1513444852d5d3a26e6bdcb256b2f21a7c8087c1b0d1a4566d03f7a3d9a74e7a175619d7972f86dcfc780d96d9ab5db91c885efb614fdc96e0c884bfaba05dbe438e585b463b520ac1e663fa7c6346609864c08f4be31e60649ff22fe6b1005b0cbb6b3f22cccac4d58c5dc18e958e9ba01a04588f8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb36dc8ccfccc29d49633c79012a361680da1734ca5dd12474ad86da5e033c84ba0dde68c0c6d4b52b5cc381e280c489b55becacec353cf10b4127231537cb547362024025c2b1517e6dfd527872d43afa0789a7a08482f5c5c993387c5e86ae0537b5fef072347bdff9073cf504a5c37c461d073ca33e82d8d1b4133c35620de;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e0dc552fee3a669a790c37ffe774c3ac241376875764134e6d4a2636f0fb04dc2bbba97336af79d84419fa6cccd80294194cb6905ca5e0665a73fe10715c645c2119fb2e4bbc985b47f31801afab3d7751b405eb5cd4f230edeed558c686910f3b1a067d4b725a483a45e0576a74f6f939179d1a57c1911a35582e955962053;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63fc873c847d21d517a8b2c54e3a9be6a1ae29386085033f7daefd02b58b45bc07f84d6a3c57ef6eec5cbb8e387ad3b49ba70fd4ae0e9ab0589813dd1ccdc7d01b13fe1989fdd75dfd4449f6076810ebabd588e5cb558365acf71d7028d7a1e4a712bbc8b28b1a567ce8fdd4613d656d7055228dc6a134a82557115921374011;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71c4895c9d8717787ef224de3c5948eac9b55a33c0ef84c8ac01d78af3875f0612e91465a97915aed449f60438992964d0d33f466a39ea4b19ec0069a485049d19ecb6839dd2af9d29e9b8be7f7336c8c0a16e666772dfccda8b0d3de8e24436f0ba4eb5e996316cf50ae2e8571230a5831b20ff9b332b3d7c9321de44469398;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f85bd23cddcfd73723ffc01b360cc6da7e850ac8e4e6266c209d241fb9e558d6cd4f95c17817a66fb6fb69b9c5ef2f07545c63a12898f081e2b7ad9de3bba8a246e2811f03416c405b3c0206a1622f6d79e32e4959515db182645dfb74fbb966ab722f3230c66c4769183c3d8ecd3ac94c0be5a1619d8e1a041bd9768b8cbb3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0908e94b19800513e6913292839c0f43663131293a4e6ed05ba11778504f9a59a79db41e7b3ee6d1f0d0dd9b728480c170ed0f1c7ae6c5c55026a124798cd3d210cb7746860976b120d431531939a7102b39b1acfb1c5fb7a5840612a2105a1223d9101d343ea50518b2a08dcaf90a735905a506d4a0b049ffc91cfc6267b06;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89be0b80891494260656b805d88e3c16fa58c88efb7dfc61757e4d1f618d402fc0c8e4bf96d7a59e2a1049e73668a4974b8ff984571193adcb07636a2b9e648763ebef9b2fd93494f364aa40c787092a6adc4d57ef9d7d66ef95294507090419e317dea222e9c8f6999649c42f60f0309cfd1178a598efd7d64f68cd27814a97;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e6f5d0110aac3492b9a1ee18660c3c419e354771ad2eb3d9d332cba5bc2c814fed3b2629e71680293f8426f14c768d74439f8a9d2babeff16410ebb33b7d8a35aaf4f65b5eca05dc6a7a9a9e923efa3e76b249f8bcdbba3cde54fdd3211fc41c895a1a3c511dee8a82b27553edb2efa23328983bcce0c6aa2f12d167cef1f9c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h263b8769b2491a06a224e80c91ad514797fd61c6519fabb2ae1bfbec944d4c4920cb8ac976ce260edfdb1bcd649f99f8a1e30cea5bffc0cda87a66e8b6e39566e4921511f775c789d76f493ce6c9097821ea8c04b5bcc04753681b9809cd47ff48e60ddef1f4b1b11896c93d5437f54542f2286504eeaa566f3d28a4ddba083c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b752dcce08327576044ec75a139535902499461b68649f1999420b8f6ce53797a2f84e1b4e9889c90f459f74bb75b57b3d57cff05de7ab11291082280d57bfc73fb2813a0caedf1cf46d6f1c621eb7113da3498a47c5bb89bd53085c7979b6c2eb3b624a659f199e0325285ce19dee1199ea9d94c49e8a2e489169dba8cb997;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9af2bd8885a24b30aec13c270a8deb6ed60d11957ed2485046bd071e0d6da8193259fb042e3e92033d1e07f829b29c8136f1000aabdab8033a20a73f63937581ca0256c9186296d63aec2306cfb155d5338175589dd4bb4e9d2cc9258514a7e6179e0d897d60696caba4848b81871b3304e09ba69c50e0a988ee10c8c6009f0c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90d89bcdc081d69c4562cdbe5611563bb2e875963dd9fe1876882929c2cb5237493ce7647b7770905aa648c34c2266f8a7f3409a856d5bcbbb2c7106ce2a63505731c387f74ab04b41fc1e53334980c047f8498e226a83c982195b60f046a4e91968175fc3d39afbe10cad11e3c0e178bc422c66547fd3e0311ccd8a87061992;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1bcfecb33bb98efb0b4aacce0d0ec5353bcdda3470dc5dab40f94687b95069e477b26420a9c459927721b6a356cdf416913a773f36cc276e614af1e67c069a7b0218f5bb07ae12375ba7073de912a56822754dc169e0a85830f66aeb7dd1e92d6a13417f1ac1313f5b45839b788457b2bde1c1315c83206ab416c5e7cf38534;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8518792aebb1874da9e9b9400665fe5f3b5ca5c4080d1244d21529acebc8834f474206634089fd5a19d95b1cd0b10c31538f6befcd06023deaa4dbdc0e1307bf88276a73f63009a0e0946fc5fc33575b417444a3d58a95bad3e140253de68bbeb760d8ba83b83fc2e8f1aa09c6c92c76ac83c0c66a82b5f4eb74ccf89b62f8ec;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23a7c8231a7c6abc63f94bc3cec244e6a5f0f838c2914a1f57f44e129763cb4deeff8b97c1eda57460789f516411baf61584d7e32ee77e7a74cd1e1675b236559c658f588c41de1af39fc706136b8c6f6f7aa9be4e963af07274de18fd802bf8339462568394e7b08ce4a073eae525d8e2c463026e4b0e2166deb99493c5bd8b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2966756ca69b16564643ad906af6abc61ea97cdff4148c0a9b57fa7a1709882db2470ddf39953dcf6d37f3a67f61e474d9fbef2759de5b193d4fb3c88d1d8d64ddb1c8955cda4cb5c61c30daf6b41e48b0fda4a2640a0ce3c5a884c8d8db3024513b08b57ae8fc699a4812f7d085526e59f8852df5bc9db1fdbaf031cf25513b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8be55d8cc5c7685c28c1b88f59c9254da35cf8cbdb70493ed95453a3e905358ee06efd6798ead3f1453f00898fc9c5e72d35cb6e86047b3098f36cec727bf69109c847a25b09adf34fd3e53e2208d4fa80994aaae73f24336a375ab40d67386742887f3ba9614b274ff44315d18c5951acc1d82fd31ce0a4416ffd516d974aa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5b2da9d3d5bb583546ccc122d340cbdbc4a1f0ab11a43d79093076f42e1746860caa54c4ea060085f7e7699eea579b1a8e75108863c3fad7d4ffcd3007baf8c5f3e2463ecb11aed836521473fa8d64690395a45615d6989464348ecee4782cd0cc38b098eca2109602b0ac3437c355f3124f1b66483a2c605484394531b5f17;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15c87575cfb4a20fcf1deee673c97478ca6e874841c3330977000f3f645d4d5d1c4f0fb710578f2dba3f595ecc4fe0481f8555b77ca1a2a190285c0141afe4c337ca8a08aa0abccd76270e6745fb5a3be7930fdb978b6be979a644ea43b6ce903f39c9797414694fa7bff39f5b04494c265c130b2696eea46a9fbc2e5cbcd73e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h643627489049b597d09885b5ca4a817c50d48c321a8468d3384631d5d8c97b09ac29da7dd7558974bf13f5e8abe3eaa83cf0f81ecf17b6f16e67ebe738a725f64857fb98fe447dc9c506b1dbaf44c060169bca20fbacdff3bb35ab58cd6a65d7d034badc827969416e0cc122100faed6620843c999aa1b52d39de2ccdcd23aea;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c6f58652e42536dc5273b20cd8d802f8f85e016cdae545f621cc90084b7ba64de9f8375c19b3ea331d04d1ed228bf54ca9e45934742d7f06a667f2ada3b06cde5ae06da88e81bf83effa775e3dcda6a520ab26f5762ea5ec26ac56d1fa14dd4c598b33e98c2eb45141303f2b4a29c858f3124bd8411c7df170698a29790e308;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c353191be06b9b7a36a5aa50929d9ebb9b6d3e1aa579b7e78ef7b4bdfe311a46dd835c3099cacfd694939a41164788aa3784480e006c3a8c2775293e4a3f028a8bd9cdf37855e84cc68a5aa93f9bf4ddbffe3f23d9ead7460b05daaf8901a8447dc6032fb16a863e13109d80db84718073a743762ff4bd2d78b7b4ccc526343;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d4f7de6c0d75c22ba0292986a5f7ea8e255d3c4fffbfda8f5bd1225d2118dce0ba06eeed4a986a1aac188cdeaf807eb0faa436002c90a66ecff554039f3fca7710d67852f24a96ac224890823df2bc9448471586a494b5d8024a81de1a1411eb633a325c1eb0013fd11ad8d9a6cf7af6165fb3e4bbdf43e6b06e9f8f9f63a42;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h491eff9bcdfdb42d58c07eefcf2aeb399f5b970e0964ed832d4552468741271b8374c27d5bd569fa7bbd1e248007552dc37e9d89124ebd0cbcb9e2e74c909ab4861c89dcd212cf2967910f86a27ea2fee265623713f1da85cfe25f0da30600fa28a02a3c89dd0f7171d4c14a12eb681db0be591108bfc8eb839b3d2c2e6c3d39;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11858ddc37296939484b6cd221c7e1514d84b1ab4f7f8c59c88189548d64bfe5c659e3888ead040f8d4a8dbdc9eee3b8338cf6f238a015313f622c01a87463a171d2ca8a542f3a5854a63eb7326909972811dbffff9674225827c89ab80030b7118fb86ca129459cb48dc3cf664e81506b3b93ed838eb502b82f9ced78828ea2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5be5f995afa3c8a4b1c3b5d6a74779b3a39ecd25127f605a453f5c4f1d7d0e53c77e46759d11c9f4428e1f0d6a9221525670448ef425c9b61d9ae40f01646e7db4dff41a85a60f862ce7dec9a4ebf95bf21851db2d37a9d3c9d043fc5d2a3e8b2e3421681acd95ec076faaf7436cccd1d16ee21cf78da09d23fab5252eab0da;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7cc18c1979d848cb3f04ad9d6e5aa01a04954e33292e2597fca55d63dd2ce071d8c8db55645e689a6c971db092b01308172465f38be7fc96ad0fb8b39544cb8ea253916b8a681c5aa4ede431bce064be90fed18a5c6e88f083cfe9be7b3703c66794a50a6a2b51d0728343386b649c26bd2e48b3fffc8f42818ecd5fc003d81;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f260e2999023e62b3931b29bd062c885f47951b729a3368610df40f61b9277bb9122115cc3b9df2fdadf6f58bfa8a2a3072f24af84cf26d0c7757554abf96b4a569421f02c74fdb1217b24941b19923525702a7993597f8a1d9174e4e09b1573e5378122b8fea09c276c2ee8c0cdc9f776c640adcab949c5f5c6044eeacc034;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7158e4061faf155599334532843df22e065371844b6f1077bdf5fe4155fe45879f1b4cc7ddf285b23b1cc62536b2a2329ac13bd39491fd751f6777720d69871801976f9c8c43a42f091a3d469861edfeb03b16f5aee4ec4c0797e00204f31ba9f42200adbad867941c5ac8186ed0fb85908ecf73953b3858f691dbebbc8f0ec6;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61e1c1eced0c5e5898e880a5053c96c51ee451a71ca9e3f4b3c76e999cd4c1713141a54e126f001bc96334946e1fe84d5c06a7f3615ecd841655b36ad1effdf669861c8e6196f48f497db27914ff13f3965d7e0bcb4a190d21ba72e050a65ae161073c9efda5fde14ddfbb44a93907b80e9435326034d8cec0a86c9b862af18e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb6c6faa500d99b14e83ef7022658ae153d3d2cfabece4b6b08bbff4742f89008e1b97caef72a7cd61b15ac2fd59cc80a79fcef944c5a8678f590329af4fa822e70f0350c4124dbfce9ff1e5dd9745c8b485f94767064c44c6fd57f01d76ceeab3968e337bb6148f4679bdce3d48fc5937f2503f5629ee4cad67d0f4e98d4583;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf31e52ef089da79c26ee23fd5ae54baff115c920bc09e6cef79fca7d29f34307446a33bc7bcb10b0bc2b144dfc8f99cd6f02e4d487f40f0a4ff6dafb6b854cc159a356dc2e7e13e330b860953ae28b8bed1c842037c52a1ed34af12ad63de43b2658624dba7e2a065e86fba103e4c0a5780f3759d61b7c535b4bff12f2aabac4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8547face1d5e321c396abebe767470c7cafeddaec028e0024610ffc4e83f937724794291bd3ea6403203d4e016edbcc67990120af9d41410cf5c4e236ab417753418f7c103871e478d50e6dcd9c3d46bcad8fc6c44b79ee771d04ff73c6e8382ca01ab571bf67a276867d49f8885095a561b5f1595991d586bc371a78282adfc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f90b3652283ba89f42e6f12361e5df9161d3aebbbe173f8ee0992ec3c8870f1a6ae80ebb2234e6f7c0c433ec69c24a6dafe24771c7cee1fcce08a08bc5f05a5091428e637042951d04814804ccddd8303ebf666e3f170047bd004dbb4b0186fed3e26b4ea00cfb8b2ddfcf1d3db6c86984b8dfc4ee029c065419ff4b2e2a5e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a8330a60be5df35e87ba4cdf7b651956fecc3d9c55425c31eaf511d8aa5f66719f884e5c6613a7e95cb22cfe09d52a63d3acf4173171efa160da0dd309588683bc3cac117076416969cae2a82851bf09c356c63f0b5f34048c49588c77b784fb85748d3006890341082a8971de297f5694948d8b97a63c5c9bf04a424048c28;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3aa92fbdf30d11131f2082d5b0b949f53bf84a06609c106a06345600318a8e58bfc4220e32d92d14c0edc997697bce1fe485cb01e22cdcd53eae5a8ded8df7e17a480ea3869f03facf66777eab2738f20e26c2acd151461770b1e3f32ab321ca6f601ac2d3611a7c0221318c77ddef67ece5775e49468562e63bf6b72e01fcf8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haabf7976dd0916274fea5f61e6c9f34cc636dabb4af32dc8bd410e7b4f896cc94be0e4665718909890fcb3533ac436b2ab99f8ca411c12170f0d677a22fbac8affb0952b1f8eeb1b4e4aabc6db4f1d1a9e801c939b899203a5d480ead09cef84853eff48113bd039bddd59995c5e5f58040dbd126a9f0c9ac93f260d822cdf83;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89910e8dffead8fc8dc3734a0b3a17b20eeed75b5a116be38e55ea8620afdd4fdf4e9beac0bcc8a93405554313855a510016ee9df4af0be6255020fb4710ea718b69306f4e4bb6cc06a9301f210bb33893502cd505e59b474c487f48d740dad67b6cfccfa19994b7c52bf125a2d6059191d7e734682675c7194da568db9fabc5;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7fe693c57fe19d37a8a963c926e54470d9cbcda4a77662dd51ce399abaa5867af57010eb3bd7598531e49f3b22af2a75afa739706a74ba842ad8bca3ba1a6232678501335172ef376613eb8e2c97ddfdde7824b34eb65986bdea95ea384af0161935bbdac408328615d310a38f2dba6423e69a9c73b9173de3b25d887d42be62;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he99bff5b336131cc02489f49e35d38e1a96652b5e79751a4fe4237fe68be0a9e1dcb6a6f0ba7fc1f0dae4500244ecb6f0997a11a07b10e716bf54f199f69ef5d259b495efe411b64c9841665bde32e0d6837c96d629564f2dbd052b3257e19cd1470c4a5d866b0f597ab65d07d70c3faa74b609dccd166adcecda5ff6f71f1ab;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd2e93b36b43ea7980d171d84d82a60aab1a5b6399834b139d7b43bd419d36cb05f54898592619660931956b1225607025e3f78d5cf4345122cad20212888546d147fe86abbc00934681e17119be1a917923c4442ac85a29ae7d5f8c39c4a7a42abd1f935f5037dc1840c6ca9d3598f42556e82adae42a90df178a0651af6dc3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h706f3ae8d7cdfaa0dc954455593c381550960704a5e862b568a6f86f5b492bd3c7354a01e74066c70b2f6be67e7f6e1a8b984aaf980e35085d56eed96c15e5741b200f190bdbf9b6c386461fbf75fa25e83715301dbb83ea62c410b3fa4de44bc5aa29efff3f50afcdd89e3460b7573bddbd08ee22c07660abb363794bb14483;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56e06f2e2aa24aa90eb30c77d4655a022edf50707264505bf7be69dbb48ed6e95000ec8b321838b41bb01890f8cf2c4281247843dd2cb8c58bf56267094880475855dae30604ca951840e892ea115fa0955e669c2b2c7c42b3474b6e03359ca098969b3b1698386b0da98c93f5e2a03d0b295ee9bb3c0c2739c55014b1312d25;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13c2b375482a1436b166f93d04cea1c6a0c6b3bc8e70dd3559ba53cff603b8875ff0b0a2fa7297930b0037c3d594b1f0dbad4eba56cf8eb282c85cdf989184b312921826e71d1449bca9485992e12d0812073a8f30f9d731cecd55006d0063ea1f0518891fa278905011d11e65e1e28139abb9e1ea6e5b4947e949a36260e3dd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca51f66e0acb20a8ded6ba735552d3110e0b9b33a5b5e705b1854912fd1b1b13834aa71199a89f6f20c50ddbe05b45acc7bafc97d0e55f22c50579d893cf9efab2b1b0faea62b7d69087777f371a96141b825aa3e639409dd950c922545bbe7dc46f8258c7f40c73cdf93d9a32823fadd5d3772ef63a6199a996a56e97ea249f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cdf227cef71946a5d398f0a95e1e09c41b310daa876698a8e6782daab53652cfc053e4ad2ffbbd65d4d34e3cbb1b4818755931cf16e4d22494107110df549b03fda9ae80c28cb718260248fc25c54a394fdf1998ce55e6e0d690446250ce99a863ec2d825561e70a460c356b6c711b58e4f79f5b826c6457d8863e34c8b1ad1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b9be2a00910f7c088eed237e05ca966397d08e0ebda239be0b683e85f9507c06bc328857808e5e85127dde9021d0160175da5ccd29c967a7d8223cda113e58c7cfaa7ba129141d4c8230e64578bb983930bf7cfd770f30ec9455508ed246d771f955545c23007085d7cd0bd7938d30e8d443638326deda16bb87a7ab9b02bff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb0d8b2ab661968188a8bc450f48ef46e5d9d09dcca12665c4ef933f2a7f95503320ae752a7ddd9b903c88c608f2b1f30258f72336d3b32edea4c47712378f2b34e289c85f3c819fe701ea315214114d601b3e4714bc8886395dcc393ef5704a1be4cbf91d5e934f955e30f9df13a5af374f84b449d65189d585451baa24d376;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ddeb55c0b5ac30a793144e7ac159109ce2b6e7d8d018cfbc57971c80d048f0a07804a4570e4950838956ccab38295ac4ce80c3180436006b0080d34ba2295b69271b0dbced5f2838ed22e9022dfe177c9603ea98fcd803b74aa8c7c8e9206520a55818461743a4318439284caa4bb1e05726725c36219ce948e99d71b89b374;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5209fb03aa44ea208370a79f9bb333b50aa621c00e248c42693e034fdf9ad24dd4c6595703598e9d1b4c02e04b5fd67b68383fe3ee2dd12a38a62ba805d2522c8d8d3b31f98fcb9b18a6434bff580e3c0dcf47aa07fb202fd19eecbc8a00268f2d0191b5970ab94ab130f75e3dfee2d0c22411c58031e446583ff90d92755df;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h848e7486cf81018c56afd99cf5fa94320db668c0b20b1e240e044cc464932bd4e23a3e846382fb27b41b44ecacce4d4f818397af986a5774ea93395a7dffca73d90e9e4df61b6fa6a38e65f9095fad2538e27a652ea4a3b19abd171d3d8d9e2f68e2842decf11be4c8ea4bc7d7babefd219102d063ae36cee8f7976c0de82c0;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h601d603ed4554a002664edd459767b35efd48f30284f86258b00f5481dc536cdf45612c7a44d35ebf86805ab5390f24c7e92ec254f4c2a505a64831961d980fcc487ad9cd74609f6735744b8724f6f7efc6cc5dd90c16ea69063800fb45c471e015175beb7b5714acdd6903d5c31bbe727323d7db450ee3908e89afeeefa879c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19dda6cf350db48d8fc577dcd49ef439e5f0d1ac11dc6bcc4d30ed010beda3ee46dd31bcb4f251c0684182ea36adbcac9c9300fcfa4895b00bb39b9a8d78414b42a91cb6a4867ed3e03d46e4acab97ec17953cb985a9a67833ae5505eb90abfa3148577bdccc0bd10f98632a3ffe58659978b25f593aabce298d6b5a3dfca92;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb08bab661f8dd202027665140eda2cea1c573856729ce387f0253c85b540f9feaa5b65ed5ef1247e2115f62b319166d4440de35289bb481a94bb1728cbe58244954bb5f02d2df4171bbc87eae9b12e67dad81513f6301ede9d26e72670a8212a9d8e83623dfba1363f13e17b3b7a5fec941d589ae219696ee4fcbc92476fd34c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h221cd82585dd29f44dba746a9d3ff7d65490c19d4214a9e10c5910682aeea3e41ae195ce814af1dd7364191e8db469e4eec628d41469491304966c26ecbe8cf143a3016ae49b7dd6613bf36e702500e787a6cf330997a211c62805374214a32352d24138b7fbd571f766d048d9ade950b446af90df6702d4d745b839a39c5d69;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59d1eb339b74ef11eaffae0c149d5e4ffb3f102275b90b46cc04840d1e24000a42af30092af7d451abab935b38fb205494c90f0d8368fa9f53c75ffdd47a1a88476b9bae151550badf80b04b902787a9925eee3b532b5ee4a6e256f7f0f9ca37a121159b7687f16a6c0902d76e19caa8a61c60bbf1099d9f73d2601053ce776f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5e7c6125837b287eeb63830be6e6c3b18304418a85ed93658bb42d99e7646966637c631756159e1bd1bd6a722b747aaa3236234c5d058f6f3353ce06c99f06eef99e32cafac174cb4d22d06c02f03fe961edf5c6e3cedae65863ef4d38bbcea0cfa36dfcb2d2a4e36f3581f7c3656b2f0d8122e70c545cfe339300fe3009e10;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7919898413efbaf10e0fd4e0414c81597430fe7951aea17202c0691cdd38f03484fcbba43d563da0bc2b6a899239055dbfb52b4d091cb65c96cd3985d6ef898c9efc7b748410128e79de5502100cd690378bd02f465b4ea19c2bd64ff498d4836afe9ff7f57f3650a2b5a574ffb3b3ecfa5f1a88822b97e7a381c360cf3b945f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45e24ac2f183d498739c20187e373eced757a89f64d037a71ca672aebfa92f00bc1a2bbe3c1ac920527cdcbc5081778e9113fa0b1042af2ce0d30923b3415c4f17a183592f6b19ae8e424fb207609ace843afe083075e56f09a161711c3783f06c441331705d1f2aa296e72f9796278b28cf1b86835668350f2a5bd6453c6e69;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48cbd94a5bf039d1c3809b0e5246e926469094c3141b684c51c5ae93b9d3ac11d88b19edee10632019cfd265a615cb790dea2cafc38fc0ba67335a5b4ea294433fdf174695236b377752a9e404ecc2f08a91f4a7fcf5da234c16b47a42ddc742cfc8705ea95a8b7e230e958e315acf69fc027d34676372f6f592243a7eafa48f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h945331088ecb02fe268d97b8ff1ee56a5a2d3c3c6c2aad6279671c4cb1192c9829dd1d1a5eaca05602067aefb1204d06ab2ef4af42d4680d8d696d1acc68bb86375fb8e85dd98a3a8ba316dee41470371d7c5037d2328b5cd7151e4bc0ebd664ad53304e9695f26cf70b54e69dcc51f95d5c7a516aa12930065a82b1d58d8a7a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb6512b2c74646dedf8be9cd9735ef2190f8b15d8bdf0ebef2c1d0dd5fcad32b6731bb5081f4ecd5a9d9b4e75663f4b055196a5e12a7c0fa7e44183e49f6ffbae53304472dd0e1d3bfca6a4ffd04e60b36537bc6a83de504e7194a6effd768246d8d351076a33b0be49b85d168013753af928747598b3f3bfb13b7a4d827b4b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf8bff5394040676782284afe4928d85f1614fc456de5e5f396b153c1c8ac6b49dcd8aa24212aa41ee3593cbfb2c0193f58c8b47f3e677b9c7d16e883c5cd7c796530be98569c7a8cde0802533888d9e624c85dabc43bf62f9953019bf6c06974c4cb08d079b65270cc592f68e17c1cc311d73c2e62fa17dbd9c080ba021e517;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79e1a1d5a9d6eb20e650627faa46c8a3f1b9a9416ae3792f6a0f51bd402a1e526ccd44adef7d2d99df7e06ec17c4b5640ee6cc8fe370c32bfb4ede113a1471439f72639467d322b7c1013bc906f11bab47c0e563843f36531122d08a3492c15749c0eb36b29796173d0a4ec675a2c5a52d2fcbde36615d4494c7cd1b939eef29;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h844ec32035e363f189a26bc8937195d574f8c9e316b1cf5d732393e810302c632078a0a59330cf8c242a796676caf01f0a948e3bdcd97621328669be49fc65b55940af8b0e67fc99860f501af4191182e316660759b517d485ae5ba3d16a9173171034c675acdf73b2fbc6baa707a1b7f850b3c92e4473fadbc573ff0a53e919;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75cc762c41e77b6b202854c4526a2b55f3c70020f0f5460bd75b1e5012da5cc5d4cb6a94ef8d3380e84fefde18bbf473e53c071fbeffeba5ed8db585c354c95f0114224f5daa752e3a7a839d9bebc3c2c49598e551b902c5a96ac48a9cbda5233847c14c23806218e4a008a3c9d42c33142e89758437901822d5c44ce2964a3f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h631452e61d954086ca90e48fa3610dd48a0da60e1e50036fb9d4f05cca0dcff22b645d4fad59716eddcb9baf3b799f0dc9511d5b5301d550e9b5e3d29ab4dfb628ba247416f3cff446cd32d0c2b5989029ddf8eff64b19baf9d254f926324c4ad40a14af6eea0dd170fb44c86e9423a4960611e68cb91fa41ddba1e96b6c44c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9af312dc79a6b03d907a85b9f3678c5c04e4b5d80d142dd267cebfc01bee249ca49248c37f96bc60dd1dcf057a173a69440c39feea47e133c69e31c622db14ca8a3dd9faf39c483808c70b1ccbd7e60202c55c0a36ec1e6b4ec94c393b34ebe133c05a8be7e85e1a0bd39132703aef0c4c5ad26bf2d354e41fced5362b7e15c4;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fda92a4f050855da80162d7132cfbcb22fe269edebe4beee05387c4b5c32d2179163c265f0f9852f8cfcb8c9b5909860327403170553b0ee9b7d20003a1a25e3ab44ae6abd1d9376808004ccae8ebe3b5e7e7412683a2f85b9724aa54fd2c094510f8266e7bc4dff7d14191573e653b8d97ac1f0f0397139e7ecbea0579df6c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d555a57ce4c730ccdfd003e38818b32eac64c96c9ac949edb94a9b3332588e8e0b972d6abbff3979281d083280b4fd1935e77791dc486a233e9e50e4b7cf26c9cf67544ec5f629e7a3286d8b3be33e3469467663fc8b1814afc5db7c2c6143eea679f1165f1b0fc44e56b7407fc7be8733821dcfb9710234272fddd620d8842;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24eda8a7197c0a4f9fa426f90234ed9dff1fed24289bcaab37b37d55019e0cb38461f3f332bd45f5417c0b61148aa523f0fa70f6dda63a58d9cad97db12bc72042666c63770bc0fd38e964d71fcde54c5e55b5878bfcda4425e0072a1d5a06022d2abc02bb295a27950b30a4ba59cf696e8a9c293412aa21d89c384af69c2fbe;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h936839ae500e3a7880f14db4d5729e4abe8ee924e3ce4a1929129eb76c7cbf4f050a3ec91712be7bf5de12ee4634c11f366244583f59807bf8d8e9484387f916c6ca4d5e1bfb1c8b10dc4e99e839fb1737a99d571c247a83589e5978c77f9bc4573b95a9d3d967a6b63f855b85e7f71623467c5c63fc10c49cd32ddfd7fc582c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d0bc477728071cbb107da7f839a61e5fcfdc833a19e5a86050ab8d95cb82d49ef5ff53f1cef746429a679f545951281dda12695081a403666ad8b6f9907343b036cabd734f9b5ee53c4982b835a2bf5fe4935426df254166abe66c0174f63991df0b860571ce739773ed1aedcd3c0d83ba75d095c389617f5ea245b136edb51;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he996ff0cf6064b27fb623ff48c84305e9199bb24dae0a43df2901f0bafbe61a70254087dbdbc6417caf2245b6435accddbc3e04e148d8b2b57f3b916aa13baadd7bce2377fc42a6e4f2bbe9fca9a6777da6a389ea16586a9a7c0f039586a81300aafecde67faf6000bb1bdb14b98842d458eafeb50983abd735f18438bc73f43;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51afd1952755d040cf32a70d13450c0985e3b4ceb537669fc78241fcab393231c5c7ef0d722da88651db4d3b425efa728d00a37b1b19553421838dd087340ef77c7c4a9bbadf3401403c4543c09d981e8f2a48acc94fde94f2dd45bdacfd611250cb611bf220b4b1eef69ff88bd5e624d6e3d3066a9d472f5d90fd3089707b8b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc4178d974205a9cb484072d782f8535e09939c4807c910233ca96ad893d24802cb79057cd6aad079f366544701f4b2f6167f63126c59e2281b0b8a81c944bc88172a6d7b3eaf9724d790f749ba89707772223d67adb77d5513c975e5bae5c00c3758395e50357028111c312b30e8983e650c8c9fcfb16bbdc860b17e5b9c375;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2159694d7733688dec5c606a496251c0d292e684141e5350a28aef6506ad30cd4d1bf3d44471a2bc3267661f4978bdef1273f7705bd2c4b39696f593ea9cf77bdaf754b0f18632f0fa164ed42103c4095e2d9534fab09f00ee2eebb1a0a223fb3b37d63f688865dc43db1a39659232d19db23bdd5a98f9dac81631112d0708d7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65d0ea814d90d85e9b4ca31165471c720a3900ff260c59c80784f8d29c9c5cdebe0661e2808648263409a7fcd4d71c6ec9322b4e00be976f0057da774a323d13752464f011512060f57d2f0b87831564ab65d55de629de922fc576ada7f8cec7a9666a12af7635b697f57bcd21395151206851fd47fcc8cad660f9023ff8b743;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a250afe7073f9a8f162f7b5a6f1440c7b3e2bd620fa9a4cb059c412944b1951af26712dc5e567936cd0f7a073216130528c4790bf53854316c01650d0423de8edfcfcc0ce5cf21ead6741b500c6a9b4ff6822f095e995e1337f236db285a0aaf59e16900a152ebf4bde96170120f3ffa19d5a01f185c357d2951ee1a17739d2;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c67f03e407b22c47675b4a90e9707d71df046df4dce6bf27a559d9e61daf1a55dc7966390857782394d8a9eceb4cfaf14c9d4dc4c872f943fcd0836fde5b4defa2d056d4af570b64ccac117626e44827fda53978a5da26fb9f9b2696fe26d597b62bfc88160b19cd270c75b14e839899a6bb4a554811607f58d6589160e5a00;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbc4ef7f428ad67b91c4986b9aaaafcb794b555c74906ff36b011d77ae544a6e46dbb3d682887512184a91cf486d06ab9f9e143007af4783acb3fe50a6042a461d3a880a0025fa868280de7999a0bcaed8c5717435efe35d60004a73c46fba6ce97c85e821a3c51b6469d9ad1126b3d4a73215c64dc974b8a0ee14b881c5eac7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2028241ba773b12ac665738015d7f21db7f10bbbf4fef648539dd931c1acded06e82b01af21b4a67d575c8f7e5a764d21c0b7aa8b11329260760e743f61e022da361b003caf9f94658b5dc9e5effb58a01a0fc2253d20a974a12094f53ab8556e09f9d5a4525c554ac74caa4fddb98ccd0076c69a560f235960c847f044ded93;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb31fababb003706dd8271bf4fd631bae51bbbd9f2172bbe13661864c379449d400c6a158beace63183201ff2c6eb442f9d591c341d8dd94e68b20b256b67629f3e9601eec7f453d95b63e274f5c9b6cccf45ba3f716fff328359f7a34c6fdcfb7e6f5b5a5a3b5c87d9d2839954fc5630aa47eeb3ac5ee7734392d9f5f06cce46;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed21a52dd56e6a7028e5a8673088cbd2ac42516ebd35d9f9377bf7e7354cb7f4a6f793ce0756c54c3b88a967e219dd7565b254ae4905949cab967441f1206510b7d356b9a65ec622cd609d711696009fb376ad39981f9f10fcbff9fd79042d8bbd55568a83d91334b085ba3c79526ffa373134b56a820dbcfa9fba413d765015;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf66ce1803b00a5db9a8b99f17924114e6d692f10800ec4a2315b68e06f28352a2a07f779c7700263fec49523174d3e6d16185086dbd18c3951fd911d80fb088bada90f036a2507f6d785da18d5dd439573c597299d1672c8d9e5f5df37206e9ef8a7724b62a5652289d45d292ecc4d5282306c0d2149440a61370394824b1e7b;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9ba01fd00148d9e2b8dc9bcfd8c3c01146e4d28643948bb9b67c5e1b1135868c7f7cfcf222bd5ea602bcd1f0b7136251fd5c9e2850301ff2808a99890ae531d471452a8bc7eae5ee6483a1ee6ea42531c8681cfc8cd4206abe4c70e1d63256800e86ff1bb09903d37fe5ff126fca1c0d6659d20bf8461a69209b6f4869f075a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d6b0c50b2e966084e86310676c4e589934b4b443947ad2e4a1b82b971f331dd99dd34388cec18238edfc9d7a4a3277a6736bc4f5fdec6adb7d3628e853bf1991876d29724f29441274fa2c65041ca0e1ce8d9a24c6cb6fd924cc3d9f179576fe258f2f992372a164a423fec05d42d63252e6071f727ecb7b9611b5ddb898e03;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19c9029b9d06a49eac1572a828bb21f651217ba8bfb41b2c98a1a5cde9e53aef04fd9ef0b60849d3a24cb9278a4077d8b53fc4c57deabf30293c26de0cfbfa7c7085d9314bbf78a9f2a5c83bfafbbbbe179ddad80584e9d3680aacc4fd355c2d3e3bc243263155c5d033d9ba2b188f554a10c394d07e064065a31c44c00142fa;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3d85b4a5c6d7864b6b2f581e04b31064f33f1d83f3d39ebdb5252e804f0b0e065d2a8a14f2be690f6a5c5f8244417d34d50d3ff1267f4b3fb1fe6b21dd18ba378a94417f0162d86e862df5a76694533844110f5e99f4fa16a7f1e3653d93e75593bf3fd196201c4447a260c253860dd2e2f0136a010bfc3a42128b01b14af6a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h505199b739efe2800f72f6be1ff470273c19b5a35905c7a322daa174a088410ab7930ac6c595b877854cda68d4f9d13d7cdced8301750dbba8fec1edcc9e99e7bd59a4386186ade5b5c1e7b6bffe944dd6e9e64ae1403914445604eab2c87387d0494349effb7eb15ed6362acad72352aa53ba6176806581bdb9a2af3cd62c28;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1faf144393615e0aa3345e49a87195ff8017f053dae6f8e569f754c42f065b5f7e7f1341c1149f7e3b8a1b70572d40b323cd6f2624ca394d26d22ecdc5f258503cdf82ca7a2f8ff13d75e2e6a3803cdf25af41af13c52120bca73fd24256d37d54bc92417918c8af0d59ae4e1db9463dabc88ed088de9dacec43ba9d5c81864;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0146e7d23a5f1e639a7a4cf9c85f01475f7c39a35d7f9863d990c464c54043d0b5f89300581190a1d4c4aadf42484ebcdafb0dd2dfffcbfbb7b748d2b42f9c00d15a6e4a2ad33d584d8ba192290a1c56f241d327a695d120d6c49ac6d78e2bd16f60860938832c3f8d948405b6a188862c2c7664f0ed5f3cac5e7d5df0eacde;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebc5cf2bff51c11dda7c6df57088fe4f1eda5e423e944468538c4982348772c8809a60d1913adf585adbe1e151e70b716e4d931bf4966b4fdbca8dbf8ff60a6b2dbf1d91642e3310596c6cead924cdcbe15fbac7d1f3694a7ef9c62cc2a3945ba87ca016a73bbeb08b03ae05710e465735569251d54228cbd0cbeaf53409dbcc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8791443fdc0c9a1976e1f4a09ab2648eac51f111ca5b32f68ce0afe85e15f92bd85070fd26cf54cf7e60538a6eaa342dbd8120fa11c4aeaf9f93ed59152ad6d1e5ec29a367234ca776dc70928fda713480367ebbea777b68770d6f7de94b24eac7d7c60ad99db500f7652de8a784831cf357f1ed54bc47f718bd09de2d09e882;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53ac972d760a865f949f1a1c20975afacc84a09d1d8170f9c9523095378fdb01c8faecded1a21a690a0d9ac6f68f759b5eacef5ab60e925193974c07996af5e4cd16b0798f74a95e06603266877b7a79af3d6e123401b477ee16bbc1f5793ec54ae33c7462f1d3e52a0050cde7a3f32db5560eefc0df9e2066b1bf876775a507;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcaf9c145eb5cb1bd651c992440b1b5770aba164295e106b114aaad99fbda458654a43b5e097c06cdd112630f6f922d271c3c0092762ac2678efa299015214ca823110ed59f2c88a0f99ce5e7022b771f46708eb9dd862f4d7fd943b9afe6783c5b343fcf0ecfe81f1aff0e115dbad073cd0eeffdd90f6da94bd74628bcbee728;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd33d70f419d4dd3f7ce372c65c22788a0ba77089a0eba75bfc8ff4d1fe152e2bd156223bb6e9f68045b7b919da58311901ca10426927bc993b3f35f4842b8f2d679a09e582ace33689b657ab185bf70484ed8d13d4cb9c49afc08a0dca5f6c6a71cc932fd2e22e3b8a8a13b325e238fff24b8d4a116a9fc41c465cfa9d7491d8;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda4f7905817845b3d79d655157409c0219a03eba91d75e2ba1dd8049c934295eda3f311a587af3e45378f0dbdb056b79315db92772f72238464f0702d2a94858ca932abc0ea834eb485438ace4a89caa02f89dd986a4442626c90451ca1505f3ae33da84431cc468d2a86d2f81e9769335d99daceac9ae23d6d4d84a591a000d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hecc868935339376befc705ddae302eb9e7d36f37068fc6ee283d2da794cb07f10651952a35dfd691973d179820dc0045184d6014ecda4cbb49d86703518f1abb2a781567098a54d424a89af591220a5dd7e5fc0099254a7d53ef4286af2c9ae38dd8f8ae33669edd3bdf78df1854091f8d33843e469b8c3b3bae1f18ff06e68f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93b349f3e3d8b812d1f695647f1e1363629f7c1aaf1f74e52dd36b463c0c5c800dd7a479bbf0d81cc81e7e527c113228ffd77249fd2a37b7e766079a76ced57bf811c8e13c25049b603b05505698bc045f6f2d9472be7738f9fd44cef324978bb2b7068fb70cef9b2212e5a5165bf5dbaa39372a8ba9e419a2d0ce324a8c9680;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2992e21219bfe4d46508cc8df3cf8885bd5602713a779e1df1c497378e59da90708d627b9f6bf8f3942b411a6b2b1df6f2317de3cc6afe5d40897ac35605edbe36014990831024202d6a70ac4bf36ecedddbcca70c0ad4579fdf841b2dc384f2d3eef93e1fcbb7e48657509d27acc649cfd3baa0ba6c3f08b8d6119b112cd143;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha26f56e199cc93c302d5bd6eccb39e905bae4f53544b1634b9a11e8dcd29553844c9630fbbdbd3e865acbe343ce312bef64a6c6738dd3d0f8ac3e3856b74ed2f5ef9e869bab1b73f4869a2145073d60657a93f4bdd7598aabccfa4e607a33662b74ea3e298f0fe3a86ebcc26add5ea7efa7afad503fbff23a2aff6b8e1730c7a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f5cc6bfcfca220de8a5b06c20cdbb9772502000377d77b0acae0d866ae292a72ee8b25c15e8059fc7c7bf0d5d53035ac34c71ff241601d88d15157a8a6eaaed82133e1ed44fb965553a55ade1f0a841598837495357243971a796f0de8bbe9a32266e56560acb018309d05b238fcbb72be43af46d8b0b130d64c5d3f51dafad;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b9ab70dd414b57886bc8d42359c2083bf5e9d228496935fb6db2967948cc2699545671919e9e805478a9effdab34eab60397b960836b71b48df188c8e8834bb1c7431641b109843bdbbece0f85c9d067cc9e96454299bbe74b5375f4964402d86d47843f4bc5375fbcb31c8a56b27ed228230c3e85ae06c7e2e7bc20b992bef;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c1ed3e929098c5ba1bcbfa1d2eb1a087aebdf6d7d2ce75b5a24df7538b76cf4fe0a1dbd208462f091c8039c1769c91f732ae00f27247090376f4495efa4ddc688980dcb1c11ca54254ab1f400f1bc2a4882c5fbb17292e312e6434617e7680bcc7b6c19669fd6525013d10fc2e00e5a988ca008b1ce72f934e3b4686a0bf040;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f4d8222018f889290801c0d1043cac4b5355cba3a27eca2ca1cbb1dcb384bdfd7d1bbfd178f92fe80a100e22426c2fe57739858aeb18f0b5af9c887f8052cfd3135e993a6f318e8ba589fe8f15a1eb189d18cf943ba03ca2170c3892d59483def7e50c726708206fd352190f855cb116099035a4573994decfb4fae26b9a32;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3a15145c83223f49406496b57a07c8b091b53877afa1ecebc35c1373a435dc3bada4e15ef760fd214c705666b711a3909de43d5fcb9a7252f4f4ca3a26ae6469cce7f4f84bd2e0497785b2e850d6b340bc31680e0c20438e5802d5b5919f8fe1c344f58860a8927a660dfcdb94c76d5b0fc01850c3fa14e4bae5c9538d651bd;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h852ac07e277dfd6bae948d82f2f028025cc94f94edead1034e5c6017243cd7b23c84fa6e4d298274b7bf6307adde2a16e0413999513462567350fa70f0ff452fdcb71c2dc585ade9fd62f624cfec316edb6fb9eac153502de01261b2bca417dff5284f3282f7408623649c51c5c12204fd1d33b18e6dabb38b286e376708d0fc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5967fce57b1b4f988a8a952f0ee25990095ba92c4a99a99a91bdad97d5104cb72aa06a4fee7ca936cead632ecd5b6591f4f7d8fcdb8efd2f4d2328d563bb436519dc2be3bebc64d70326b8da244211ec011ad223395ae7887cef39b718b7d37bd3d63d3ad37ef7549e9cb8af2f7fd4138dba6ec74804d075c5555ddf446fa3b3;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93f855159af2f5e3a04defb5f25613cf21d79656da219a903493289ba1a9c237c74f24f436f14e9ccdbc368b702d9b3d36bdafc47cbe3dfceca6b85191cad24f2bb0a2d7239c03aafaf81fedb700fede92436ffe1fbe5d321c80b03414142b838705ac50bd98af888328aa6e78b6ed776f8b3b9b3b27044dfb241dbe204a8bff;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h166cc7ffa9db8fb597ef2df5c736f62c9fb1ef6e14bd565d9a47e64bae1876a0497dd10eb6fa447020ba53d907bf666190a39de418ba09f2137a8b27bac6d61df55d245e2846c81f1e921aa060182b33733fa1f3412058f9f19d8487d0cb5903dec505a0af3a8034030f2bbcffc09828b72dea5da3bfdd2e808a5cc408315655;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b75d15c6872d1ca27fc88fba4028d9761102420e10100ccd4524e111a7ab021df9f2c665a0269073f57ce6e61f7c7cf51b72b66d04a6d159639b76e9914217c6ce5374ebd35f656c7006db9fd4f44ada8f819bebbbf12d6cf34ad7d10af5a5ce3b787bd35386950d5e4158598b20ff6e770a37108797e66f85a74b5f84772a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9c88f86b05e760dc86a6b44615afb5e90b78ecfb5cf45f9464149363c9c491636e9e36525303b64d897b1cf45352b1ffa0f19efa6865edeac47382c81ed2a41b90d7176221c5cfb34b9b0f6781051f5e4df8379acd1c556b73d5d59571363e24b387f108bfdbbb5c14895713a7e304ff13a3cc345b8cce748c3fab533c89d12;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3465bb814d5969ce380292ef0b52c11517deb7fcab7808306b2e9af8b8265640973a8bcdf2cf5ad57071b4e6a1ee26f1bb0ce9c293175bf6e69dfa0f8dae3425ae6a0409175e13d9b0ad5eb28cd7a299a823b9f91a9f692653f27c96a8facaf8d2b15d5e7f8f670f4b7085e217afc450c62e3f3bb20f2a0ed3a4bd2eba7621d;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc95806ce5afc02bcc9b71e5ca6f78ce4472fac88523d9de965f46b6da65329585232328b9cbfdd5178ca5756e4427973aae7ed2c4c2d65ecde5669d185eaf8eb192100db32a0be049e9ac62babb694a24d7848fc049180dfeb978955b423c9af4d29ef5fe9636299f3e983a8277c08613742c41f74538cd761d06a3a4b5180;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he85cd86d388565a6b052b81b19500e3e436d2f42dd4c12e62f86f78d78496921d53913cfb6df2f7b10b9dee2b301c56083cd1398ceb8961bb05958d6404829526f8b1ef1ab89e159e53ad521251ea85024a2bbecdc862e94fcf71a8887d5779e883c322fac32c2cba05784b027bf390b412306f6bf723eee8997f51613ba179c;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cb215c842ede88f9960bb4d5a6f3dac945afc3125b6e7480d8d7143f3da43acb827013a341da39c0cc7d0bb3eb7de8e525b32ce0f89b323abca1149721091f9a081ff13a5ce15cb03874a2d3e45210c1cd56bd73b0bfe70318c900a7aae611e75912c50c83f621f8d4d60ace51d8c01399f5889305af4b5878ea5454472c1fc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h902155e71770e51e897aecd598cb72c66d17e0923bfaaf523598f386aca155842a4a95d050880b4d46a7e054516df6f3033443bb37cf3bf43e926b5cfab931649d2955518fa514f69e0d169eebfe6815d4161803dadc94367ceb4c8971dab7e7d31f16d547df9190ee2eae7b2b05a3fdb04a018744b7b15053c9768dfbe7385a;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97fdb3ff58671538204e21da4e60ca62cabb454a9e2e78ac8e84bd1257ca5ae0d1d718e68ae38936d5192989c92665bf8ae9acac4f5be47241112ad00660812148ba644c18171b14f4f2296b72edb31132db61ece7a295e90de91ad623b0e49c56626f1fb6c9228762cd97ca58d8c2628ccca578c64cc00bc2910accfa382b0e;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h804a05094d002bc586eca84499e9147327787828324347f74e201f77c7b065cc7a88555cb1b095491c3f990edb599b52f4754b7cea4f5d043feba5783f461f99f6c345cba84b77db85c757ede71220514de217ebe2db22d848a39e21b627ec5b1b508d20ecc387b4ae93850884cba4e53cc80342f7f9cb5e7109cb47e1a55a84;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54d09d85b3494bb777bd5dbf27267c236b20d86d5dbfdd5d17146a36c5ca7569ef50fced4022fccc5275c62509a4a8332a3bc1d7dfb50ee6010f6f643207a95a32c2778ab0966555b6fd738ef36582be2c7b3f330c8527cf453f2b11b9df179b0558f0e3f66d3a2af3fceade255784625c2116428c2b4296734afe1d15eded15;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb988f225169e24541340f327b12923d7ff295ca15ed7b0f3db4b59439e01886c3d06138f1ab0ea25985710de431e035d2d677f64ef5a15234fdd79b9cd09a9af2812b82f9ee6c3fc5fd7de09de14150e3c687ff8f25fe7d74be8d705d8be6e6dad9f385b5fe2fc376e7e05ee01861055bacda9f0aedb183b57c269b17933e65f;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf64560360c19b6a790bc63df56fd5ad1b827a18d12829a7b5b6f9609b28572adb5c443dcc0ed7784658578a1bc8cd2e3d6bb9ab5b299df824c851cd15ae8829f640090ff18b1e839a334fb3550122c6476fc543d17aafb497606c0c09ffb4a270a5b4140c2175afcc2dd2fe807c34a5531763f0a2275ca27add518afbaedc78;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca2ae902dd65436677d3df6efbdf9f42d7ee1687fcfb20700121a3d2c08daaf470355971438f488129204be4d731bab081a9efaacd14a4127061ae6c925dfd7aab58987ca4e0db359be601d1c328e62d911c2af862ca71457dda6f481c1084a1d121a5259d5d66312b840dc775c9c7c199710b1acfcb9079764afeb99077dd64;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h847b4f9d5f9936360e1f41cf2a104791f9426d9ebf4fb0e5d4b0ab8447b71483b5ddc53ad2c250b042bc643472cb06e6ed303ea56f1004b80726cc1d9903f41c6837e97399d5c8567a1e49af737bb2e776438ef3020ef8dce366c4ae344e7b8e19902922eac1e184d7b32233ef41768275ca9cd2d62037af351557057e0192db;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb072b64d4eb00461e219e0186f6b5f446a3fed68837b4e0c24f0a182d9d13719a703a6557ce4e8d38fb6c8caa899d1738978ff7c355ed78eab81202c46a24211e15e95ce60db4569a1b10df958c88683b8caa3a3dd8149689c940e9a203ae0cdc801a10f464b6b947dbdb61af67bc57f6d6dbd5c93da7112eef595d677ab0633;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h603206357c75b0451d3cb752271f4f8b63bc64ed68b054c4395f372846ac808cb5a1023c62259337dbc8099bf217a28f20732d8a5fb2ea3cba719218d5e7c3c377bd1c0040a4ba1465b1929521bf24291a43bf707d8d612d1ebff372dccc27a50ffffb75d99ffd38af535908ca87b9dec4a383f20ef9982a6f20f7b844416206;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41ca8305f0ad245b1b18dea48823a4b7d5861891139cd2c0d2490273106e5b24ac13f4d36b223685976b60453c4b2bce51aef6e1f2d9b9bc220bcf61e1a46ce7e3911e917f99882f3c7e23c39d71386623a24a47f19b8ba12432d4bc9b8bd9a7ec5db0a0d6d6034d6177eea418f980f6a4760162c939a2dbf7c5448895f30a43;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89f3bb6271a4aa344d3ed4d6d4c666992245f99355344b0fda2478174e6878c4b4ed8123a0c838886489914ddd9fcd6dc56ce5561bfa8b842b63bcf42233c39e224d7f60887e17efc772dc4500d8cd722f0e583ce16a7572edd124ebb5b293247cd4fd6d92535b4ac94bb0fb73b3aba99b3a0bde6e147cd2ad1f70eddd683706;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haccd68f605ff278d23188fcfb01aa7e33b5750b29f142ed9b4aa390280a5e9f6053e3b4696145bdcaf74b142e81b8b0fb2d102ab8980ea0569be682d0dc3091d58aaf8b1a809b0a823a20ada09bddc11c7c544367be2cf112b646b37eaa86583012a6d625d6537f0b30a78512427df04056f0630c9a39f878acfb421b9507929;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6b3067519f07b5f5a3dc2512539cf2d7833fb36b391fcdf3729cc97ddcf0888f257541e5fe1c8e593a1dcff27a674c6fb38b9669ec13e2fddce9dac4063564fee9c5a5d449cb76f88b3c5475e188e6520a97beb17066cace6308b1ee1c8bb8bbd28be251a3d25ff04d93ac255cbab17367d6b9b91b3389f2cad03840ccec799;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67806d817f6847c4313d7dde395f296db27ccf388004c491ee6a4be84dcd06073b3fb0aa138938a850ac83d41bdb519be55ebec9a1c97af5d369dd512afc4c6c2cdae197c79c19c43aa778076b861a482d319ecde80397172ecd1a169f7b8a988815512d7e74f35447a754d077556351cc32fd9702f076e1f4f188c8632f83b1;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2f777bcb6321f9fb32ae4854d3efe5af50ac90660900f773e87398c5615ddaa381f0807f454b6120ae071c4cdbf2187226c22bdc97aab4e845685070af92b9d7f616b73ae98643444a2708058f7e07e1a4c4c37941eb535a83d4ba95421e563841ce5b1e90aa244a6a7def5d4a58147d636cbcf0f3283ffa53ea3f37cd93b12;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h614585b34a53da97ff2f27d5f2e4abec510f437eb27cf72d0f01da563041990c256f01343e76f4793d854b25f77ddcb1fc77969b17cc91e6b1cd09315bad5b4a1b9276316b96428abbdded771ec396be6f6d284d2ef95bc38ee619e247054382bb1dcaff3d01d9b96707e74a76609d152cbf718b2b5c7671c5abf83dbbe9e801;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb01c0dffb8abdc5cbc33970da8620a6e3c5eaa3d4340e55f74285ddb7c87c5bf1e497dc00f713b51d59f9cdf73061f038e8ab0c671976c51998c83799d303ba62eeefa0b8daad2ad0a77f6b3c039a30d7e5c70e0fe8ec92bcc485bbeadb4a78b5a81771bceead6315bb3cf043738aec02f926da1fdcf4fb2f3cf8d17c2a69060;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12ae1b27ac237d385469273179107cdcf8bdf7695ba6da079d33da82fc1964eda78a643180e63d65747ba8c50bf1295d8597d94525d691f59d50584680ab43807787b75db46283082bb26ec596875f1289a9c88642d959fca5691268a092981dbc4b4b59576b12ff475c553b74ecb3cd7d505410fd0a56478dd0039e5b64bfdc;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c012fcc972d43f7eccb7eb10dfe30fe389d878f51ea6f4cb9833e59d4e0c65862d0575cafcdb3a6bdaa221ee294ba90d0d77690ca7e2192a97cf347438f221e5de574d9bc03bc718baae5d525609d8ee0b212e3c7159bbaee4b91af989c67177bf9ad595468b201db25582de9e3a2590f9e58c33046f1d94c299a70c2329620;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc72c249e17b3af3f16174555197bdd7e46657597ba0f9509c44775f9c497076911d99c4e8f1304663ec5078f045d0eaaea03e6dac61b2608c8dcfe05e4525b6cbf1f7f93f666bb0ec06fb384ebd4be0a33a1428e9cc5de7bd2621d2a71fda763adbe62b288fe59550f9a9b6ffc4c126deac326b2177654552bdeeede0f9436a7;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1584eae574c61133b2cf2a2f6794cc68622c05973ce34101c46f1e598dd984e119316406f93c0f9c0106de4d4fd38fc22672822a779d6e53976e3b3d9d0c0e5bf4d3bb9f1f8915b65b4eec9934589d87e1dcc36e7e6bcf16e24615922401a0bda3cd0dbdd90d342017bcfb6c14d3ae6a39d62057af902b76f1a988a325e86477;
        #1
        {src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf842f01d24576047effb55cc7b9ee13b555b01bbcc2b402eb92411db2c27dd8851ca2e07b82b1f50a57cf206372af8f9a23ff2ec2f6ed4e287ba985dbedfe615dae8d47ae0dfb61f474233cdc3dd0916815f62f20e1d3d1062fae9b23194aac9901763ac7ade205edc61c74ce5e9f15439dc5a2afa50f74b38b5ecfb9397dbc3;
        #1
        $finish();
    end
endmodule
