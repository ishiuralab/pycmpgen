module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [7:0] src9;
    reg [6:0] src10;
    reg [5:0] src11;
    reg [4:0] src12;
    reg [3:0] src13;
    reg [2:0] src14;
    reg [1:0] src15;
    reg [0:0] src16;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3])<<13) + ((src14[0] + src14[1] + src14[2])<<14) + ((src15[0] + src15[1])<<15) + ((src16[0])<<16);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffffffffffffffffffff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h109da3a3df67b54e39793;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d8c6b7437a95f05347d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b1d1ec0f20f0fce70b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac990b5182a2204bd052;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b231c35f9f9c40988817;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf3905cab8d4f9b7a4e20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4638bd3d7d8ff94f105;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d7f1b98761fb15add46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7abcdefd74a7f34d101;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10b237483c4567a52bcf9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1621658a9b13e1c9b8076;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1531e5ce37f73ed917a45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6bc034ec0a5342ad272c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bbdaeb7f14b43cecd896;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9733ec84efe5383a3ebf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ee87e44f5de3a48acc01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11911377e78a21f45fe5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha248631096e7a1bbc789;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f9b1ef40f8bdb1933fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8b0e002d405b98d91f7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac855d0629677f1c88e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h62e6960837bb65b2e0f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c5e4647f9713f8f6a1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aa425f2a629d4c9996c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1233b5b0af7b56cf2621e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfe716e69f520a129c6a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c755f8283677fffecf7b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15943d602931236087e90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16147aaa5ae7e443d8f4c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c5610d8ac2e13f996fd0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6d3ed480737f7ffda22;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h133deac920edbe3d7d4db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94ecb3579a162f78ff44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6e3a2d7c35b7dbfeadae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f7d197653e0d76b84a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1602acde0d5bd2f36b454;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13f96f8c6638588eea852;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4fda2761d63c82dfc8ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1877c27514c513a941ad4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd229f131b1d538f860f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h159e453c17a3416188c53;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e3cc93e43a73f872c05c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d557818a2223d7381f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d5dffcaf316a9b8442f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h531acdcbc693cf0b2c80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9db8cf862bc12544cf0e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114c1c0ae5389b9f85662;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105a0e37c02560d8a420a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h96028977d37530b2a7cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22c3cb3768df10e7a5f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfef490c831bfebc33e9d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d4faa4ff9fe77c49c13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1270fa7bde009967b7822;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ee356943ae5fbaee343f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h808906e9327bb16875a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12827c17fa7fd27e79443;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa1411b0ce582349ae6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfc165372e85599c48062;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e7ecc13c2662a8852ee0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha805dbdacbefdf1b8d36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1042c5ae12c38a7e2e02a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2979c2de5a542981c2a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h136806b0c8ba0e6fe8959;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c9c2d398663fd5fa171;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1376059128d3c700c2597;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a9afe770e0d6319ef280;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6dfeda805281ff5e2bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce6d8409ecceee87121d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14eab26a1f6a1d5cde0af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0987a4c7fc8288a8d24;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h86536d002c39403ca2df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb665542e62574ea42b84;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3fa0f0d31c90afd29695;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17bee458f5c9ec56058e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb283a56aefc0287587eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c270f914db033738259b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0bfbb139b1ba951208b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16bac79c2021766b55bd3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haf193c46585391fb3832;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f0de5231fbb58fa3695b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d33bf09554a324f40bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f558af607310c1a69502;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffc526bfee5c66e26e64;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb90040a1dc3129c687b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h98d68adc0dd2354928ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e20a7d0cb3050e88b79a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h126dbb6d5d7d9988392dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'had01e8ce7e97133691a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed56bc9b28490bc82c63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1964fc40d27ab6014050b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8c6981b2ed025e6271f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed7c0522ebac883f0351;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea4f10c363a5ce9842e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ae0d42684589bbbf93d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1375296678297a368c911;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2c085951ee805e57434;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he77544833652ed6607d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h685df03d86fff90ed9a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9fe671095af954bf1807;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h142bc3867329ee032c97e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1459d9159eb5dd7e50037;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1334f2feecb38e049c696;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c46c1fcc2ff8f0b1c314;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha06e17b2785be0a61b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b72681f4b23e280b175d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h853b37700707428ddc5b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bda70f7a563445ca5427;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h37ac10f9da235c88e5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h40f21a93f30a26144ffe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hedc107e44f80139359db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dfc4dcc0402006112e2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4746e9bbc5865e4bb57a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h167ae2f55edbade681967;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9c78b181d0864f6f69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be90f9151d93d938ce2a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14e52c66a87d068621cf6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h75fc685cfca326369381;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1847ce66255713f938403;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1878c8eb9a76d2e9e9314;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b1e028048bc0c5fe9664;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1730228c34097b22baa0c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f84f9b5d5bd165db76ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1238b175ef13e4210f401;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16cda9f7bd5677aea8d91;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dff793ae7f243debec2f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h96dfc6ffcf989964f904;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf854885cb9ba0ddc436a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he7013655cc8e3dd08ed4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h128f0550249076b57b7a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1407df4359364248356f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7df3de97f1c24f1960c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c36feec8004b6554286;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119ce2f056d1bf1010415;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16acc51a9caa5343b9c5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1075d7c0086cf6377b693;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186e5d8894c5a1c3f8c5f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1857d9b51d27f9d893b1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e3901c1faebd25959b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc9e829027d81b1a767b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb77cff3ee85d97f7f871;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h930ab28b9fdc3e37259e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf70d4c64794a4685c9f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf6600538ae59d7990b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a95a02ec4f2e3695382b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12220991ca0dff01a611d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b41dbf52b150d7f5fbb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15821c00ba733e973ceeb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h181e315271de62e7c3442;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h172794c82533eafba00b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1359f7f9263a3d38b4001;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21030d8ede977e5914cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9027d4dfcaa811cf94f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18d0dfd6dc3a6696e891e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17b593f902b12ed0602c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5274787ed36e4d93feea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c188650795db36866afb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c6acf41e79dfe5249f6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186a739afd8c6d982f38;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h183d83838ca060ba6147b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1da4850e91b2eca904cf5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15cabea51b3294c44e307;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h158274cd0f65b9f77bf6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he49d97f184d856a16674;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h141ffb70d175fc78824ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9997c681e3916ca3314b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b70a3c29e70e8bbe481e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea0cad77d5693995def4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1853085d3bc8cf1c03021;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7b84561ae4df590d762d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15fd57eabf26100f0a2a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h184a17beb96fc4538a680;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e267a6a5f29fbfca7c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c54dcf556caa31e3e8e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a9dd8dad1daf5a1a7f54;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ce94a70ac0e611b9e57;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb2b4c756f93a8d0aaa8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbbd46454dfe17f835b44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h71f7093c29f75a0d51a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h155ef7fc55026176e7db2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c739d3cfe36fbaefe040;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119d11d0ed322e59ad79b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e23c796f9c43ec793c2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15456d1ab3f575666bd83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e235e66d1db4187d8c3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c33bbfc70a3b90d5c8e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h154b8613eab7dc574fde4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6d8892bac77b0b401d44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127e8051afe427ee90a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc7ea65251e354d6a2cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hedb6b543a243664dbab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1234cae442f5064617272;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d900e9d70991447e543;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h744aa4fc1a8653845ed7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7159fa03d0033d7ae36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd77e1ebac40555f3561a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d4d49cf09f16d7f880e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c41f7cfa615e37148c16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1208f39f12109670219da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c7058dd94818ef0ed849;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb785ac73f30b5b9e1315;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f06342ad3da47f6af0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h951ee036809a23f1dd65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12081703be588d7ea658;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9cf008e672b431281378;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19165441fbb39a4aa7d9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1880fa0ebbab52879c654;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a09e4f7e97b11b71abdb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b85dedb02757f8ddfd1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f64457672afc890e9db1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8cdad52ec33bdffbe0a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3c02e12c5e64330001ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bd6c8e79cd47633f7df2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf2c3b5dce608970083e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h64255d2cc7d589f6246e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19d51b0480dbc92621e08;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5852679d264f9b0da67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h49eec7945b034c543da1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0e32879e4534eb603c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11135fcfdea384fd9ee15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3c94f1b4b98a1a2be09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2e831aa7fc160296285;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h450c4a13833bf7574b49;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h383dada3f28787cb0291;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8be54a5ed7c6477e63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ae7c614e723fde75a23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'habb10ac7d3672b888010;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e4eb4924ca806fa252a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h106cdc0bb618d6539c347;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcc60e020921625be3508;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h99ac1c46d697c9b053ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1540af9a2bf1607ec652f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e99f41c87b03263ff61;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb887e54ae82b1a9c2e6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bed960539efa5d9d23d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h191048aeb47b527b9e1ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1332e988ef09031f787e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb99d37ddff4b89c19724;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178ffc2cc29285331f422;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e157a8e0681a8d20b643;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h334115bbe994ebfc04e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aa10db0b13e38a8d128c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13877afae3281b9a73c6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21c76141e5e6486415d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13e352511f23c2d7b8b43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbcc88e3cd28f538526be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf8a813893aca94967e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd6263a388f3cdbe1f468;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7967a429a52011bdbcd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hca85cd189f611cb636ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d2a3eeeb84fd2865bb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3080eef7e531072878d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h157216bb7d5c845e53c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0b224428dee42ed7d6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heb6ab5676f522eec0cbf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hee424da55d578eef692c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd9f7feb94057bfb292;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef541be6ffc22960d47;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94fc37ab7cb7855dfc33;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d722adfa58599158a0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d7546588a0b02f32dd0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7bcea3917c94134d18a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7095633faaabc851206;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h184dcad665b81f2356953;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he39cf2a0908c3c376472;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15cd92e12fa2218bfa596;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e37fa080147e87d3a23c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1e002d1084672c8d119;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb6c1c278fce141cdfc49;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2c90405ca303719b7af6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17121a50a39040949e5a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1401e87f7ef9c670be585;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd2c309035e7d040bb736;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdaeeb5858026e511309;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h134e99fce30b06f22a193;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12b61b505b212aafcfb3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h79b1fde4074d31395da5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h80bee2d019cd55fa6d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b7f045db6beedb908c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h45d2c6b99e2987cf3dab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h167aba5ad827fb046baba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8303f5c28b02fd2b42e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1221e5ea4c1e6605ccdec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h113831167e76d1fee8378;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b1364db92977d7f4943f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12591bd637d4ba343bc7b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ec139d357c6980ad46d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15124ebd3e2ea6de3f10b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h154fea7b59e0ba361504d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19225bb1c5ee4ef86be7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d0acc209612bc0212ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c071cbbb9a90ceaf8973;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b14d2dcdcec231aaceb4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af13e680495da4f4dd9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1052495cb67e18a11810b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e3a8f2693ccf65eb0b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d17f5fe8ec5f24c451a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b97ec08485aa87d052bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a4b70e8a27aef11bcdb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10126ed73e0403e9ba86c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hefa7a5add43708a6f846;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19bd951ed4610953c335b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h111861480ead847842fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf40224eb26d06c3b9fb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e0c0c20d0b8dd34a249;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1da567ee666c9a6e8030a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc76e33b06825d39fb175;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h59b396defa68a8f14601;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he7993e63f720b1804637;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eabe0c58c77fe4d2b77c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf4d66889b366b11129a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd18cd3327d83b81d1ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfefba1249fea5ac13079;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a559516f457fba36359;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8db1eaa9fb4e4ed4940;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a68529a7d280e252326a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b055b00dd2c71d7e121;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he4ef882fc80fffc041d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd987be1f51e821fcb325;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c415560e576ab8f4a481;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf746105f59ddf728230;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11394929fb3b84e5822ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c08ca1a6f5a208ef53dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf28ac96c669a7d0a59a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb24f7bb2300d849954bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51473037b6221eb9a1e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b793650566b6fcd47b5f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h161e3dd40349a223a93a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b78304e2cdd783e417d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h24da97edf14ed5362560;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h769447c8ef8fe7c8de4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca619c56b107ceb92980;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6a8fbec7741348e3552;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h165896222da8fea63188;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cd73ade7829324ae2c99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf5428c846cb1a6a354d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11db8a1d5d7d62f85e0bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16af46e939a85bda69e59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1663c5bcb43a707d7472c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd76a5d8d1b09bb8d71cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e44d7fd75fab59946b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f4fa7a122d4112f09f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ec8fccb9f816651f6752;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f446adcee3ab683e219d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c0076194c3b681db516;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb2c9dd752001b05d1ebd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9739b3bc9d381ea7ec72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h330f1c0172fab6b116a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a09223414bd7e92755e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h84dc3977c39b9bf043aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7f88591cca48df63fa2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b7e486fa39cc06fce99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1da81a9ee4a3a2e5aed63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa52d9abba99310bf046;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1715f55502d3a99272b23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fdf93269117eb1184cee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h324df041a8a7c0ecca7e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc1571be82d45dc4a687c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bea022728569160f1689;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cb8a58f51ba8179c62db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d8eef7257c1b4eda112;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h540481662d6ef4097f1b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8ecf1136bfbcf21c846;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52e28c911c0e932638b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18d91993305a2f968f27d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4869e3934864e7c44e1f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18add2e2a3bba09a5d083;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcc2262d97f09d2cee888;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af8739a84ec9785f7d6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1325faaf77dd49b7f29c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h164d75c19a5daf5d94a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h153048dacf0e9394fb6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c11b0e21a3aac4036ec7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ec63bb4ada59067c68b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115445a0b017447c9043b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ecc63b102ba1fb75bfc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d74c612dea905fbc225;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h74c6d99aeab48cfda38f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12b3d56d953b7828d885c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h181525ead3c8f7b9334e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b912f0e67641f668fea9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h164bee4eb8ac65904e1cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4645d68e7112a5a337e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c42f0c6ae1dcef53aa1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f21afc74efd1b3eab882;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h176d4d85077e8940042df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ff9d62cb42d0f47b3360;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18a12877f801c4c8bb8ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe0a5eae68a49a101627;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h193d96f4b6605f899dfb9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10ead158929e04bff971e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1973c313e5f5e82384b2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14a04d8e10aa9facf26a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6621b99f92e9a35284a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d761d2ca19c835a94bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ac50522a0a1d61704ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h870f12a0940ebf2220ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h198be502719f56a4778fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1176c1e4815b7d19d1318;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18f4c36c4b3053017c81e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1919aab0341f0a484918d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4238e12662c8b870a7e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f900f3fd584b49c0af99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h190c2e9d4e6f8d6ac2907;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19745fdb2b279f0c3642d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1da1e1da2f73f12c986b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aa65dcd4e8fb4f048aa6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42739e52392c33119d91;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb143d7454f1073f35be1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68bd538c755173ab438c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h155abcbf40ead7ca6e66c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5d04ebcf27d08144d12;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe38958c2497b0df0e52;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h126863593a2a46dc04fc0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12035865c46612d88bc80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdb2ce6836065cb15d83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b33829923d43857f4c12;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h525bc5936a4697d0db12;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10b23b93ab21af9e40f5d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1992d6cd5b020e3eb1e30;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dc7580746991f3ee1d9f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f039248cc664ea807277;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e2286c661f3253129bc0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h99cd6c229b4632fba4c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2f8a99f51f130ef21af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5f6db0a248cc7e99e57;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10b63c355b183b2474b90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11de8586551128b964f0c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha31f06f5c6cfb91c25c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcd1b8b6b77855ff009d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13aab1a6cb0fc4c1649df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1872a79440994aa425542;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b96bc463cf38afe976a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44f5ba199b6ff89530e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e6ca9649582a0c30389;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfa4e9a38abe82d89ab7f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18f9e8b6e931ebadbed01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf64c0653e4ce8b687f07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14f5ef7a384f12e75872e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h128256d3e518671a47d37;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h502f12d0ece4bdb2ff99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11da719fe8e9c93203cfa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15999e6ade9bd92c9662;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a529ba0be79ef33e886;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9f8ed59c908cb7ed14e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcc3c6edd2289e51a625f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda32e9f8d0caf304c4d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba2564f56012ca581ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h23cbda572b8b407f6299;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5aed780cbd942301ff82;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef467e6c2028d83afb33;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdad4cec31421c30ae595;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h285b7bad798ea41611d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b5f28f2f3508c8a9b54;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h128fc300b56a8b1aa9285;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h36e9c1fa197ccba15cdd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8a8a4dae7c44fa1b260;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h125ba13d893fec5e63c41;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e355ea7617580ebb663f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8317b44bc7e15ab19ab5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h199cba6d4bdea9d81060d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1711dc93e60840fafbcdb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c61f88fd84f422dd0b6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h107755caf33d28e97bd1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb08601574fe2023d1b0b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h90ce3827bb15716e550;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h126ca358c0f345c35f664;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0e6a50e9a4557d6431e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14e4b97e98c62bd698cb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd5c025ae9ea2acf9be14;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h167f7a531a1af0f2a7f8d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b9537bc51d010a2a37fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h70fedd92e476460c3042;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16675d52e87919c645c6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5200fd002438f7bfcab6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10566edc968eb63c18655;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1650086cf2702cafd7a42;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105a10c3e03a0713a46da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15375cd54fd44d0e2d033;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hafddfed564887d278575;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eecc39a88d8a874bc49b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b4efb7f8efdc9585367;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a8d59a30a52de8e1b549;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h35632ac0061e058c5599;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2328799d68a683851626;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc89f9876e2a4c34b3888;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he22ccca036e01dcc6daa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c8fc3a19278f90f9b58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1921b9968f5edca398c07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'had6d428d3d398424628e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1170bf0a0bd70ec63aca2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6143141ee10d742dcdf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ae197ef3bc58fbe98af7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h70afef6b702e84dec40;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123c760fad89774efa566;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f6d3d45b2cb94699aac2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5941f4dcf469459cc1ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b8ab515df9480ed2ecd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ff597c48f8650beb9d30;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h431c2e38ee98f3dccd9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e813cbdfc96c81a012f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h281e7217f019cf88a36a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e27351304a14c200cf9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11924e5e9022bcfd57179;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf21473de303d9d331d5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c1f9a0d58ffc9e8ff5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb73ca03d7835d2b51a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18cd49dc0cfb2ae550bc5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h627907d4319bc2886803;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1edbdac5c150b9cc4a4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1652a3987ba55ca356f06;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h588c04b9ada15cbbd022;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h154802ec723ef67f29291;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h139568d4c3dfd36ebf682;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h193c5972bead8aeea3b68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4432a9b1a17d77c64cf9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c755958dd4ad0901b84;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17368c3543cbfc07f731a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f74be503ae7dd873fc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1597cad10d546d4f80a34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5e6148df20bfeaab02e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h82dab195ea02ee52ab31;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9341d6567f69cfda2aca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f8d29831f564c7a5996;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b4b3f5a748c33240083;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fd2b40f7756f04cc8f29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c6cb67f4bfe6dd00493b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f8788f83a16c322901b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h145e5e9a427038feae7ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1202ac4e06b8d069f4e6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9b2aec1f64766994014d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc1deda27c5bab9444683;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h575018f1a1b90419e2bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h37f55e475d7f38306062;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92bb148b6c1de4dab8c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6fb0ef40e73b0b01545f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e8f5cd321442b2f6105;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h72ab80f9c7b551e7b3cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1339dc4cdd8e3e3fb2e3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1065d475daf3050f28d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc0155eb78d6f2f32ec09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2b18da0f0965aa686261;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cc1aa1e46477241ea24b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc93ae59f4f0a239b36c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196c20e1273c94bc7b97e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115a72e7111ff70739525;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd47fe108e89fd02d733e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14964590b2b748720522f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h65ccff25752f5d468370;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11eb771fa3f51f89c7539;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6ebaa75b33d9f39092;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1867a2d52eb70b3546b6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140f39fc6c8b0f1fc3a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'had77dd93fc7586b3a91c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h109d8e35b0b1a1b940070;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7e02ef1e3de1210c23b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115036d9a64443b6fce2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f845d7bf543357e10cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9197085f5126c3c07d97;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd17949440a6c28c04943;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8a64cacb1a313d5e7bc8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h677fff42b7757c04f46f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19704917e2975e003aa1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1010ff9f1559ff60c265f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd4e3a14330ad3bd3545c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1616c81c49a2bdb54b4f1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2426f8bab8ccae615b1b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc520e5615cd76b49371e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d48af97973eff0d76df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1436e75e86f0235f54b5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c535ac5d8fdb975700d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bba1724bc1bb3188f3a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1613b7115bf5fa8d72b03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c042c8a0932852eacfb9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h90fce9ae30b7a67ef910;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h61238ee2d12f22e90acb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f14f35f6927542362e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e59e53a36fa76f0322c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95465bdadc58ec3af3ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c6e08adc28f566cc1ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9bfb5d623e17ef3e9f96;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c3e578cb901aa4534ca3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf3448cde2d172cbf1213;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1daec0250d9f7028e4da5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4ea3be88a299226cd3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f9b4c9261bb73b09bc1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18aa1962c4afe63e557c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h197dfef4d84909723aacc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9f1f9c8152790a46f2d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8ee1b2fa718dfc4ee50;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db2a4093dbe65e1002d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4012ddb4621d0854b0aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bee56d917cbd10352e90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178fbdcc3e33136c9179d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f342bf59bef41f4df23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c1686799c8f21a6a858;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f273145ffd70d1bfcfac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda9e90b40773d488e91d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3d2703b3586bb0302e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1fc8ca604fbe1b85df6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1deff7af9597bd17e4fc5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3c89f8e1ff9bcb753698;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d9e9135c4a9fb266cbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60fb351a23c3fdd0fce4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e11d76e8487cf268683;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba5940538c118f172e59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha444c63fa6d8a31b31a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186900c75a02dbde1f2f1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b1e5c8e7faa8f7bff63a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11badf539eb461700a0a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h287493f6bf2769516bbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15cb3f98c018255df4249;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1964c872a2e0db6bff908;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h96c4433d7fb87a0a1e50;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e32cc4f5c60edd08f62a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he299e120809d3b2ad115;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h277940ca8b53b28905d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f1e95c8ed6180b7ba75e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19219223ba3bf4739ebb8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h193cf8eaa7b63d4166ceb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ec7427b90a0d9450e7e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11512ccf4a1befb6ce802;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f6c1e9d06dec73f35518;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc9370b7f587e4691dc7f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1108f5de3b226e2bfac4c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f0b100231b34167589be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h144d47a836cf7ffdec6e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7256cdd98a05d2ab6742;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae06a5b7dea8cda4baf7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h75835692ebdc912d53f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ea0a38b0d3fb3e4a581;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h84edc49073ae0288343f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb815b683ab1246ba72a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1836c20cb28eb5ed63c2a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h533021efcd963cdc6c79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hffbf23bbdf2555c1976a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c31f4ad262b2c339f5d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd4263cd987aa42d33fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7dd8397d26240fa0a36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a397ff3b96025ec254d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c4cf8a6f0138ed76aa1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcd6bf8ad9dfaa96321d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he40770eabfe456d686a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h70c680e1b146432616bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde94bae99d523dab0994;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h990fa86d70e148bac72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14bb9e00ec90f933478c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db68c89e2053cf612aca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10823e74492bd5dd493c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h110d3767b20807b37c751;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd381eabecad4d95ee52;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1357862f1c1a9c87de5c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h96da90e901eebde9688f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19919e0c25a9d3af6b71c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8f3c097a56001aedc358;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d4d47e8f40471873996;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3632a01c1a4e74ccbfd6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19c864665e363021117a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6d3719e067f4d312f42a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'habc0aca795da1d38dc77;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4cf0d489c1b66e7712f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b1986f32be1de3eb9173;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c9c6aa116203d4d646b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce1a30eaba85d0bc9856;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h164eca2322d84d407943e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13f7c3af8190954617002;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha29f59480504b7aa86df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1866d4448b5344d131de6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9bc424a7b0c1aa3d307b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1247587efe765d1143f62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1877adfe19ac9b3203cc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1358ec0f8924a81bab13e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h131c85766a0d1910c7d9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5dc81f9542d9b3fb400;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d90f65d5dcdaf6ea4bf2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha270d13a671f522748f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ec9d8488b8b80713bc07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119b6227f84c6fe3153eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h176d52c068bc36daf49cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33103934b30d29c9e093;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h74fc250922e485f0ff18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd8491b3d8d4b5a98916;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h758f7a6ba0327ca03a66;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d8bb4f8d899d35a6722;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19fb14624f07e1125f850;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha18608c907f594aa006;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2aa81f2cfdde87dd5fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h112925a255823e1113fb3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cbf2fcd8a826dcb0d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbc97921f2c70fef990ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h72c870c8d488bf05153e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h750f8b813a7828888e07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb4cf40c63314d4f40fe7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17a3ed84a55ab39aa12ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h23aa78f0ac514547937d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e454dfde4de39c0a0042;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19c53c35d4229b655a85f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11fc9c9d950621c2b7bf5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ab9b9d84177ae9ccd96;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h587fac353c688d7dc604;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb928585ff77aad44a30d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d69b9c6cbd94e776a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de5e2eee74dce86a1824;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ddf801beb4f01cbc804;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5fa1ef470836dfe7d06b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h954b3b24bee3eb97312d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4344991d66ad73ffe58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13e2e18e3dc9768e3123d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b2ef89a97296b56cabc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b2dd36745118534a92d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf08d94ac58af61ba6cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h152d49d3cceae2342b761;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151dd234b6f76df7f83e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h149063f089bf2ba167bb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2e2d8f9446e0b1b532b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14731911a9b8632f13c8e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4773e3ed7609c709a998;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d392a02a9ea27d391e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hefc0280f59985da640a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151f56f31747323d7bbac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104d95b26497e6f246957;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2225faf3d3ccfcc55f4c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1291dfc08493f7ce8aa6b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1afd833cdcc0a87ae24b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb08f537793d97f58aca1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h109bb634cf912a9eb6176;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h55d67ac33d0712edafd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac70abcefcc979ee0db9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6a3e32d37515b375052c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h117cf27ab841ad0842a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6ebeebfe535ef5d9c10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h25c3e6309cc0d9d36405;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ac4fd6a0549851a8ca1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha27872cef9f16b09af30;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h688a66d38b566d00d25b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f358bd16a1253b900afc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0f203d70c2ffd5c2eee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115737a93d9e45aeab0c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192a3f066b694ae1f23ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb723e4657498ac2544b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h75c674f65035896d06fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he102ffc644767984dbb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef573ec4eabfb5dee087;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18038f84970f44f8c38cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h98f593f23a86d662cb67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2338d34de1117276291f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a308a177d1816f50b85a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8f0de29ea2a678a9fde;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec523629f3b47aca7f10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h73ab043b63fd33fe100c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e55b28407b2da2d2766;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe5956996f2af3da50bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10fe2adfeef0872a8c084;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf328c46647f3ac01b98;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h169bcd08e39b7f8f72f29;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h147fdb025662cd9a4b02f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10ae33772f3a28e2f7943;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11977f32251c851d30e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h735329c0befc29a19ad7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42f857971a38516f4b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he79080e630d698b9e1f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12aa5474736f2c1f90342;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a6d06c3d35d7b5fe920;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfae9159c0efe86af61b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hee7c2c3abec930a3ff2f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a03093312da711d524c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab4aa092d27da774e65b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h69415ae1fda7f4161128;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19711480a9d13d69585a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e64b2f433b3902153e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ae9cfbe339a17510c17d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h138d1a062aed540725e58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed5aae9670dfebdf28eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16db05d6a6855f5ff8898;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4cae13b1df83b2e220c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e5f7432d830cf68044ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c30f9969b99e6681b5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5d66169e6998fb70c13e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15688ce9b611b45855683;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18085ddd9ae518c90e1fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f21a503d864b57778b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3911779af2487b74250;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1753ecf13b55b29a10be7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h49bac625393a49a36dbf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e34dbd16f74de57d86e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6a55b4837ec0aff0daf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cc2393fbcfa0004b5442;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1468af435d04e03810f3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b135b86001a9fbb1622;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f65a23b1aa74f68307e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19c0bbd296e1afcd4406e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha57b386ebefacdf94203;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d823e766ce0b076d5a4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15dc275b098ec041cb81d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5cab3762c9b4efad371;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ed3f86bd985757c818cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be53d166ab6537c6eaaa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a3c8092d0774ef177c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9df8803f06dbe9ebd141;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c4d738ea17c9a890ee58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd47ac79f5fd03965e6d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3434bd7946ee9807afc5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha471fbfaa77804b9a26a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha04157dd50dd3eee39cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3ee4515a01059dfe987;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa523933a436e251a48c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c8d7693c8398b219469;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11991fb4a5f0a89ed94d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1338fef5095c3ce5c451c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he14c0e9cacf9fe5af44c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h108a183f28f2716aa6285;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3f8456493d180ea5976;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h74aa7211cf88cfbb9949;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd7fc1a99453acd800f6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed63d9087404056ad58c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5436fff16439a239d71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1217e6c42d1e004457d63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ca6a823989d24a2edb7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c004e25818a133860a86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea00b9dc6d6dcd56eca2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e444fdcb6a76be1c26d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2a0e0e5c943d3b956e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h137fcace57acbd49b08d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92b05c25cc8c91df47e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19baebf4fed3fd6b14faa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf1a10c4a16bc85b9f50;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha25643be29b7269930bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf0af94ba9517042b0fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119c36f353e52d935f2cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ad6c83c3d5511d1e98f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19121d0e50c11e493a921;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c048304955518c16d128;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb601e2ad93baac0b9d4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ddce500369b8836d915;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f7771a34eaa1f81eed3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18d2fd9b6dc12742b180e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124cb6f382542e054a4bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c97b88f97fb593b707a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3401fc15ae8bbabe65ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c19a687c1d49dbae0a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcebe62b7c5255da67845;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5734806be6aa2c825f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b5100169b9d4a6d361d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc275a0a72988eb813d22;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11985ed7f78918cf5be6c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19c5b1619834e5cb688de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31b9373181b4b67efac7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c61b2163dc9829442ff3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h193df768b638a25afadd7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ad5eafb540d75e6f855;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb714b727701445b85914;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf0b43307db8d95fd16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1905d75ca4d7068f37ec2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13e9ca1c7669ecdb6075b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db3c0f637ebf8b112f23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d4c98958ea4c3b203b3c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b7eba5476bc78e5e148e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7e561bd67320d06ad4eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14557e5700dd6b98373ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0357deb2d5813fa846d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1033978e48fa2d5194362;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb6193695c78d2f22ee89;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc0a9e55f472d9c2879a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb41536b66f14c3573b7b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ab02dc59235865a6e90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6336688154708c95c4eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c8959b4f182a5eaf00c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14057026917e54e2b5662;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9c29c33a08620d1503c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28015da300e81bb0081c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hadef1cac22c548020e01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h275ff952a5c091eacc26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150c6edcd50165192b889;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4f5e4e91d15969d77c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hafe428e489746642fbed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h50195695aa85b17364a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9aebbcc4fa9c2c1ef70c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1071396e341635b8fd907;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2cd8aba27b3fe56449c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h112d6f9994f7590a55abc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8749f5c9e43f108203a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e18d507cceb7abd6f011;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf492f50628ab064de5cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10fd8ff2c55442e173e7f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf81cd2b795a316ba8d01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19eefb17f615e564113;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11b45e88b5acc33a04fd1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b4d11fe6026b8a8961a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10606ec0cb02c66c3d35f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53c478057c28f6185578;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ba915b0fcb0b2f764cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f0fb9a0e55e5c72d0215;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h61714c0a0cc641f652e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d81b0915f26f77cb601;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5d4bec3c5716ddbcef3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f766571b4b4a28b1837;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b5bfeed70ffcc513ca42;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h194592a64ddfb97fa7114;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h447306a070d9169e5144;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c07ca1bc29b3bf0236a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18bb90f4bf4e2964d9134;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e3eed726a879479d786;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e057f12a862e0bb9d6ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c0915e84ed0eb1ce7a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9ca3690a341611eb502;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9dd8af4df859845080e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33a1aa56d3a49a39d6c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1697db623de31785f9f91;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ceedb926feafa9ba054;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha254b990d1d83d34cf64;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h213934c2527dea88a580;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1270db9a9f43c0d55ae1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9600f4fb5bf2af04650;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ab265a3ccf6b07ff011b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6fae45c17a32f6df73ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18f8b4d397c14fedb421b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heaefb33c8926cc35546f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e19bdf4bdd757b12f14e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h378790e39cd1dfb2b08c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18f1d12731f3b8c6160b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h149afcdf06ef478635d90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2cafdbd704720e5cf98;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h64240c0e6bb8e698ea72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fcf89761f78ebdd1ae6b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14e22400a378e494d2d1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f2829a98a5a49e215f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h154c80d2faa7f36d6b659;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9cfaa96d551a30c045ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf8a6d56a88e015b4a195;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c24a1457e946960c5675;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bb526c49890bf29f6ae9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a76cfae24453d19c4fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f21a2a682754e075696;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9e455227d7e7f50eddb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c2810102a699947d212;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2897d8a706a27b26f89;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f51119bef7a21633dec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h753681f9460b492f2a45;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83bed479fc73c4395f48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h183a37dd6cc1841badb37;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4dd490b6d74a5063b495;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1201fd4d62e0888a0e01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12409f1c0fd626302603d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e5081718037cd4403436;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13fec4de5c4730a457d79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he34ba34fafa4c40d0c15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc7777f47473027cfe0b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8db83cd1a6db712fbd8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16dde9ae2a6372b44c83b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1357cb1b4b30b4e5298f1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14f6dd32bdbff4050a8c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf3a1e6321eb939eafa01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h967ce4b7c614c4abbd6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1600d22dd4ff94ccc2d42;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h75b0260d521fac25e78e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d356a64bfbd513d8fb5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h341a973459f22c17c567;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16e3ef65d604ecae0a1dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11bf07cae56fdee2016ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7147bfee31d2448aff6b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1981889de2d1157770567;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fbafccd83df44ee5f8e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dc907154bc152c3bc118;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135d7aae871220090f88b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6e3d2c5102d39723f1da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1750263d7c8ebe23e913d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbaf0f880fe1e9c68490a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9c3a172745e90541d91b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ec3daf4077ede9c7679;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105bd7b23c82833d83818;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14286a6e7b63f198bf796;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1079040a9b22337f87194;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd317b220587b3f6f9ac1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he600e6a786c7472ab040;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d8199e2448f1bab26a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c04a68a3ae6eb9e0819;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8bc6c3c724b515c9f960;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e5813d82a4f5f93bb6c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7569a2af946cb6337ed4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c1c40a1311daf130652a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1201f24c05eba1279b0d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f1202ad0c89485ebda3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0d233cfc1fd2d2e393;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h111891c77592b3c5428ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f4ce5f73e74d36bf0685;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb11dfb2618ab4fb6b0c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1c86e0f2b48309d23e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa0c7bc44c805da066d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fa48539b97b59443e04a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9608ae1bdc41a8c674fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12aa590c97f946c0db727;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7133f38752577f5ab770;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha1d801afc3c133721b20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8b1c7531e7d97cd15427;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h687e4778caeea6f71e49;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44987bd7b3a74d74f3ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2f919870750f64dd522;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h110143d320607651d98f1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc337eedf0c1a079bb378;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h113ea1b7e7a49a70c2a2a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e5c5825b6f872360ffb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19eaf377a3a7fa19c7dc7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17539213c37d637d74875;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h69b7eb29d46ec36c1bef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d170786fc4a8e1e3d8a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h348d9fc57b731cb7825f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h117d51e396af84ef62f10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h24d19e74a276cbacafa9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fa9eb43c77933b2328;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d866414fc7b93bc81b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb224d855e277c7522c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143eeb6a47ee8b7cc6f8b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h81d3343c25a115370310;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d35153dc4b9b66aab36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ecac50dbfef3400febd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b1f497acc21e9a6aef0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21bd01bf5e2650f5bf5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d57029c4d33ae55cfba5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb55060a6637a65ca3a1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d2edd5a47390040b766a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4bcd811d851a9519089;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb8677a6f412938fe6beb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf39d409109f560d2e4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aa0ee42b25fbb22ba5b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ead478470710e7db3e2;
        #1
        $finish();
    end
endmodule
