module testbench();
    reg [25:0] src0;
    reg [25:0] src1;
    reg [25:0] src2;
    reg [25:0] src3;
    reg [25:0] src4;
    reg [25:0] src5;
    reg [25:0] src6;
    reg [25:0] src7;
    reg [25:0] src8;
    reg [25:0] src9;
    reg [25:0] src10;
    reg [25:0] src11;
    reg [25:0] src12;
    reg [25:0] src13;
    reg [25:0] src14;
    reg [25:0] src15;
    reg [25:0] src16;
    reg [25:0] src17;
    reg [25:0] src18;
    reg [25:0] src19;
    reg [25:0] src20;
    reg [25:0] src21;
    reg [25:0] src22;
    reg [25:0] src23;
    reg [25:0] src24;
    reg [25:0] src25;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [30:0] srcsum;
    wire [30:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h603b5a24b26920782b64ab77afac7e4f43771f57e33c8e25c6b013f507bacad61fc5ae5d7b0766f75a293fe5a06723e89aec18b219f97d3c94c9a44655f3e59b4af1ca70b4e02b50241f4c21438087f323b53432b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd48c3ca75071954129b87ca0d728983ea979db807d4663fec871896c838b2c1b96863be623266a39da090894eaf4c8d4af7d708a867f41cc40fe77882b5129bf66de35713450cc9e65605a632e32f14fdc569c9f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f063bacfc8cbf0a5f997d963f1377c38c8f01011e68d86e9e1dfb851d3360a0c7a847d97afffac6fa1acb58aeefd2f3f5d759508fb818fc442818cc5ba1f303e4cea74fd16990cd90e1aae48786cdff69b5aa76a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf440d2f9fda0f0183799376bd3ce5065742b4a29c4c8d2b1c757a75269d7899aecc1daa83160f81fc4bbcc16703936f642d18d1a4d05dc65c0736f730c73a4d160c7e5befaa395924f0dfc31672758cd288db0556;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf625bfe222ce2e55f919f069cece3fbdef9027a00e76be09f57a9aef26fe1c67a07475ce21f2aa4135bd1faa25895f3445dc01a8d8a2b85ae25e5d9ef3e77e070ee73fc9d5ca2221627dff5c00228d4764c40c779;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ca4b9a9b56b3d23764f42fe7f2e7a9e182955013a0f05d1566bac34ce937e5977a14e7b12107ce7ff8096cbc3cec2b04f7dcd4da38d387fe73b87e930c08a728c8fa2755582103f77ed4f531d585923e864e73e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec158321c10650a09d0061735401f5ba081f44303c5163d51c6431c08b37e02ff41e0512419db098b2fdd9f4944bd36a60534547608cee9f83c842d5689cf2719013a7053025acad105e5b41afc9d1adf18890de3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcabc393c7b898f2f9e5df7edf4da9c7acc478115e6a9dfa38e2bacd663a6f1b145aa52e0088078b35038cd0c83818f4a0147a4ef4a31a624ad25be45fd014524dd1a58784590296d4261aee2009fc806146e5e893;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37a3bf91ac26a95e436721a4a70ffa395b09e981245ea8d16d945f9c90d27cafb0fba595e106e650d723fe17e0a716a5c114e66b30b3e0a3a56a6b50df3af936231ca2faaca623ac48bf3afa628b7c2c10106abd3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53f82e54622b7e122c4921f735d6d95c659786f683485a99464a91982b5c16ca0780878cdd38d29b97e246ac57e358aefdf6579d0aa03533159338617c2ddff8667838a3a2e13d75eae3ba88dcdd32a82d2b271da;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b923ffd98a0093b6af080aca42200c233339f6e3ba7ce5e7d211a5246f96ea5118f1e60377c9997e14f0d6c368902d8e8615d8b88103451c9f4969eb3908f18593fb0a399a49e9b9f69f938480e620ea968d3ffc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd732d71eb6b8d909608789ec83d6f96ea76968e7b2f3040a4c60b0cc6c8ab6eb0e71a3e3b766b251a286262d85cf1cf8673eb31d09fafc3563de068ddf6740faa60f4fdd2d17bcf5457e4112f9800cf172aa959c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c113b7f600e77610f06a56b69135f5ffa474ba0bf2cb3c88cfad000413b1a585050a16d027d7673b748f6d356beb1cff4b52cc5d884ef95c9ea2e97942addd70e3db40e04e42fa9db664510fe299b6664abedeed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc2875ba6012de887bfdb6045d3f45edb6cf75c3b55652dff076abd39766e50a8c8f564841b5c573e972194b8eaf1e0d7d171a10f7f67700aa50ca6ccdb9ef1db88aa107f6fb2958650329fba251571eb4bb53dc6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99ac0ae97c5b659207a175a4d2d5a12fba566b8b777214cb433f3198238003aec29f8bb523fd092a1058f90918b0cd5eb35b83274d0eda7696c9e600c5f9d816adf7ce94bb79b2e0cf4e90d911f103c52efe92fd8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46338fdf21b63391e897bac1c44c3324a62de006e310d3cd943d049506fe95e5775073d596715ba107d1984529dc518c7b942eab56d4acd43926bf13dd1ce9229e980737e0c7cc7a5c90324c21d1cb6281dae6653;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e228ffa9e3733950633e1ad441b5ca28a999714460729f72796dbbcc4473ef3d16ef42bddf3bd71737d8908f324139b640c5a52431cbd6a3cfcbc0b783d94bf40a1762f3a53d780d44b387bb8cee4a088bc7d3c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3fb411472231ff8b6ede3eafe68b61e43184ba5e939f8b95803c397e4e6bc6fe9a3879d4843a74ecb3718be2f75bae2df351ca71761e1b84f77aeccce08b75caef23c26e835f12d5dfc6e7204fccf933d24928331;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4b94bde8c263dc97ddb5f1dcfffc9e0ca261b1f3ff4e488298b8fbfe3f01e96b098bd804e1838540e722aaf271cecf4b03edb4decd4de4e3c06a0578d926991ded3a1a710a76192167f703d210d1abc6e1e076de1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4600f43b80420d7a877050e42cacf3e556de8d3778f092ec22c8d7f7eab988971b90e8ddc33d65107200c62368138000d170491bebdcd81bc40aac6ef362a967ae16c5999c2a8105a5191df66287a2027633540b9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc837ce542fdf71455858296ce5be9d14aeeea8794d48053e69027f9186c6a3beca88b83183207540d6f374888933ced3fd8a152a69b5af0985fe68a3f13ed02d30b1e2531adfa6538735da7edb4e1e6768b2a84bb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h121ff616757d2ae483f0c8d868b0a00c480dc1653e959986068102e220bf855687ebd55eefe09b8b97d9c33d879cf4a646390f5a828491a7151f3e65b0fa73fd9fab25f06161e10c5bd91eaf7d30978cc866a37f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99fccf13afdc952972e47bdbe2eb339d9ac8ad146d2acde6132d7929bd663fd0bec22f7260c38bbfb31586e2cbcded1d1c21683801001f5a9a5e4767ef987b19987bd32299b16de5fed6e0b2e00ddff70935f494d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2dd72c703ddf211a42d6aa576a83c8cfd46844cefc770ff9f229369b84da490406853eae549bc05025a22933ffe50f200f482249a1c99328a4526b6b67f864f9cea71de7cab6c22e6fef99dd9480a879940db67b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h30c5cae8371871455123a0baa005b306b69d8bd5b1b9cf185b98a1ed467005aad151c688ba901ce062c7e198fb334fe4ea80fe31918d537d87236f734b28ab4277982507d448aa1d1b7eab445a350594cb7719e0d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf51d4fe791511772333e251b389d82131cf94f388e3abf02638a076d0ddd4b93db8fc75ce0a05c0d6605fcf1d5280bb8d0d34751fdd4d6c55042b992cc32f72cd8e59f50c5e0acbc32f6213df077d640d6fd217d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f9bdece59a2ac7eda4ccc547f025e13eb6b7ab2837e1889877508e70893ce5d61160774cf9e67ba2c4bdc322251ae123ce80c83345d8ccb7f391c763d7898bb3077d7d0b6e7f24f3d0211dcaf9f49c6d4eae3e3b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf4aba6e96c46bf7a924822fead7104f040ae166b0fdbdab896a4e63dbda85921c6417358d507682517b90ddbe68baf69175a1280554127e3332ed2118dda3023a8314bb9ffa2d0a2c691d24cc7cb797a8a2cac1d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa6a46f78c753a182c75212659edab375ccaac403d168ef2c8b634b963c799631c759248085579ef38fe181324f066c7868a7968259f908353256a2499999005bd6f240cb907258bbbb579c68d37b1fad64ee961;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41861b69112c64537f78ad6e3d74d7e75aafc0eaeb0f815d459577c40660bf67dc6e7aee5303059fd1af458f3d2f58a55faf2f773886af1f2f36ff671105f6241e9f31e5b9991d4358eb8222a2cb989377b409bba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a364d23697449125d9ae45c255d929566ea2226655751cac33f4d0e6902763e1a3877436b62d014860fa102b5eb14c67d2a2873899ae9eb43c753d472356e8a1b12d321a0f6432772ba2770ec9fe1f64cb9cb0f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h204d78b0df8bdb2ef419747c23f95aafbf846908c8bd56d450a44f8bddedb4d8536af993797c464262f5d85bcf47c34a30e4e989f1f28a9427c2b372ef0808cd348c522fd0934f315faeee767cf7975b57292f675;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7c1076e00c8317394f157f31ee0ced7064ca32d27ff39e9353218cd0c4a983e068598e9dde0f3fc1057db2d82296285de3e74737cd1a3a97126c57cf27d909d3480d5db292c9e43e582e2395f4edb54f682dfc1bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7ed28745f0bc4b01964654f6bad5f065c2fc7a0d676378c53010f3680bbb26c6e3e9360c27dd6ac719e436afb1876811392c9f4d4b0a92b4a7394d7b7136f8f232d32722cac5092c17a7e4632e565428f72bb44;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39b6e1aa5421e61ab6e7f089cef9ab49edcda366295398c12774e9465dbc141755dba84d8c6de208b00080e32468332b79e261d808ce2811ccdce5085fd8dac1e0349f61c9076ba4e66819c17718e1a14e1d49a9b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h141dd7f55cf7beefe500b272374ae8b35b278eb6c341d64d4fe69d4b9394d913532cb522a357b09e3fae4a530500b252824c7fc8f6cde26d7fdf153b4f7308bf22571a100362e2a31685696fafd5984dc8e076454;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda5966c4c2024b30e1d365feaee557877a27c607ebea4971dc6f618a31a29b58e8507b6f88f33ce36b1603c4fdef4cf21d27ab3a3881311d465a83411aee6cd5937c2d8fa4cf6aaac7dc09e6dfdc72f28e3ce48ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75fc502341872eca8a784bc2f72257e8fb05d850f2ccc71c8376e4813b675683bd06a3233556fb888ed3eb9e92092056e2aa411a7bacabc17fc676f869b1d1862d9db646b2d1a5443f132375dd6e12d471ea1b08;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf67eb0d44272940958e4e85c4826ddae39eb48325e7046ce5739b9541ad8ffae6c05386cab01f54ceb35aa0d6930421f46fe99164d81749a63b2feb07a4b1dff6d57ddcfda042bdaa830f684eead88d500d6627f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21674ad031fa925d6e246b1e5421067d0ab8701e4e5b5d072273085812798728bfbdb9eb33441ccbcae95757873b9ab996b116f31e0205206cc99883e90c89900cf4024ac2420ac93f34e14eb1cdf472b047a199c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha641704b06aea9bfc20a620955ff2a33579646fa18f4836f3964814f36fe5e5682e1a9a39b5df1341da8d469042bba5a9a52406364cf12136034f25366eb476132de788a15442024cf665b537d73893f3991fc9fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2da736b031ab4cbdafcc555341de15c2b11b3304581bc41b570be8c7f7c9c1efe9e7e77c45ed5a1707edf999938fa32fdae13ecde3df9996aebf6114bd5d830c9f157830e99a568265880d5aff7dda69f1bafe13c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha60131b6c71a6fc74393d0459570ab7560346f1d6b66e6790e8418d294694ef16c3c8061003111fdf0d657a1d39b707fd9f9177e029390aa95754213b909e42ba650e771bfe5f39d1c1641371c2948f5fafd5809a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c6058c3826acf0f038d8b0246e1dff93a141f8a0392861f6699cb551914151cfc06f6e88e54257322335c00b0dfac5105e71a0c1f9e3fee4f4b6cc0200a5a726fa347364dea66e9bdfcfb094ee25e9c6fdd77466;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67ecc4e6cb3b5d9b272ce0d910db752b475cecfc1c76feafe32c81e40ccba9642de228cf65616a5a486fc57b88379e89cc47168866b2b8f3ba05a1e1ae57718c3a893f6599f590ee51bb3d31e27d62c73bc304f00;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a45ff0560997bc54ed4fbe62a3afb93a6576f067a80d7ed85f3601bc857c3cfe9a37e8943f26d023a100671540c4f03ca1e0ea6994506e52a6d218a455c641d366bf67fdf1112d14de062aac09ef2106e2250ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90fa204a4d0aed21c7220830c615d89d7be34382d3b33c4e3cc5f631bbc41b7012a9651e8857fb75706234014dc70dfc95eda034ec39a3272d4ec55cb4ee5788c93bfb8cdd2f4b7748e85b6c49c877a10b7dea15b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ffa400140c8e9961ba414f5e1ed673d4542f1eebd99d4f14b1a631230190f327baccd7386d13a55e50869d168f21c7577623c661c03a9ced73ed423a741efad7c52353e95daf5cb73e186083b6aea8f3493a2e13;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3791373c3c6e324df33d23fd319fe0af632ad8cd49ea24de5fcd378da61c41196b9f6dbff09b94796cd87f79903544a24f9e01e7fd634acea0583405bc5b150eebdedfb27677c72b8b3bfccb41c2b7e016aeeed35;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b0c886d8f7772e89f6e3250346b3dfc17da27b8a7a45ad0cb8faa85159eca3a90b66f7b3c4d1196654f583dbd8f1804502b7990959aef73d4e322bd628eb0ffa0d04fe2f2338a5c6201177a3e24867070d2a4d46;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h759fcba41d02ce2668f18927dee71bd9c2f3dd8421a99463a94c08a6f487f10d5fc7bdcbd881b2bba1759e831bbec8a9042292af8446fe70d51c875508fb212b76a1daed733aa925092fc7c17a081eba1dad10d73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d7c3ea9a7270feda7cec67f4eea51c457dc883c586071b68205a6e1d84dd0da419cf5de869499ba5fb9a2d65df3b73a95bb2cfd473893346210e019bba5b6be4a4d9039127a5ea77b1e311090bb792ac9939dd06;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf692b6a503fa1b7e146b8d4509a59128a308d0a9ba76dacf62f089295cd1947e810df4f8518c910e018948fa4fe767008b3d0e81095c0945d444b89996b05cbbea87158259193bc4d3c30bb103c794581ea5ca5af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6f32ce09849668a90bb0544c61ff4ec8120271b2c42ac252b6bdce9900ac848a7f7800a40239c4e1a4f0de7767ab791e7232616edd87f4744153969f3718cd2a88891ef0c24b75c5a26c1275375f194e1d7a4b4d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6c5ada3e95612ca722b37aea90a24ee167d15597cbf3a2db240976c2a0f8378f031c4da7a5e63c363eb17ef1bb43783f333cebb88e5da45ccfaab74fd48f7e3cf94b149cf2660e5749f5e933d473af8b5e4eb3e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7cd132647b696c2c638ebaccd8188d2b10133e7a1c3fb0751784dc169ab87489ac1865b60f8a01c0a9c59ff1adc47118043fe2f60ccfa5785d606f5721912b611ff17c4546c5b903460c1aeca47504efdb1c4541;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68a97a7276455523ce243511925d794a18d754a05920c6b1951093649053417312214643bdabf75927da846c493f23315fa639bd5897c8a5c8f7b28766e1c2ef009162d52421cf8e6cef924a2f4a665fb3f00cd07;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45c1aad6116856dfab8b29cf716c204c29042e2581ada6c1c53d9f0f5fd3edfe0d120986692e9263a7d4bec59aa443d689e40625f6277a92ae976fcc475f744414188f7e8d97421f4e5ddf23d3c69a9faae7448f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9266fa9485d7e69e7211dfb8f1eca99a5dc7e8344cd045948cc529984622254ebf521deb1cf48d9b6ef6fac5b19f7a2c4ac656576d3994a50ddd607f183261ee0fb65f0be4d958b977dbaee43cfa1d17b596788be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haae41765cc066233290163d22a7837f3162df13d8618ec7f9eb7b60ab3b7196140acf7e509c7c761df4353c215fb609d99e5282b52c3717a9c84a9d0d80f31cdda76eb72481c5d9ed90e0b098702b01f87ab1f2d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6c6d1bc3e8b0c3514c5de3575e1f5ed7e3471d89ecfed7c2bc1d2a666c0326984067bbb7f4b5d2493d2f7442f7d1136b79baccb7578f766596b108c196e75f8fa935d404370cdcfd8182dd8027270eaaf3105aa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2dd167b6ef492dcc3b689a6cc3f30f846acff50335d57eeaa3e82417bec1cda80d9ee537ad266871a67e1cb5f749baf1b15c132566e626261153185e751b30a2377d1cd05273e84d8bb84396265e2516ed872560;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8815a3d80e746a7bb8e1002c6b93d31af71171b3120a3528c257cf7cef6824e8d955fd8bb0f3966c083c184605c08d81092503811928648c7302d0a1f1a35292042b191c6e3211fb346e5d84cea028e085fb968a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha97ab54881be9b9e523c0fcd9f544ba56e0d8fda54ebc6bbcdc76b8a8a08c14df32c43f0bcacfef0c76704183295e9dc1b36c0c90fd841b99d15cac3e3ad84710e9e46f07331cb0821239673e126eec38aaeee7c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e1f8fd8529f46cdf891378f360e51220862206843ef39b5e6f56320281d8967d30dc35de4932a6d46caf7b8d27448cd5c2fcf1087307eafa27dcf5d4f90a8db9cb156592d6d30c0e69ac5244290ce19e4a36ae7d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ec1de66c40a924539786579bd4d793d8eb12d8778b4e3dd3dbab5dc95d298a7a8392120733d17d7f6b552274dea8a0bf69948737998b4098164be20a85a45eef9fc6c7a93526643da8de7ae2cb6b1103ba5cf56b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf34c60dfd6d7372a56c844f1eab7de9e682b150c3c6301e8f9aae77207c59c4b9a8dc11d49e1d652a7c55eb674b7e312a17e326262e46d677a13038e626b3b641271669a8031198269936c4eebd867e76ccc0623;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1148ef9383326661d6bd8a0d0ddbf5cac68a3c71f5a079147d0f69385b022d6c711103b801c2ffab5db3bd81fc17689cc0a98b23ebbda45863c361df19b914824da08799c9118bc02282d34081ee10929368ee696;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ac7bf5b64491883e9bf32c10fb971ee32467f9f279f0581c0e7a23086117b4cfda2c89421f0f96358eec62282b57f627a49dc275828694a61cfd17aebcf0d1650e1420e1327480333b78771571ff4d6aab52939a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5205794e6b448000069354d09de10e4d987e1baafd2559001c712258fea0b6bb8ca3f9abe87e4220d87e21f622f525990a2fab8f22a6fb024b4d568b240cce1bb20305bd4dc47cb032c619246060b07b6ca8b8e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19dd9ad4cfd38f1996df2816b4d6f4c93e52429c068ea8c8c167a2f9dd1717d2d2767a1efad3c0f51b91e0fca4c7c33103fa4c1fae8e21dad07955f5a6674709a5353bc6a0c61772fd21a0f27e69a442286449da1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95e8e6a62583db92e272174a2637c895892c7cf5c2db47991284e63a52d943800b2f642a8b54978b7bfa06ef77edd9f82dff37a69109f32ad7e74033f1984eab7fb1e3e5386f6f5d888e81d905643af9b4d5945c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81558970b999748ddddc1bcd0437dd681f9d46ecdbe015eeb95f56601d0e7c65be73e843a91c328899d57f1a8e34956328c4b876ff1098365dd59fd2ec814161d17719cbecebae998ebcb92ca3422c33b3d181da2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60d8db224fd5c85b0ef3ad5fbae90c3425b7b58b12d200535d6b28f308b2d785433807ca2e64f978759a3bac311161c0eaad43c202cc2b23cbe46613b2bbc98c96ee5df97962d96710c8737759e07895dcc5461ca;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e816320ca705b26fb75effaffab2fc5604040eec1376ac233c2ace042c747d64cd33dba51f9ebe4f09c87d1da9fec3aec77f7dab93a9b8df3f279292fb19d59d3af801b9ac82e0afe8fda21b85f977cba15ae88;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd70ee58435f3a2cc66d1e75c3a992644410cbe24130e9f97ee3c8d943a58c8cf69e08153608181809de1a8b0963b0d9805c676187ee04a87ccf440c7a2a919b263b141c3f3e24f996aae91a44036b7c55a066b88;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6bad8b908409695d795298c244bd926b548059bacc9cfe8a62dd7b82a22676b5439c503348a8b410e07927ecc2abd13d78e76fd769e3300208adc70fd7761c863605cd424923891248c722874867e63f9b020baf9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa646602e5e62f7f5d54a6249113a3a39d16bef143d13968faea91ba848e3571d8205d404237765b4bd411a88f1d78a31769824744f9a52f23e68a14fb125ab0f1bafd6c85bab4ea191bf0679eeecce159caec67b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c0711e468d0e9b4f3ecea0df6166a8a8f9a076f136e0730630f6ff42bf701de38685124f49376340d8898167c767fbea1b9f0b9dd8508897680a16dd1bf14e1c0e09a73eef5dd98bace8bfe66673754108a32680;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd406ae99b27f9c07a622b86abad67b9efd1e5e3ed12d56889227b49f51df748a243c9f16750121d17e598d5acac2aa40946526cbb0708933bdbb7f7dce4522b04fb4f6d22ff59b4143d528e300a2478d1730f9005;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9393a289aaf76acd43a9e964e6b6addcae14812a73d8ae98b84af7c7a115324e598c783f64041f5bf39e8f1fcd690017144545dcc423c69805d2d301596db67fb55d621ddcef11d52c2d5007c8ac08219607154a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha87c4cd654bb83bc465081dbb7e0a096573b7c0e50da29969787f4312a08f4074414c49d9567d6b938ee4fcbd01c0d576bb573d58b3f73a5dc1807e2dc4a14fb572c1284e82a098b00fa18244583c7b0d8d4897a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8c92eb938189282ba7bd76872739c294128712ed7c0e3996aa399273b99467f072c15f688f8ec774fca99546fcb9b2d7bc5732523eef9f0bab70a08998fbc1f944520efae7572b3bc0e48a659d1a67db824838f7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6be9b370658912f9c93e0c890608b09bcd36b38920dd249279fd5c342a8863774619b13c7e06a0a069a138a3c31fe71c607b62046b65c4329d04ad26c6207083d11929f0bceec86676f02b5cf31717b5cedeb0ef8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc69566dfb97a9f9c76d88d4238c6d65c7db1c4c6c67b3ab69107c1a039f7c6e75acc1a4ddf21b7720326f5f03b3a029322d44890d36a40a990af73b40820c59b4b6bc17c89a43e7a6240b8eb57bb2b34c8d6b00b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdebaf9351e5797bbd82f9c2d3449c92f89d3e0301e9ed06bb76a213730e6ad289993a1bcd7591a0491136d925181d66ce5a07d9ca304cca47506941588569f7b6e285d1ad27a450e26e781c03001635e283cbd491;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h100983207b299573437f2a0e4958d9fe36477a1e021147ac5414ae91883dd52b179f50661eba890303700ecca07106f1045e6feca6995defa97015baa8ea710b768bf2668c87cbb8f76046e77ada3e19cd2405880;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39e036b8864e6d603603ec9baa8fbb4b454d10d75b886586b89659a88bf693b76cdd0e7efc3573042c4e753dcdae649ce20ea03fcc2abfa9b1baaa7bd3bc73f68d16565b440b9677bb622ffdc949c6276d4581c21;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he50da7ce1127488a232208c8146d561a3ca63de99012e7ee533a46a1971be174841a0ce09dd299267e7a5e90e255af60a277e2ce989a5578e03e36a600659dcefeb7b1e716410de76cb803eb4dfbc7531ac9ef2a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1616bd700fcdaf2b0682edfed23f77abbd69bc46ea5cf7368b8684e858e887cb2407f4d3d13216d8ff455586aaa0c982a9b66de9f48c31b91328dfebaab17ce8298b7fc751dd3b9d3d54bc36dba906c4165ec6d75;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd50f074afaa030980cbe2d2ee1297a3c1f6af7cf76966e0b1de9e449fe61c056574b04d035a0eb3328f31e624e8cc1b162ded9e15a92bf62eb514f3c65d0ba39bc4e4a22c10d823c73065e4a538491c022cd9389f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0ce1d2b0e073df69db3a4a3762e0f9e356dbad5e9a6fa524e775fe1ee2198a16bc598e561ec3299d2cf24d43d97ccfbd8201b7ac2ce6e4dad3570730a3bb4c64a47c5414bfda99c43480514d0c8244d6135d74fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h229f7958be0d1c4d69e7b03f41b5391404377584244bf12fe4f5720f980b932ccb67036830af8144fd0d569d6f0ecb807fda7f71e5a57ca6f6dd8faa189fd433593a64560f9a4e88c67220bbc6ce124cd9c7a5d78;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2557ff1a3435c0fff23eab84810f27b895ed2728880ee98c5ba73c75723c0b15e371aa87eee524d08af7795cad2cb6e9b706fc40641d7b32e9ea4c4b18a64f949308ad371ab25a800b0f058a05d44a2089bcce038;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h383a0df85bfc6a75618151b3dc0eded1e245b045eabfd11d0cdb6ff5e92a1cedc830c4c2fcb3bc54bee1fc8a8836b037ef1acec3e2ff069387893625ab8c4ddeb22b295a19a81041636999b3b8b645ddb61baf96b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6aa7034c60983608739af495fd84bc0c4a319359935be40c789bf633c757794d22a221ca711b3896224d84366099e3d0174f7efd2a0a513521815751e7f2ed8810c1440b98dd16d0fdaf0d2101ab392336f550f7d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3100755c4b2a61006441bfb328c220cd3f06aa1b74fa8214f1f58b0d954330971e3e9fca7c11416b90518c77bc221cd09a0c0904d34962836667bc36f7e563d3e0370c46d6760e45c0d7e10c5a5589984c132d8c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8439b2071923845ba8dd82c0719c6f062cea714cb832fbb482145f2f551be2f71d05094c29b3cc1ace4d6833ed7c55b4403a8cb39a8b3b3f8de9d77035774ae1902f4ef704c6c3b36c835e490fac35f9ef5ec509;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46848dc6c52378dc14e0489782d1e4279e4b5e40b5c3c035a164697c353f430e3e22a563073182a076c06f43ecf26d4a9b0dbba9210e05ff4149a0829337b05b1f16ff166d73452f7b9f435e12cdc08fb1da3b990;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h293a604cdf46f4e35cce03f1f793ae2ba9d06c04217d660ed9feb1f073bbe48c230bb74f75f42a9138dfd4c23c94ac5ec4c1c6a557896e94777d5f99fb99f9e5a24a47ba34a6196fa0486ef9edf78f7b326021381;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a82eca457bd904ac82745656a5ee276238573c7b2a1ec97e20e4207b14087d8f59574b74a64b165d76a62b08632ec257d0715b1051c8b651006ce46c5b4bb38de82babe3b8f9af51f56495338a67b2a7b9d35f41;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31e21c4c6809551793efb5d18aae076bcc176ea0702933129f1aa1b61888f3bb63e3e825f59e9919c3f8813f65f0992110baf7cf063f2bf5201405f0c19d3c9b5301cb8bc854071c588d1b693c8b7cbf28aa62be;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ab3ba095b0f8ab3dcc3994952cb560882ddb67f71e17a021e81cc01568ac9cdd9ae9bd0924abcc35fa71099f8e7bf7c510f2ea54c968fe8c2c1e1a415a0eff1b22fd58e8004e225116293e7e3834900741fb59f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8729d228a6a68f48eacafeb8d3ed05ffdf62458d1db172baf413fa50b66d2978d815d3067b9cc7f32db151730f913c7495a54e7e6ae30e90f54b98e5934fa7a2eef096098098ab819674897f35d56ac1d5d070ef0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h608d3c47f217c236bad10b6e53ad40a361b58bd2ec064060168d692d9afdd729cebe75972b14d736aab9b6f3960635d2d1d54f83a6feb6855a00bc322d1650fed44df4b49ee0ffe7abad816e109ffb16a91ee5fac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d6f31384c27fc89708166e21574f630c50319a6d3228a7db1b161fdc75a3e49926c1ef7ecf6248077c5ca9c4a314b103446124342d453fd9ab932d7d9a3c9c1623d8bf81ee23c2313bee8483dab22fedb09719d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb18af69c8252bfcc4d062027c418b109a9ceca013a1181c0e4849e834b793c7ea3d2e374799812be2d73f0dab186c17d21912ddb327d3856e4c389e975d3859f4c6a3261e1db86ae2bf02629333dde0ec4d515e57;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f4b32119ccafd30c558ce8dda2bee83ff7e27d33b64d9b645db2b2fb3c421b05837ab0edcd48d23f893ad1130c78bf4edf306548f43d688909ea73c9775d14e854da06178d2ddd0efd130ca00bf907b2a3483c65;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc17729161d965c4359aee79d85c5c8ea4638c349865cc22df90b91c74512cd26fd148a174057885dad20f2b72e29fdbcdc40360de986fa56bec33d7cd5098d3bb0fd0013b0fc0c15a760e47a4d4c7385a405d23a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6d763504fbd70416d678475ee23d0a1258d15cea67e5e288f3bff88d66411aa765ababcbdc32557c5a5d77c4e0963c9c3692936bf8c09d035915eac7f708e8d82eadad67581f9909fc3b5b5eac294ede5830d3b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36ad36642cc9e22779dc70ee0632e9f30ff87355d905c24c55e41c265654a16cf1b538f687f603138da1a818bcd97e24b8226f6478705b665cf4c86108e47f8aba0d3a0046f1f2d3fddedc1c33ae63ee858d32b82;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7a53bd1988e3144d45640e8fe6a9da6eabb4b908953de19c3140471178f14043d943f1b11f6a9c851e8eb8274a452ec8436b0a1f7db7947cee6884953b1d9886db0c0193174f1ee4cbe3a464425a9028d8e51263;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7aaec2e83c4a4e9a8780f0d2b8bfc77f467218c08e122d85a464de3d0d48428ea81b04a46390957468c40ba16dc09dedb3e0a036e4c94d06e260a3c3b77fecc24c52cd2416aa7bdab613e31b2666f25b749cc634a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h727229adb79bbca4d43c633964fb3368e2f7eed367ce59ea151c6a73a92ef95e5c1011ce2ab259786fd03fb968fe859028f5edcbc3679300366d673eb75bbdbed76c46dcc5bb032d0ab2fcb22c1328fc349a17092;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h433b801f1315793bd0e305135aa7aa0062487ac44fc7879986a0bc65b4c9a7469f62ef4d90b3921f5ef5fef01b1ac282bd27eb3ba17917ce26d791eb9455ecfbf454f79560718c638e44f8d274e123c3f3d6c8220;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb25cd2e8eaf1869a0439691530f78409fcddeb62819dae27faecde470c150a19687d5bb0f4bd2d2fb46512a5d8077d49cc2a355707b392e9108c901f2a8814fc462ef2cb5167bd695de34f30c367bc12a8bb481fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h581c3625dc89f882695b2c63450ff6ed1b68c78d38de88238e5cb89493a01121c0ececc3be6067beb5c0679ab34e01127d02ee0f01fa290103c5682b010fca240915d306f658173d24a67d3f9f2fb70636a1c4250;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f137f8e24328fe8f7c6bca7afef6618ba0396f952ef0f208aeebac6384b38cfe59345c8b935572d3bca86ec3ad76938883f1e393dcc9667925ed78b95a390d50301eabdef5c382c74a0068134283be1399ffb570;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc71ecb78ac9290128bbcc8c0ebd53462f3667d91a85b2ad3927e82e885f4041887562a9ccefe61d3a34bffa394a4f5605d4c90a4551cd68cb894be536b8cd55aa2e5d7d16c7fe6d600fbc54dedfbec8ef385e9b41;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70becbc73d29cca84885febee8bfec0911565bbf05585adb2dad918e30a5fa0071ee75e4bba1a7b5844ce0c5a2e9bfa9c7611d7dfe4ea48ffc7c81c0800b1ead67ee4a56e952c9371f815029314361ca1bd6d4ed1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc3e45800c4281e765c8548252e55e94f97a6e0de0819d011e358f652cb9717842b6cbcdd911b58a7fa0566187f0aa17cb10b96e99f0f6a910497d5ed5f701ef2ab274d6c0f0e64cae018bd09f6f810eea37907ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15873016067ee478959159e81798a01a75abf1d9f3598dc9dfcc891fe90cb2111530c8e1f4322b999920631973671fa568c8b9d03182cc33f1912945e9c62fb1baa4be27cf82c67ac32ea6be3e46adad4ed998535;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2df67dfea9858f28cc3d21423c6cb4a2d1784cfe5f5520ddba829c381b152a20e500617dd62fbaf039b014236bb6ce761b03db5d9551b6fb2e8ea5569adee6296943721a2a496e43a24114a7ba9b40c3b607692ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h190fc4234cc7a9d3345bd414f7090eb6f2769c6a0c20e8626d8f670c8185faee6d487702a562d821accb7d7511906ef0cab1447fb6a7aedde33cce1352ac76a7c75b50898bac4bbaf4ea2b38e0e7ef8095fe69f06;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72f6a7179130e0a0cb29a2844e42037414fdb4a7a77f719ba99c767d7545ccde7263ade0b197e5fac323ea96c6c9141f30aefb56c01e3c6c3f108c799692e8856cee38155dc2e32e375ad5c600e45ec542ba2c7b5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac6f7d49bb6491a99b5c7958933122f6fe430b7139a0f70fa7c8fcf2ef610fb70ea98fe75306ef96490c3a7189c71f5c4b2ce58c0f9cc0c1d1910cb7b1eef89bb8b24be9a7c054be67db40e262b0563425c6e09e7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbbf7ca190f3194ec6542a8490274511c486fca390cb35b39ab8912f3cb3b3e86a27d63c92f2a5c5426497d3838b4dd97dc8d646ede17bd2d10f14107a4156907ab76c85b3e756cedd5fa6e0ccad6c950a3a8b97d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f057ea29abf497f0d01a2cdcd1d25220d2292905eeef7051e000997a5c5658e991eb8e16ad502a850443d3111116ef8e8d71ce44fb55ec9662e02d3ee596f54cf939d975879a68b65c34428da9a04ef19bfd838d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfffebd7c25b52242c31d7da2ce8ca9fe082165b67b7467acacf74bf987c35c5883459398a3f6d7650b1eb857a08009e92362bf5145ca2952d6c07637f4f697cb644aed90d30ba961b01adc954e5863781ff71fff7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h33d6e727ee0cf9b3bd89008efd6ecc56ecb8a76d148468b578879ecaf538a2cc00a4a2f824cbaedff423bf5b449dd78d24f3c2f3aa26ca5a919006aad4e1d2e2c1d43fc3f7e0860a1ac766fd26341e2523c078078;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b40c6b9dc318492af57dd9396f65a3c3d9e3471b9160af1e1f4c81dcefa74fdb644b8c5b685d24a00485f08530359abcc98199181b36158b11a5ebc87a8d3cf980bc4cb15123d31086ad3f178542ee5fe28c9a62;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b4e6af0b0fc57a165e6410aeecdab375906f9a7c9e55cd386b3928355de5eb39db1f64634d18e040e9dced49fec48c2e586512f5bac08ca350e122a27ddde48a1f439e370011764ddd7d4ca1fbdcfe2889c8277b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heef29dbd30ee58324593763135d46733f79c9976dc5008711bdd1f8be5eb065e8e8d46df8265988b8a0d63e0a5005adc2c109980e1c44d72ace6ce286312944fe0c3c63e9a3baf99d6ceedc8ae25364286e64313c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h977dd51f93325567de0e07cb1a56c82c85a548f134d286023c521536259ab7a45457695e581dad1f08a6bfe7233963f038e0212cbb33cebc7b8f106f63d004965268a5da3cc2494f3b887b5b7d8c4d10b4f4f862d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h986b4da283815577aee4e84c5840419e527f36f21210f11b7a9f4e0dacaaca6495bec7af5f9d318fe91e746c0f500bc755ea6eeaa2689f0134b8a1db6d9a3dd509d64147ccb471d179bb597d35e08d4feddacae52;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h800e463fa5792c39f82a0bd02ff668df7fee09627ac1d77cddc654da8aefc385aeaa89e26663e5ac0ee8b7cc9efe0fedb450758efcbea21e72000c29cf40548c89746b6b2038edc687b865598fa0b55af616a9b20;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb65b09e1c4d85e68ac1d5786f848e8a422e2a3b2af254fdb443d46cb03af9a9aa2a78f788f43433eb7dc49ea6cafa3967fed6f7ca509307d789e9c0cd6c594384b3c9e7974bc1fa71b908b077eafc7274cc9eea50;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ff2e53d62d843557f8bc53a7efc22478c5e344b778054f4a286fb563aed51c3860e09b69acb7befdac51179bafe2cee196cce1e7867ec0b674c0781321f65b983a790533ad234cb9ccba336c67df22a5574cff17;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he33390187e21b268268f6f63daa3331f6beff1145d35605e23313446043606026d2133809ebac748a8d4fbec48219c46321976a73325c33f04e224270dcddef07f91870a56a6e6c6e4949c3238a26d2480087a8fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41cccb4e2694028b49ddb747763db672a624415049974da3afe74f8bf5d019c10a359f0c64e2957b38aabedcf96022dcca7d7a1578708f88b2b4aea9576ae2a6cf403977f3b3799036b873c388eaef99cc0c31e95;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1326cdea6520be286bd6ad274306af56c17357cfc4c298cd7e8b22328902414ea12f67228439bd2bb43c09b2a4bdbbf61ae76483816d73d33da555de1cf4b7bdd22c8da03199ea2fcfd8b0ad552ee3b56b3be766c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddc13fc149f22514deba88798fd2f5401da660af34b478b3a11d5cb11684768f3e33b0769cd87465e6e3af88b99a5edb052f0107686a57f78b49f1bad025330a649c8faba1dc1724bf3f3940757fe600ca5ff7a8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h615149e4c3719c08034afef3f92181f527507fd85aa5ec3815d5b0306960929df95ca57e48137aabf44f4cbb175cb415b2cedc862138e58fe872d9da329825fb3d99489cda865af61049e849ef62fe577031cf3d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he8978ed121927b8e1c7d21963952e1b55d9da7716456bcf932d9b6665f92f49c0e369b3e0cb1ded2489dfb6ce8e6ba55eb2f8143e5c7d826522053673023b15dfd87d68fe7c0f4bf7e1f425116ce2df0c4d1f2693;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d846b806875ecc38fdd6d4e5018b93a76a913797b5fae155080907a44c1b45163ba19eddf399b3ce68d8fc8e16d233126e5d983941668127ff246db415dfa830f6f6c9fb0ae68e0241595eb2460acbdf17d24e5e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b1c94902f3e8b1f1d4d4490f20af34187bb2dfe6c5d402a10014ac85ca466d1bbd5fb82e16613ad452a8dd490ec1305f518a6eb3773751acf1449c1ef3eca9ee5e572b4fe06f15170d95262915e8b9efd427641b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5141928a85a20de0225a06d74b70e3e9fa78ba91d43585563be28dc87431a785a8fa66f1647ea089cfda027bca56ce0c2acfad177d656a595f66429c32dcc20721ed1d06307bc3cb574dbc34246172faa8d4d2322;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5886a52ecb8e4eb6bb3a00ebe1dcc3dacb07aaa5660e7e74b57e02f29def6056bd5f45d7f5e2a598615b3831a82e6d0252e672f818bc47f0a9e0e4d5b378c659769108b091312d3d7b6e916c00a5a89c489d44ba3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcff373f910bf210329b124f560cd3f92aa0c601e8a730c231abda779e0c2ab8104a4c494422130dcfa4a40421a8caac5b4035eb4f6b5ac54d206195171e2159377013ef54b4fe37f0e0c0a7a74cc0a8a479c0e3d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h797db28b42778f1994d06db9019ea4657464a56abe3f2dd1b404629a1eee691036fe10101860ac61ff1d82624436213d335b60d4ce419b15eec93fed209e61cadf1508c114907f9ee114103f1c5dc369183357ba5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb316d3b4b90da4bdd3c2fc41e462134110094ca4704004766ddcff9e2402fd92e4b315fc48e202af1fae0700624ab286032b1de52c364c3752b272b7616a54fe262c7f18af15fd14f10bd72f817d9fc7bd5146f95;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a115f85acead306357bc330f00bbc6da9a125784b6a34b3ab9f6266fe23bf7b49baf3c84106794cabdace22c9076af7d5c28b7409519487381864610b98653a64132594f81edfbcd3ba8259d04a6a46d9ca0ba3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h391803829431cbcb536000c3f7d9016e5431a72855d91e103e19aa13e957aacc32831c299d00f41621c95de29502e531dfbe4b6c9ca8772c8080b2a4232fef59efc56dceb5b3b0bc71d722ec535ed813bae242bc5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d85f1e30754b5af11dc1901e98d8edacda54c1ab8296c8ec2dca294cf1946277c06fb2744172526ae11fd5c3cd935cd1501c01302e9bbd939fedda4ded26657178d7fe7abba4208aeb81cb0c70128caa46fafe35;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h575a1193294df3c93cab768851f1ee0cee3cf1a323fbee33011217a7fb5c5c0517e6680e9b05ce0a238a400ae92a90db66530ee0300f5303ce3c59e1aa05dd3b1e961995475cfa3a29ca26371625c291a75848ddd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h986672775b8810d41b1fb7e9ef30d5168f9f8dc0680ab1e2ff4cf0ab3c04ed1c9e4cf8c4a2b2a9d65ff14c3a94e587ce8c00fc17658f05a6695153901d317ae7709ce3e76a6d0d221318b87e6834883f0d8319abd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7d41a659292bc5c008b6b4212db1ae7cb05f8014add02cf88c6c67e5000b5ac26720fa4fbf1547156877e640bf31db8bd93ad1d3481e316678da02bd73d9d7c78da026cc1f8966dcede3c2ba38726e415bb657b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha359a894e7eb331f43f178d6defb374e8525eaf4c7df2228325ef2ce35258f94506923481bfc8a3ea8159d33519275c8d89e26c53e70ca854d76d4721f7f2e96299d8da768e5ef14ffd5aebfe5f5b4c2c9aa3f3f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38531b57e8ae6818e9e0c451289c1c908c95f7f63c78909f64a06d733ee0364f1c84e38a5d74a07d90cd7f5250b1f57f2027172ef1ea8869c013d802663e60b6bc4c272253c97aa92d63182b3e1c8e1929c57eb0a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79daad04777beffe8267caadb98f4a7eedf39f78abd05d56b702658484a5914977429575dff4a66cabfa15dd1f7e5705d840adfe105a37406622d6071200b48583f22366544f1b26abef99a05f43368c89ab9cc43;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7e5a22f4db9b438000517af88c2502d469f0dfcbd4be10cbe28307979a4b92c3cf14bec555b6d02e738faf2dc955336bb2e0f805d5e21bd97a6159befb58bafe3b6b40771e83c36e86b83e35307e2fdea8778a47f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f4d773e745b59407cc5bfe641474a62d09c85fdfd3706dfebc39a3224a15cff6919cccff8fdba119226db993f69bfd197aeae5f65bad2246c6ab598d5b2e2437c5d6df8526b9420d20d120fb992da9730191139f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e327b4f4ee7adbc01d05cf7887052e75f1a6ef87ba5b245dc034b08b8add5322e4cc624ab91d9addf737377fee15472b0730647839913ce17db8b655c62480e78ef52feb8f01b5a1cb49c7dbe1ee205a642bbc93;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf91aa1478f97dbfe11517baf53edf78ee5867434432c66f480ed940a0f7a09d90537d20fb475fbe27017382321b2bbb95708de4c95d09feecb5cbdc1ab1ed96df0e927942c3329b27cb197035e4527f39777a5d46;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a85ce9b5e8002e869e1e1cbe06d8d57d8cdf60b3222f9e7b0b558c9ea681ce86449539e740b585bc2d53c1f51d3e1978a1417190b8322d3b7c7db2b5b09c392b7518dbe452bd5a616b2bc569edd788d780364c83;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6a39e96b359096eeb9da2af36f7df4661f7633ad61ad97019a15a2d62526c312553de9fe2e5321e3c958febfc22e996dee579806da40da7271068b2120f74685ea266cbf753e425d616301e8ebb3659b6ae045c4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77c1de62e07cb5487da4f0c5164fbe74798bdb326e4f69cf030b2c5d83fefc87e2b48c07977041246764bca12e8c4d99d3b448b4958b5871cc170e25a751e5f5466a622348886e5d184bdc3014dfe11977a36d8e3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb04b50ebfa15dc895bbe01e51bb9b3b805a89a58837eddad5ef98e513cd0a8f89f4c9df7f4f9ae30748b00aa50bcb7712b5d816ce49e1670b82115bc8dcbb2027c70ea14133e3a98e8096e11caadcb03669c1b06;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f655d349c139652e4cb6ca4822ef6368837b6da41ee6791e5bc06a58fb9384fda70ef147ea9277af79e9dfe9e588be1a296fd194c5075697242f1799a716eebcdd7ca20c6f30c70bdbf0d7fb6ed2b9bb1cf6a03d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h25dac45575158adcee8685fbf3f60f0119e32d60ed52f25b6baf0a7632b7b9f0e2a5feb528431db48a9062dec9b64d918da86a6f87d017001ee9a2ce7fe98f73baedcb0b4fc162ae67b75c0e7e750154350ecab17;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a908876e524f83f0a41dc85bb65f604fcc71ce69f67a06280fe23b9db0f789f5985a04dfe5428f4e59dabc0afa519d060654239e6f68f4eb267e59dfe581b22f2ef464c787a33ee575e035372d08c9fc67c956e7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddd9a96903eed0fdce24f80da4695eb0486e1faec9d5197a6dc559386c8db92377ca76414407c66860a3547a26f0e09bc2486992c2c615aa6fa4e66e1b2b8bd1ab4b0bc6ccf43055e0c662013bcefea140e7e2220;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf13f9044bed6c90cf8680327e76260aa1e1a177cf8144260d74c4c51069091862fd18e723a6bde16a9766579180167cf34bb68aae88befe664f1c9409b9a0fa92157b50f80a62f3c945f728484381cb2af58c4470;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28aa5af5a456da38cabef75db1c6ef29c93f230f6258cb9da50276be54829079d60b0512b9fc477a1f7990f12326c78b730cad482a4d8fef10479a16e263fa2b758c23cee13087885806d20d4f5179d9732cede27;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4cf3f4adaaaddf3a4793d7ad2c0e534733708eaa984227bbe07df2886484ddee921e40b7051a06a3af0ef30e32bf72bf6ae66a5be6c7e6d6632620e4aa1977d62490a555a5da676dad002321c8b7c1bbaf93e16b9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e83399addd9f2bbf92a5b5b024a5a6ded1cffd128060fb1042b00d5642376152b2965c0c5e9b08a57949188fc35fc0068dfe168f691d17b729515c418d894ce69580408e10194e996f4b23265465d47900691331;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72343bf4fcc7d7b67736d0ae76e2c20c92e6bd6ba867c758fe0fe4ec58a0063fc74baa3a530a3f0a1ba12730e05c8038356eaa3a71773b7b6aa5f9f4bdc9e9fd3edad103dde3b102f1d2a27e80ff03784eb8509e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfaeeaeee56ab32581097e85104300a574995051443b85b574c19a6814aa6d4d9cadb097869e6741b003ddc7e095b3d86a1877037ae8fd1b4904fa71994c589447f366eefcc64cb2f09a13dbdf3b31603e293f162e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd70606dfef8bd0686e6b6d99366b525ca07ae2ee64b7cd56c5374fd20e22c629c2733b32e3bb5073e9bf0aa274af5779e7ab5570cae83175fac6d4c1b3db5682e38f447e85c175d208a5f352fa8e3e639508b97a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc852b09ad0f58d8c09776799621f77247186e92122306534fedb7b04bbed8253f367b360c30494484beff99cd263c7a6659f34cb79bfd874e99d87a55985b8ed2ac1920570fb75e249796d445d16bb4f8c1e702a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef87606237cb6e14bcbad49abfe82599b14c5aadc00bc3e06af5781340c0e02237dc636bce2a82d2c9694d23880adaa93035481eacafcbb18a20956bad84257146c422c5f7dd0bb4f6675c9ba7479d8242b40c570;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a18ef9bb215f2da0d0c8c532222e50820e8b4dc7c8ca2f88a587f833b92d84b8adaf92d851970509edec55317f0545e2b2f036cfc6d75e201cc579f1f065792374bb948a533e7ce62aafc2e72880172b2d0c3019;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfe5d356419a0cca2168429a401c79f11b22808ff04be3f67491194f2a500ea2729d29e734567762fcf44989870827f6c017343b02015ff2a87c0f853c1467a3d1bcc31ae31678692c1cf0494e65fdcbfdceba75f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb50993f1da198d2d7e1c920eaa61ae36fbed179dd277bc84c2e3ab7af433815942422af4275cccba52f8850fd71eb5c988e994702032618e44d5076194610dda3b0987447689a1f19c157053b7c6b43f6ffa8470e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h491e0bbc19af8869016cd7593e985350bd66a7c244be4873b32df4abac45c72df931adc8b4e52c2762db611d4228226faca8bea3fdb9742f40ecb2c428fbd3e8b058be6439633acffee345e059eebe85acc52851;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a53f927c4ff69ed137fe96f157af0f664eedbbd89249ac0448af229e8bf237d8e00d12816811b3d39be514250eada1d4ef4a4fb9a6b8f1c9fcb8d729b6e5564413d365c9c80219b7f2eacf418e2e4ed3fd8c2ac5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3450f60ab5b8b38c6df677a3115a1428eec14ce054884f11422ae4a749e67f094f2708e61275aba2e5e0ef110737fc10629ed7d7b66b647ecb4afa0ad9180729e05838faed3431d15e21de5f210b676d72a800b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacb7830b5ba6b651d70e5eb767375df3cc0f177882dd82c1253869d618750e15e3ea15627de9b3d49aedde25845dfd31b8f12fa5c37c777ba15c24199a553f0856aad3154bfbe29d4cbbe499bb201bb87e6b38682;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb9e5db6321f67ee9355131c722444d90342eac5f60fcc094e273e5ee7ca14adcd1c608c584e861fb04c2bec8813b916c86fdf604ece5cb8b6f7e88545a54e49ef4639134897c87bd68d29590a5bd502448119ae4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf54a64e33dbdf5485cd21948f9a50ca3db38143f130b3e375691f58f439f1f9e8924cc9b6b3600ae399e17f6d97df4b2146294db736dfe2b7eaf434f6151c1c39550c6d357c58749129f1cbddff1f73bd526d3d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h142be3d0a6f5a724d140ce0ad25cb83fa8d73d851a8599576fd7fbfec0567cbfa88bc2d3cf9938ba58d5a50ab833b2f890d9cf99991d77a0e39482c6542a2a3981b28aab4cbadfc087fbd334016bba162e3cdd386;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9a5e779895b9a0652b33c388c74ceb03b3015dc9334fe6721f48884411a474682af7de9ffcb796f1adb82b8efb40e673e0dd092eead560edd412ec93dcebd0b38164357181d92bc23a58766ef4266d7d8af02320b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83a2203a9c544b79ac9bbd5f884c38ef7de61269ddfe22fe3d4cc31a138760f880c3174ce624f31b6dc57687d858e0a00b749b845b7b2d21e9ed8e417500cb9e3452d4fd44fb7e4d2b969dac62ca1c038d29ca04b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf88f413c8b2261682fbd6c422d6333bcf36d4c2be9b18188e458029b78b47abd4d5259c4c9dcf10fd8fd36a6706a9d60b7be5240ad9940b2883f1513be2585dfb96623bda8bca8e48961b8573413f97f55ef3a860;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd80e060972a623da876cbc8f186a15b0563e725845d6922a98584894f47677332047d5ee0f2804ec78b7fdafbeec217f3b40f1334ba423f4b377999a29d696c60c9e7c255f6da0843c14991310b95a19826de57e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2ad4813c4577889ee7f5a41303735b825176e43aaabed2cbd7db584f1656110c9739d079aff8c4df5f8b4b315f56e3069fb5e76ff237c5fbfbfb0737562657fca6a90b27e5c9ead860f504cfc06a7c6fcfcbcf4c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ff4cc2741e36e8638f96d3ec3973a693e65bf76c96d4597e2c6328bb92aee54113240ea0bed505a4375ee59785693cf995c204bfccdab3beffabe59a01d5e2c11a7ba0c161730ea46ba19e586a5717c10ae6a0e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h212146628b6de80f6eb0b93f738e9135ad5332d41d3ccc6fc24139dac8d888bfc9e8d48c087c02aa04510620ecaadc6f1256ed4d2b4a19557dea2830508e12fef01d0add26f1fca733fac7cdde5d949e1c58c2306;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h266900c78db4e1f8d3df3d2a3f2f24f5d0f9a8813e5ec98c0b3d0513dbdbe6deb206f27151f89427e456e1395ece6602fc82490aa721de1d8325081bf9efb0e77fb139bde13872e3b7b984e5475ea85d1fe22f9e7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9209dd4368eff9e76c274eb9852676f5f0dd87b5db6b79fcfd538c7eca01b8b78f19bd210de80ab6792336ee29bd0d8ba53f2a6ebabeff3f95a41e78819fad23ac585cc5c95b8e1cc78b3beb460e78fc176b7ae5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9824a736776b9ed42ab452f58f43505bd31e8fc5c2ebc7d0975cacaed218fcd440a28e39957895b81784e3a3fd21085ac3402dac4dcfe6d59814307a388af9f4e6f82f6ea9714d2505ad8ec181823f8d6191da75;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h308de94a79656b54e7b0879381cc179a684d0c3c789fabef67a49452dfde246bcccf917b322000b2ee2e9c44d987cc0b02f7b93be68c1216f0bf124f4bf6641befc3e4d6caa7dc10631d037bcd6c49e831379820a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd3a51e84b085d8e922701eb802ef66a0df22020561974dacc3e90b7c4b00de97c1a203417602232224143b78a8ccfb8cc6625f7cddbea3a208724cc4dd1cc554ec068e478782d6b5dfe16dc84282cda1ea56142c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1dd790515de5c0175e2855d1411807210fe6a873d4aed5f554497cd6a9dcc5d49665e3520f95be97e2b03b7dddb2e181c937ec4d17ce5917c2b8abcea6089d55a92c5ff3c1a15a447bea555d6534990ed193112fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0b081836d1f6b4b23acb2fe53a9ad1b48fa0497da24971f106a9d343d04ff3db1d83a4d4772615dc6af2e5e08032f54bddff2ac15ea3cea85b2da052efcfba5798a9ff6797a2179ff73758a86c4a8865b64cbca7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8c43c0f338ebc112c22d26cf2667533322f384bd171b47cb2597c7845ab11c914a9d1e8fac711e983a6a1498d5c469eafd1fc0210c4a966649eefdf8f1b2418d2241094ff931fc753ebf1d7b6be5974cb2acc8b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc96e09b985947b39e40e11f4198fc03e86c13eb00f780367ae863be5df75cd922dafe6f0987557956b13217cfa0a5a31ff631e66e329f1e000dd5cb533664c603b7c33b9f6cba79cffd2795e5e271a5e9fdc92d4f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h14ba7b68c9fd57f8a98716e4363a87a7369664abd6cee041ec82b1d4d0f58a986a0d980688ba86386a2956eb46c18d35bb123400ac4ac0c970789acff41e6d5a131efc85482dd3244c5e148313673755fc8641e9b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1022474608e51c33c44f93f1fb97feecf059b3be1e2be546421e6ec478aa710f5de352df3ef0118ac70d588d7c9aade711d778fc588bbbe9d06d8f2619988445a51572da861cfab9c98452ad1cbfe20f583b24b50;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he67c5ea279b5dfbac8c3375887df9536ea2410596801399c8ef1c344ccb6f22a0436568642c44a42e6ecf9037319532d64afd42d91a89139b1c8c3f56ce5ae69b1900654e4c7c086196e4d7a2d10b9aab49d131a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h266b2191693e256ed56e8df9d5dd766fb68a67631b80f92c43d44145bc3a4213f7474a04871586550d15c71b39d27a8dc24160089c53923531ff37888a230cb144eece061d8a8b675275610f5f2b1737c46f4ed39;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a198a9ba79ec5a2f9a87c040623bf64a68ec401b7edf1813c57521174841573de538374449b04363bdce5873793447c7c53583e124348a07f7d84dcd8375608adfc4ce9c9d2e8a236d211036090e9dee866aef1c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd1955fa93de3ef12529e1c4dd9f52d5d342440803156d488291e8fdea382822f2009e6ccb52ad522d18216ecd51576a19603d0bbe90773ce27c21e3bf637098c6ac49b43e8b3bde6c7847d9bab86b1ee7815cdbf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h586921569506dd017b078eb9c09dba1ecd730409b396ca177e1c1c6184a2479a1ea174f7ee5d275e52ecbb3080466144a2ee6c21bc8bbe58cded05ac7cbf0ed4ff4a552b720fd40d85b6a78c03a0b313ded0da73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d50d29c59fd6b1f84f0bb8451b6a5e8a4af832ca8b45ac527d9cbbbdbb92c2bf6ac2b0ba7f162f5ec0359c30157fbaf25bdb635c25e68d6c23ef33c21a5aeae7b883f004521c112a04e63dc68fa26e0d1286d4e3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf6cfd47e13f39bfcdc4be650b54a6387ab749024c6a52943d49728c166f9cf49d9b0121f825f3fb28740df10a2baae4d840312c63845421bb91b046717643ab28d8ef8cdda9f06d8f1910d5fce6873b55924350cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h519e5572ac36689cb5481c3a99216fd009bb64930fd211cc641e8769df37fb764d42df6ea811e889e3ee154362c81e096ddc035385b0ed69eaf25291c835e011d3f649bf3626e8080c3bb53f93ea0a0f17a073462;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb822b6916d66c7a63fe2c7cfd405330d7d99ed197dedd1346c44a201097da9d4acb1ffc70e6aa59a9e97982d5bb03dbfee31324ea44d7581d225b8372fb38f323616f8196b0d33e168119595acb530ea0be6025cf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a2764470272e1a7ce03513128955d85b85bef34bbd60ee9a78d62a2961f5de64ad47774a5fe2d105d42fdce70590e5f81afa320fdae1d90c0d941d576c230d95053a1583b2fbe611edc0cd33258a2df5df97d90c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h855607d7988ccd8af46803f023bbaa8f12d3630788c5b43dd369bc81e6540e4ecbc5dd7eaa95736ca42966a76e3b3f99619396696c1ede5a4996dccc932cc270ed48e9d5114d2a3c04c34ae9f4c71ab4ff2792658;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb9ff5d2ac5e6da02e9b91185fb80e230f93dd8ade36c80d56bb03be3e269096a53aba9d14167b58673e141e98f28f165d70f740cac435ae5d4f7122d62fdf15ee640330a8e9cd3b8060f9a0949df9879ff24f90e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e350aff2abf54527a0929c49bf9a4e6729c5e4b0cecb92f99813bf7ee84fa7cc7ff49269f3db158a3780e7c632588a5eb9e04a258189a906673d382687014a680e4c943fffdd1698c960d6d37827b033d6e7e2a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ce6ad1c75bd302b7c7688eebaabc6b488600ffe8a19edf0615ca2841cd5636fb5c1c6f3e43c563553d5712b6bbf291b1507df5303b565fca75b476ed674513928a8ecf5a95bbd9f2e6c50ff8f3c1fd44efbca31f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8775bb41a43883010daf2e45da72c4454d5fa725a1df4d6afb90ade42e64167c956fa8d8121f7050cc4a9de8199fea71b1e95c65fd1b9ed2d472bc4f5be7ca808a9ba6bd030af472f1f6c60eaa1fd9021e12c0d61;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h445988c4a3316b549498fdfa62661e7a8daba606b0bf0826f35d3425b899eb8c627631f977721a2bd52a65f3652ec6515ba14f0ef8c272fca8e5718ff1b0ddb814cca56fb813856cbdfde1b98154715a1521fe8c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h980b9516c801957b7a2b58575f23409585eeec37ae65afd0e64f2f3a32d95d808d8bde27d8fbc906592582f693447d1bd0909f25bf53cc97d8300c908cabe62c1041d144bdf9fe21f7782f7efa1d7ab67cfe3345;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ef666dd035b552359ad593c7ba606a776da0d1e5f9f47f3fb7fba59fd19d015389f6dc3eba1269972e7ff90ded20d2b535b470887c8e5bb49ddbef6724fe01958dc114476217b07a8f60007510960bb2a275dc6e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0ccf28cb297c39a237bbbd8cb13ef1ea30a5333a792276452449807338cbef22e2f52634d2791b28610719d78193e9c6a4712d4bc63d1d9ab28fdf1d2dc0f6c27d7db275f44f561ec9cc9ac85024248bc30e5d12;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79f011801cb190e2f2faae4720c631a97964161d94f9b5d11ed0e608ce25220b501257bc7a720595789818ffe2c8597437683710ecbdab876f4e40d701cbce241878b97b81efc8e4537f395bbec2ff1454cf5455b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h180d44adacbf29a78df54ac4c37edf1764f94593b529f4bfecdede009bc3bfc84e230e93c850d5598323cafbec8f2b364f62232b89110eaf122bca38c3a4c978e1f602c9b03b1df5043c3c560d7edf3bdf13a9c90;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87b7673b65034c7645b8a6755837f1ae7543e5bf6a5570bb1116181d804c49cc7e630465e9e15ce16e9613be29d10855dc6c1d5cf9835210314c7d94a5eb71660dbece4290d380d37c304c07787f41c2266a76e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha70d68411041520b4b047c5f8ae3c654ee3f599840a9365beb92e2f6f6b3ef666497ae58b813945d434a893ad3189b2a18c8f34b78b2db428087cdde1bcc16896b543d59658479f225e56a9360b757f194d86d4d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48efb043969c4e5c6033da4f6be25d2ffcdbe46f0175650a762095ef118e0f1061b89a3ce6b4b2a087eb31adb13809612ddfd3a5d09de060c3e4a1f0c2e3037dbe2cb0a4a253dba275a81e6584e1efb6b90b73804;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h598d3b8a8e7127778e6e7b5334ed799163b96af4ae5a6643780f88440ca9643a86a611b461f6bc77424f66250fb80e44afdabc5c02b868515e3cfe67697e2c7190882bcda0f898c515b8968c14ca95ce35668087b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55a6082cba07530aed0b3ec1e9d24f2abc3c57129abf973c102965bd6d3696ff256b48ae870985fe401ae9940892742ee53046f3a6d1e77203e90b39edea0a6d8a968c5051c1eedc7b345faa12e38ab790e9e82d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd6157b29b4257aacf8d905b2e911e781060a1da73088f0c4ae4ee0e59e89811dd264f65fda67270100ec16bd5fc66785a33c61d3dd0139f55dd15a294699c4c13ff23a003a1a4781949095e55b1274a68c9fbf688;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15face51b5911fb3a6683b687d4ba94ef7bed6fbec7991ccfeaf31e37f6fa84cd484197d8ac89c4d924f195e57b47ea16b7157ccc2dbcfad9b746c5c84b9998db77fa6be1b871e0304b2b274b568a729ef472ca71;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1bc51a1e17f2cf734866ed078e93b0d0676654a1172e4b3b671da09910156bf25c3bc5d37267d50ecde8a53e86edb7d53317343e34d8ff6ab9f906d1fce9aeb6b9086d506edf1a932d429c73f1bb23a17ec8d5f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfea87982d4c6f505853c35edb0039f4d5ba485caad1166ae5de9b3d24e493b4ccf825aaed78ec7eebcc148bfd7eecfec0c8e486529750b075e1d0ba03ff9621faacb4ae3c4f577f4128556000660df7bd0e687f0d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb645f2d19ef8d65b61041da0ae4cc04200e8113822782e8bcd9b82276caec3af17a8c4de3d340877c7731101f6ada069c290ffac250568c5f3096a62c7fd3ba91002e281643a5b9a795b9e84c4abef696520ae52;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd6d630c451fb0a8356524101a3d7e51b8045c7abacf24eb134ebf7e3ff5bb8e0824864c20d122e8abe21f579f26dade0a77195718f0b9f8ff28c60163e6ec5ee240b1e48bdc5e4db552d686a99fc62528726f22e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab3394227f4cf2253bdd3528f28024b1013570ce57763fe2a920ef2bec292cdbc62836b014f479395a62afb50d92d8e1516b9f5d0088bc6bfb04fdc5647ff27bb79b4de03bd38e12a3d955895c9e5c784478dedee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3eeec0e911d25e935c21e1266bec9f8dc512c533b6fe4e9d217c3825cfc5646996ea54bc10e1810b39c7050b72644253362a2985a8a4f5c5b2783d873a53511d5a5f0069314bb3189121dfab3c48e06223d282ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73ebf735e57d45d56660944ddf68336171a5be415b94605ed0bb0274489ba887d85b114446895509911e885da52c0560fb57ee28fdbd42d989cccc5308a9e5fae223dc8f4fff2c52441263d6a075b4370420f8357;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50c0612dc025b926f8bbd3103f70d92da529d0955f1ffd983d9c2f46fa879c459e604c0b9d476f5d7251197b16a6f73dd26de01ec93868e347e497a452cb2b349815e3069ac9872c160e321e4bc60cf4407bb30bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha45ddf1b5f8a292490121b046aa63999dc4757d9f1d8c8c31afaedcdcb3743ced97aeed03443d26be1f78bfd63b1dbd8869b1ecb9dd47ec412533ae4f4b0a1748137435db9b8600f4d4e8c619e9f9183977b13c30;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ac4ba3d9964f6e5dae60bc259b08e926ca607acda4232a0a63d7440c86ddcec7389153d899d9efa49a53ded5993f4400eb8d99cc754d2d418cf64a17607f5ecc95afdc8d656da7cae41c4ff8aa372880d28bedb8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b850cc2c27b3101f82b0c7e9c8ee5ad5a2cab5ca06f62d84921526df034c74337bee4b254a601af76abc670880e1e9ef73ccbf762912ef7a5e6057027f6767a10a81fbaee39a7e3e74c6affea5cfa2cbd1059f3d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1e50872fb3449ae2f1a28885c6a20e9252aae0f3f7be35f6d1b72962834e96ef9e8f9366509b67853a2134975843ac304a2aac42f9ba1adb2b910bfcf7b9bfca46d062e5ed3e86cf984b0cbc6651781ef791a7ea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46909bed306be161927ef51e99dac27473b96163d3ea9490b07cb6cb0e5221e7d0eafd75ea28c5867dee2733adf156ae1b89592045d2c5c20bd73d31414e967442f2acb143674b35a0026f7f59310c7720494862c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0bc98eb68152470b1f38a8f0e58cd9506ceefb15deebb88952f86e46b2bd150422d13b042cb87044d048263fe12b48a2107568438981dc47de957de5943047f5379ce6ed3f053a052ce7a939d2485e5c9d831449;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h355d0009ba33cf950ddf25194178c0a9f760fc2444d61b05631817c29c669d1e2f5aaa2a3fbf6a245805a971e50b86e614085bfb6e6dc54c8647aa6058a3af3e28c6f46d7eb24732b382ba6e415de495114593130;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e71b9363d3e09ae8c700d31497e2d7bb38875563fad6ac6c29e20700c4888dfa251c4eb2ecaf57b895ac2b036a04b85c68c5d14caf266b8e48313d1668c2054c496d3d1263acb55976ec46e5104d36fa6112003e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63ad47c5a90216b9b58a95c07e36fd9a1dcc509a992cc4e124074559553261b2f1d20521682c62fa840cd9ac08cd3b27d592f274c72184d21656909a61de76f437206720e9be27a55bf223a4a08900e6d92f6b8e1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78524c4b34cd112a3dfdd51e2047beb97e599cf0a59523eb6d8d0181611c4d1db7421b2363a2ad1f0d01c24bdedbd0d7a34fff845b87c151f946de3ad4d1db6f37abb79fc241ee57601ead1ed3c051b0ddb9739ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9d360e42b0a330d9e24b40088071df4955b1c1bdff2afaf61500676e8753df34248eaa5bfd3e3073f2e16e594d2be206e6bcb588f75fb14ecc2ec1138eef9dd8c271e9cee837dba0dab427eda10b6b6b122824a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78278df73e2bfd92de150f1aaef3daaadaf2e9c40b5bdc6e00dd57ffea985c0cc8ecb885114a3226d03be77505e5d00e00e2a951108765d7280f9d858bbfef496e6ecbc33a6ec8bea4d13595687f8a67b2ffeeb91;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heec1db997604869211f00730994b039950f0de52efb246989cf97506fefc7d26a783ce12d8dc2ceb641da334ff8b5a6826c218fcf035fbbec02e5ea2f6e1522ae7d93fd9f1edb8aef11957b22f2a5c15021c2ef0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdd1add2df1e65eab9bee4b5a7222355c0321d1e1cfd306b02e283a0bfbe304d002a76fac5441e733eafc2363753d46e585a17e0c317f135d1231805bff8a87b6beef2e595ead540112cb5df7f0a1383dd72092d4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b6acf9e363a8d67f2b725409dd1be07c8db342f33fbfedda2aa4bbda9b45e787d1cd867e1bbdb037e6d7795f5bd72127fd4c087a09181abd8d711d86e412707bff9cd92cff37fd555fdab4c47d2bee495ffe35ac;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha941f12d47fa3b3b44ab10640ada0191103c8ed1b852380bec1e30bc51048b1b7b5650e9b0ddc546fdff4edb900682db8710bc354bd9de8a062959b32b6e197dc42ee3b277a40af6bccd949aa6e8d03a4e721c83e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he86e6879d2a80a0e33d84d82d56be2d53ea2b95706a7c946487b8fd9f4b4e14bf09e39a47296b1f75795d621d9f25ef6a167da5fe8ed5d7a1892b01e819a73aea13f05e8a59217ac04fc3913dc12d63db9fd1d5db;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h585b273dd94fde720bfca02ac527897b90f67115706a10e53684b1f7a7011bbfdd4794ce8c5d7e374a07a086e5f9be059cf17141043bcff95763d56b71336ad597ce71604cd252449a3fab57d6c7ba75fe8f2fb5d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc29503517ed5ca1a40f278c82860525c99e28cfcb4c5fa3c0e7524c80dc2f25b4cda72c1cb494a5c2edc7531ffee967a0604f5a626e0ae5916c1ffe0b7beb63a873179ea5742a78ec3ab7078fd07b07029ea654d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55c2fdd360473be30a0db6fd9b9eadfd66cbb6b6243ede09757d5dfd0e5bf5f8a6fa71eacd23f717791177ee9093c877cbdbff4bedf4ac3a3dd98409b7a0e867aaf09f5e7d458ab1354ae077c27976c78b6272696;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5d197f0fc70019f0a954d9f4c875294f0460f6278f006f42b689e53aecb5ab4fedd588b086cb5e8290885a261f73569cf1c3e3981fd2e1de122ea84adeadef9b6944316ac0db9bb3e43337221c0210cdcfa89cfcd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h65e9be18f4079d21174ade523072d8c58b59fe2c804022d8e139b5feb1a11cf7be72e0348f145ccf0924d4a7894686f2dfd4d12ec5c88cff6a40bde9e4e0737537a8a78a82c2dab2d59291ead53dc3e11df6c0764;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha915798aab5b4cec9893083e6f06f76d138caa20ae5312c712e7b5ed9231660d97c61ae437db5a7c8959605f096315360e7ccaf04346674eb1b98311b3aa670d9f1f4bf7776e24f1bc7641e494c20c045d0a50c21;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd26464feb3ac80ce6bfcef5ab386b7e99c563cc4b9ac7871bbd15244ef2805369cb72870ffb1499ff1f0e0dc47b700b7fdfe3dd430a604db3b0fb51d2b6cbaf2d2879fc2efa75643f0f945fcaa08a6198fb6670c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d6e1506287ae54409dba5a5728402aaa3b50dde9ee9feb11aa6e1fb7aa478732e48d04d084bb35f788e373bc193e04bcd9030dd0805d01d4e4829cf5cedc114fe16991c57772db8c5f59a8a28fd6cc443cc51ed6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf54bf17a0fc4147f520c71acaad0c5b459c8f54a1b51f6635da91ba5eb0b845235c473485cc26173e1eb6684f324d54b50f096e968c7e65dac5a80588e3de3c785c8eef5d529ac97c373f02a98b70d7a4170986;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2186f0b0cf1406d63e36357d58362be830b66739740cfa480aad2614f187b0e7a24f0c23fa0bc28658352ac741e72c0f5ab230f7f72b52d6b8f18560ace2f57197fd254778a400ae2b292a7324442fc1aa798819;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd6886b525dc0c8bfff44067962e779d85afecb8c1d6edf6e7ac20c8d24c4ef7cf2bcb6d655b894a61be3ba2d530c61c13e876318b55498e700aa8c1410f4056eb350b690919c4343936483369579638935872c80;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f5159822b5fc455b4907daced2d23dae0b3a3ca2019aa3be33d1ba8a225cfcab6645c3fe95ee4bec75ea93a9765ea279e6405975dcbe384ed667419fce1d3406a488a5dcbe8b031fad798ac8979ca85e43910e53;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcff5e37a9ccbe7a329ce0a5b8fc1587651e2e9e0e2772ecffd613898267c150a974683a158c62c3b7b56a6ffc68f2fdfc34ca9377ea8e27422577de99536c7bd5b41eaa508e254e6a1312213ea270b8025711c4ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h556e3e763c2ca182edbd1935a2fc7988b92f27f7bab4eec45781cc58fb808187a0ec33da2dbbd4e1595a8b16683d9f5fbc17cd34a961b7e129aac25a0d231f257ffe86b1dc136abcdeb16d71215ee5c4cdfdc2bd9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9dfd7e843dc5d45c640b4a33cdc6254d1a5035a028d5f1feecabd24fba11b8fb0543bf8cea47772ddbe9799a64ad4ea79ec4ca8693dc1037b87aae2d66db593016adb8148bc58dcce335b27afc6414c1978602db2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h236364e740ede1391196f1908e1c9aa1d36b00802c4b4ff0687eb64a5fe0bb8c6444c8492955a1555d816bec63fd62a23dd69090ba8f8586ed96ab7009ed067b4fde5b29f94fce2ea59233be06b44ea7f25a4e293;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ecae6c08466573136d734c714eef70528184ad57477f86223f6748c975394aa95d82175d234921590342f6e33d6c803afb22817dc55df90b91d92b4dfe99bd5f3985d42d719d30dd7b3728737ce77b001fcaaa24;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb567d185bb0e6e75299537621b7b71fb857a91636a692d63f92c06ec3c8539796f3a331f1ea7c673339d046a7e846f8cafb3fb4c884acf2ce189e94a71a559949ad2ba00e2c83e378d265b0e26cbd33df5a9cca7c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3b850fb7718613a11a401b8ac967e6229729d8872359bd2021043ff82451311e0e14895fce9601e56b16f314ea02a20188b7a86eaa187c259d5dc31aa6673e7166c7fdf657b78982bb165cda82c7fad5100f0cc5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf61c3f342d5ae68224e7706c7c44a1664483aea4ac8a8d7644dbb3854da7dfc4294b8168e5b78a8bd0b8b1ca4164360c2f8463705b8e80516738935db45d3356a72b57f42088b4ed55100d629d989dba9ac4d8d07;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc42be4403ecbca7db1a65a0110160b9f617f5fb2c0855fc19bd1483647b4be4d1b691ac5fe92bbef48bd3d67a15c5bf6bd4d338f293bbd15513dbad2378445bf5ad83fb81809c16396c8ede0c373b733e1a46ff7d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4d07285502c5d5102f4680746a409d9abfa85cf37af49c129ee8260001134e06fc64bb44baf2e258db3c0f7b72b145118d1c8de00a765f7010a6868db421de821d11200ef185c6a3af649c83cd0692c49dc1e5b84;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37b2367f8f1439acb78dee630b0883d33b3dd1ad2a08794d5d75d1d09c5ab23cbb079c6131d8163d671153fd08e604f8d7c8269a1300dc61a6f5a7fe541eafedaede6326ae05e037eb48f634d0366150b0d335d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c79cd31023c8fd190fe6be42794d27fc0d3d9082e03edc538d35298d88bff17169adf28112f594869b99b907374b1b43692ab57d9becbebc4af411fa4a69d9335dc9ae0caf08296beae33430692c1d49ee87d4a8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5223a745af8704928afedd9790f8fde6b85591fb56a9d9f44e935bd857d133ff5408a7dce75efd6722f3463dacc48766e19b5a0816a3f0f2999167edf001ba6ab3b41ea76e1c290f54b7ff98996c63566f5d1ea85;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f9f956f4546e27058970aeb478b853c1f028aa6667c0ec9fbe2d7b57a9fc6d8c15f5e2e37ea607b9b7f62f5dafe15cda1bd634eba475d8db54416dc613b3cb898267f3f568db61e70260eba7ff663b15a66ba407;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h45c3ae8a8f3f4cf414e543bf5818fdc3e553cacb5ad9a8d8ba2c15ef2bae11d8ffea10c4be0ee0bf81f630abe2e6c758027561aea7e71b3ed771ca09d86afb4a34743718bd5b010f8dfe55082f1b3175783663532;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2b148b4149659c21591cfc29f3642751f949db6919a2c43b6d5cfdde5f7f575b92671808ed96343e4d6961cd1e48dbb0cab8d576cb9f6b79161cf1c01566bf5026d96dea8bd657c89ff9ddb70c8c4cdf87805ee3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f39d6c8fdc20ceb92028a7ddecc2b4e7eafa08251d2341d3489986fe08795d417be087f63f6c12357c6c9e67edd0e0cd7bd589c95e2f810d8ad72abfeb9ad3f95ee9deb9f1a31bf955218bf0fed5f4d04f76e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83268ca7171760cb95b90bc999710a7323f66c39226e041dd96ead359887ba23f82bb1f6ea977771cf096fb6e9d00cee342cd45f9b7d1c70d8302af89439ed031155eafe6ef3e275c726ba7664a60e7a15f3201fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h944dc51742c1b419a03e24afb9ac392ec7ad0ca9d1718486bd9197431ed7d978fc1a42eec5a5147f4976fa3abdfacea5035cc874ae2f4ac8c02c2266dba864526b74514a054d0ac7b9c96ee882295d80f529b87f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb09ce8143668f4d08689379c2c58847c66925628096aeffbabac09e4c00167c77574c285fc0021ec5817515790f87251af0ebdbce1ac6e965e8f88b347e805965729c852dba59566a1402e0ac769debed0bb4004;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc34defede428686f7799acdfdc37e77ab335d9cb5c6fbe3ffef9a94c7f30314c34573333837dcc438d7e94f7456e763f3fbdcd9bb7f3a90a743b26cc1a525e8fe2de4eea5dedd1e5f2cbeca6eecadeafd7a27b09;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4f9aa15143acd46d5250cfcac62c14c50653370f32392c852006a0b15239deddf1265b7c1fbf4adc286ec5fb0600985f3a7bdf3e53259de88ea2b68d7e43b2517d733d5d2d6332ab04676eabaac88cb2cf587f84;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5940ff3465e1ef6529872399c57562675ea7e02c93e51e51d4a2ec5d56c4688d6dca33e62f52d86ec0b4617cac5f8affa5c1ae974f71e684da284c75644e5387976a4f7c2c62acba102c8dc497745c091d1778ba0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb35964851ba28d2b646e81e883ed4a94e3d70247e61455493eb4305a51c1b0d48b46a753ae847e9826f948b23283d87e02a79644c1f1a914e2367f7d4d2425526888cdf1e514c6a1afd8dcaddc49e1789a686846;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c53d45cec592eeef9ea34523216d812765f748b177963771fbdbdbcc9077785047127351e5e7d2b4ec6fe6ed909f4bd7c8c6ec4b5ffc58787b0c6b63518d322bcaea34e9a719a582023ada003df03b826fc16408;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8159a2d396a677f117f880bc02168f756642d6d26397649fa0ac06374bc4fc61df645421db12ee5d0dfda18841e9f55f590d62519654f1e2098d7f53a6c347ca6d23afea1dbb7d9c70fc88554aaba19f32a7d264;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88b705f02bddef628425c15ddede05cab9950f1d74c66c5c719a663c7324f9a54e74f29fc1c514d2e79a884ebf269c27b98428744eef4683b84915adf2a51724a14ac224a8ce4b4b269c5ba98aaf6213a42627aab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h31962424e5248e72107f746d1e5937c0b4fca23508ad60358bd8c9d424bd72a63001aa11d7248e95cbd89962bebf40c0dd76121762c50d7efc54ee9d811d1c46259e9e3716d5a08e6c43ec9c1b5be3544fd159ffa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb49ebf06dda1b8aa8083f6fdf3ab24d7fa1798e37683e634d270100aa091852cc53ad00fd2ab1e2382a69efc3f8dbdb3c019695bcc3c38429f1d732acb842bb8f536ba58755d5e853dbaac3fb45a1a532ea4f27a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4660673634eac485b784518523f7667c2bc9815d2c031dd942f33ea696479169ab1c0b8ec3842f68e7e0df9fdad78def6b6553d4edd0ad54778157d1eb8ce3634e842580e8e658a1dace83a6fbd0c004e5ccf2dc6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h975d802fbc13d1d7f68d1eeb9a4926a05c1872ca7e9e0a516e7f4ccea2edd274582c97d2eb2554144336a8a06ebe61db147aea345d3f0cf82db8e0f25f46ac2137060ae4fd95a4e6ac55d464568c6568415cc6e2d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbf10790fd9d2ebac23548394e075d671893096055fedba11428fd439f5afc2229bdd45640adad0bc164c196495a0370867354826ff47a44e5cdfe5d1805897529127d1612836ba171ddf060f5153830d34b4d20da;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7f126c5605a1c468003f876df01b1aeb1c5973b67934b9f1697c207a6a94605398ceb9269ee9646d82dfec55c546fb82c27b1ce0eda73babe547a563136b153b6ec7d454ed212df88955bab95399b0001c010a75;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41ab24eb17eb004ec98496d0df41688b1ef7f0da9d42b3cb13f0abe202de1a280136ebc22d7805904c369d453c5815797458d5ea3d364b908fde36a684c31d0610e65390a81943eedbdb1189a2b1549ba31651ef0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e9980e7f1703ceb6fb694d00528f5fb5a7f0813b8aa107ec34246011607e2fea6a9fa176c1d92b93546522aba42b22b8c0090395644d57702f5a4e726a43f00a6aa75dd54f6504bb6cff2594fb6d4cebed1bcda;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha22510f4721f23d2b70ef74ba04776a6174c7b14ce7a1e1cfd59ff21df79c59e792710751c6711d1a2207da8d5bab8d2490bbdb619aa3416fdf09adf9d7bfba18ffe9ef9b4d58dde7eb10a3ddc7600e84f54b0ea9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd23e8f11ab3c092a7eccc28dd9fbefd56def2e17f5fdb44ebd5036a9698e9dda2880955c5a8b1e4cd00b214f739893bb986c4614182dc1534b876e538bbae76d25194586b64a6bc8b055e68f85f4ca7eaff02c43;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb14e379d9feb3557e2fbaeb3e108c70cffe5541a3aba4f3644794b6784662b3ee152f9ab2571f2392c402b2ebb9f8833f4581a06c4456da6f1d22e7c4eb12f791430b8aa8628986a96ca5a4b00430a1f518e73525;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h929428b5b9f2803b1e5d87afd611684e294f1acf8ceee929b224942adc5e0b8fb9119c64c2fedb3cc5b534945722c27d7f425604f7c45cc413af13799ef51d7cd91101c4860ce68f41221378082cc493e79bc3b54;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1a9955957128b17647e31b221253bfea0335b95b5ee56626afa9b3743fd8ef4f079a87b2e62a404309abb0b399c2dd392eb36bd8175f5bc78be6d6079c8f26ac1c371a1dee38efbb2e6e94b28b9797d8ab2569d4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h331f9009adb5b208fbb8ebc552adb7a87c7546158b625fdb12952120e25489e43b1f45c241c998ca8604995986e15d7ef081ffb12466cf4e2ce8cc4041f775cf86a83e94fd9433cafd4e5db90e6a70381c25e7e9d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0826caa93c8926cb22c1ff1f3909a4cc9c37b384b1a8a9729e1ab38767745e2d230375963090cca46b168672b7684ee95d8b1438fbf35bc2c729c19f427764bc0d0e38c384691823eb5d79f3fea34627a2d2e2a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f4ea85d771796431b8c97168b99a47fa4fc0bd7870d678c1bb371681b76d2471d590fe77fdfd8a3d5c5f4ab205076b14c169f7cafb38e79a9a72037d2540c9370eccf93db899318fce8fa45ad60a515d39ef8f05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e72917752b1ff1e569383ec3aa3a0ed5ce179f84cfed347eeede62238e5d282f01ca36741ef40d0c3a537470ca46c348553703d44e98049b1e72d8a399de4c86fabee37b5571b003a5702fdc0f158ab5fec02602;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h948ebd9e4b45372640069696c1e9bef196e5e5ccc560e5b67e9eaa56d75c68ea6ab495c75945b26ca9d1f32ad0af0810ebe69a6a3ed03f556eb4cdec5e0e7c729ae7882a7e159de6d2c7161194b46083f02ed6ff5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5342bf485bb8a679f8d8a1a82aad631728abcb68a1b021a4a4201d22ab7697136545defec8e83648797a2e9bded7437b01025af7c5cc4dde6a044a3886d15fb642607b48e91fedb0decec1a36a331473ef510e16b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58e8f786675b6e1958ac86acd0b441109aea585aeb8a0a75088c5df5e2678e93e0e23fe8df8c52f611d0fcd72f9e815356a58f06602e6f48ed759139da19e5241412c65d06ac65197e2ae73de8e60c2980ceb3ca3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h89cc0b955c1a27cfef20bc3efdb221693309ad6afabe34a7a0d5c899750fc7ca17debf1cfd94b043fac5e8c9e577d3ff61d547542bbd4afedef5a03d8a87fa48857786e86459550d6d0f672dc6841418d5b7294f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6f0113e9c0965df57153b8b1aadce0c9ec400c7780f5ece6813f3d6d126b3b030477a7e5a5989e5102d349756b4d935ba730bb9b09545362509f718894a2ded782a8de039317b5d95750a5018020c4d9362c533b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2921cbc9478840e3ee0efd582ad7d970e8d56bc14472aabc6dee0be0f737b5f7a22f4fbe090181570ee062a7f3b722c962ab575616be1b5a321476d2a396fef51025bf6f008f21cb6a9588cfda85ed40578b5422f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85019713537b94d5e0cefd0b0dde2dfef520b11b4f23ba2aae9628b076a8d4d3f6c983e5f608069a21416c666f72aa99e8b13bd5725bdfe0acc700ce1af54107de9fbd7c2d974bf398b23c2a4b8fcefa2589012c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha80c63c53cd8f57dbbdd748866d81ce480491be5cfe91c6fb4dad4719d31cc2d1dc10d145516717665f7ae95fb2e59ce0651bb56a5bf3556924a29fb24abcdd6489ef0654e1adadd82878fca4f45a5eeef0826d0a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8d9f92be8be90b8de5dfa3ff024349d6edc1f9431f1b3c3146b89f0e8ffd70a6b0e86062ff3f2226954981abbf9e39adc1dce78b2704d0bea2cbd82c399037a564bb43a0744684fb4966a23c314fa5463322136b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24c1f79ede48bb3c78c9f4a1751ec3a1405672dcd846df19b60eb83741ffc1e3e5af8b988fac56e4923af63c478a3dcc3754a516e74ce9d6261061c72b21439165055d61140ae7ac9d32dc2b18922f7ba13f6d1d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43cec321fd36329f5c4c9c397c357dee270f74c9c89b4b9fb2e6b8b5f7d4e9a951ae681323baf23cc366266be4ff662df48c108e6e75fd08ea88e545b95cd0404fe58de6594b6399317657f4d095733dbc6267e73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8112ba69133581e2baa2a0318f06f08dd4f39a280e4198a51db4620ae1e94cd8f2b33bbc265901841c58742998c105394065f5261e33f97607c2586ddc9f76a1b7a47ab344dd0de39df0a8cc0718f950372ffa7df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb0fdfb84448c740e53d3a7c9e50f6682a6ea3927ea9cb8668233adc51a4d41f37042dff75bed26d0169870ac4a23f80230a45433d165657d66a95352f14bc26b93a7515ec3545a99d755669dde9a46fa40bbc35ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hebf2c2910303485dc388165b4dff764c06ae08008f6654dfc1a82b4db9c2c4b29714ba84ae1159398c474a37aa6734017a1224e07e95a8619f70130cc8c01b000f74ecf7c922f6a35101c71ddaa8925fef3309a91;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd294bf8f3e95a1b5889abcef5e4dc4dd14910a03a2bf37e17d9efce2555a7c64db1b1e9ddf2ca70ddd6f18714d68fd488359a0f2bb3eb60e02eecb204b4f0f4a5e3cf0374edfe5ca03597cc8143a786bd0019f688;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54ec540a5908126982481dc7b57eee065a3e83dcc14e998fe4259d4d7bd41c3b0c89b4ebba95e2f7323e468e32d87c8c939d26f139fc862df4a3ed81e981935b49ef79cf4f55dc5b5c32637fb7964c9c0ee7e8bbd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h211624261c431a0585812d3f5be74d260c953ade6f643a481de759d9aee28279a1aaf8168ea60855c841b6e71790dd5e2a21fd53bc520846e8b54fe1352b16daf8698f9c9073e578eb20acd62c7b31395f3e302fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h609816a5aef12f0ad8070fb32171a13ef2d1ec5128540915dbaed5dbcd266387742ffee0d081c426ca69d8ce040557047fd53960276fa2a078ae972768e8e051930729f049a3928e0d33bee665df4f1ed3d9dd96b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h267c9a0a138554654b4fb090100773a00a4dea1f032fe9965df996d287bcfb79d4b941aaaa980d0798d73988d81e579ad58646a66a4afd3c10a54009fbf151cbd0ea6f02fbdd0b239444ef995f488911248569ae3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haaa327f66a1cb8d3193917cdd7a15c7985c894f611b53d1d8406dcfd6aeb4bb6f87ae42e87563b8211777ae537de37d5447b58d28ad58a3d1449753692b88781046816cd5eb7cdb7ced0926d1df469130f3f4b0a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9bf1c6676db31677fc8e2dc3e9336ea75368e0f0292ec6c51e733062d60035232ce567fbc51fa08ee6d8dcb17c6fe6613a96e40140a352b14ea51e6b2939587c11e8e1e5a669fe6a121f42860f5d891237c068549;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd042f1a00de3ad2387a906fc7092af2b7d037a797e49b832b65d01af8b8f545b348ec6f6ef917afb2c40a5064ba2d3a80709f3a4dd7272c22e92393aad04453f0e534caeb8c9e2f89070c39770acbae4c4a1534a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb30717a6cb1b0eece9444baa017f5c4923479754eed904743f78cb5a3bef7c7535865ec3f2eb24b86c463ef7a3a7e7b3f96e2a8247e215d0372611d38b684b21a1cb928fc0e0354655a129c6416dbd2302ddbb1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hde1aee0fdffcd422ad5542ae7062b8830313eaff321f0e90b947941fd603ad94f82419b180f3ab20d0488bb7a3b56014c07accb1c0ce35568eca21f4ff81d086e599a64042c3fc3b7d625a5e330b57ebafae8914c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc71fdcb1d005011dac83a9177de46667668760bc2182906fe911d56a54a57b94e5c97c4e985a3102d771f9e274201524b9ff8a74626a5dcfded350008f8aedb29230f9a5c57bc56e86aa616f0af1b0c39bb5a2706;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h167a041f8b6f942539d2ac708201603bdcf058501f1c46e525441ebb370f8900f27581e68ffc2757f57680ef5ca7aa1d18197fd0da36bdf4f8c15047e0294fce26414a765c686f6413bcda4af15ebc5bd8eea7249;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2da5b5360ac8adf1aac341140e419fe04d9755ade15d178c187e70093c8b50cd3b9fa5f900921d427d95f4ab7fd689f59a55112c6ca939c81d65fd17b8f2256a23a095a4702d9b29e0922f3e9d7c376c56d0d83f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9006a8392c14b5b7398600fe42ad894bfc9bbab2ec3a4f6ba83a57cc38cbab97f50d8d0a00998888258b3278a5cb8fb59f0d43dd2a3f00999fffc57cf423510715710fd32954e429dd5cc84cd3054ce52d9a07457;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35f187d4c432aefbf56004e94aa30f65e11c9d67ed8268f574c929c19d097084eb5a74805b44480219a7c00ac29087e903184dbe1ce35d7b437ef863eecac29e4ee46eb28e4d1ea046380e2e42a8b925a72c76567;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h13caa79eaace329895992db5db5eeec0f2e78c461f97573fd33239b2d1c79283944990f93cf575fd40cf52d3f47d1255cedcfdc9715b8fe7de393926522bb549b4f699ff7f9874f08b523f505865bdf47cc292414;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9063f449fe64f6e2421247906e579d283feb3ab02c85ca02eed090934de82d53a942ff9b60e37be8cf5ce949452de78b0e88680537b9bc3587737c32b25111b065c9066a0666f54f1fd18955d885eb90361fd9378;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7000282913f0f3e6b7a2c36ff5e2a8ba0aefb383fff6ba02a1dd0cbc09b20ca7d2bf1262beaea40c6f3122df40c32e027115968e5172ca47157d0b6784d5f9f834b76e4569cf53079c6f58c0a3453e24473aca739;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6cfdf734ceb99849725905b557587ce6878de2833986f20358e96c25987b44dbbca4fb8ce26385cc251f2ac06ad6fe411fbc7102a7df9eec50abd81676e9e8f9c84f2c9967023118a05c21beb81bc3744b1bd0763;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdb287181b9e5accf27cb391a99eaa03a688e16ccc6eb057392636ea255d4664f8ba305effdd24e52a595df533b53c8a0b0e975970b760f6d2697050775c3fc0548cce385ffb8a1375262d9e055b26cdd5f2a54c4b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha332c150bead7a0598051d077f83c7ebda0b45b26da534dc381a5fdfcb1d2ef606b2e750495362841535d4f96ab60eed685eef38e75b54d6a300673dffe6b5550189d68bb14fa603ad2325aa83e93fb4c0a6c6a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46fe15fa7606f00d88ae95a7b065cf918a8e1da731992bd68774defc2f7c21bd944ccf9b48fcbe61388f17b4a97e233c69a8256adb9d63d066292f02d691bfeafd4567dda471ac107366735c94cb288cbd3ddc334;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e99ee834f422fac9824b52a0b8eb1f53cf70258ac837161f042a6c8c6abd3550db7e01fcace43c315c91b7fdbc724b9924f02aaba59dc8c3d2af4aec41f4c23bf949045d1e521d8d5eaa9ed0d7aca28cbb0d4b7f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9fead32d3c79e1689025965ee5b35fb8c32fed31f3e94c4c438388235c629b599f9f1957eae88c956ba988fdd385baac18ed027bc49fd8305e1f40d7e260a79ea2ccbfec45b2ee836bcfc63101f59c1587dfef7df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h931b0d54176bb328fbd924bf4cb32f80a199e7835c43320ee5abb8a2ac0397fa8427daee243f62260d31d3edb753890358cae993d10cfd7bbe4c2bb10b216af31441afdb10dc2ad6f98cbde49053ddb244fb32f5a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa5f39bb9ec4b90d09773ae5e96ad844bc9081d9cc35a40ce73fc60dda88cf873f5db1bd66e32a3cca9d169739c7b8210454d35a58c9d964716d342cdca07631b7455072c2a61cf9a1e0aa5e4dbabfbeeaaf94dd4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5aa6391560e8177945c1ab16de904b7f07356acd3d47d45a1703c840d502eff43856e998334df633ee5449b0c2361bf91c3e567ff9752dd80d97b5fae3a388df9aab001fa1a4ff91c7009ba43b1c56e5b39f4c4b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1506c6294eda121956169ff16bf22167952f8d3bb792a6336e2f83162e1a0e4e6a81a93e94129d9b153c20d4bae4208927c645237b168b5c4bde1b5582d93829e7a815b263ef8568d860768137777450a5c39cfc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h691a4d4bd198ec58efd1ddcb8dbce587f761105e3477d37faa096e849a40b2a95ba2b3a40de4d27433607c044559baa1dfe452d5655b56b2a22a536d85be918457213b7c028a6de152c092016aa5dc8f9b0b0cb34;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1dbba6669a706e5a10c42c6630a5a80f23b4e68fa581ebe9e4e47bf75200eb972446446bba361b034905e1ca9f3b7339c6f271b0eccdb878427c5b5ddd734a9e14a3bc21b502d6a48a9495df40c8598b8097c504;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc8680080546f0b0dd973541f2cf8f568effe5a47fef9714a9a646ac14aaa724e1150a046388ba00b6b968f5fce3328b364b4da2c4009104b77a86e33e73da5eaa91320f8381cb6e4985a7f0cd4dc57acec8f4c70;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7080e9cdf8a323e27a7c3ef96e657e6ab706b1e1604a16578e19c61715a0c05a152701a31eceae1ed56a5f1c056de39a27f5446724deb8c1186eb33e7b5915d121b1af20ed6916c9b7f3041ebaa55a96a3454995;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcfcf4b5f48123f921e17bba6257cef55edb4610efbb6cc6ed5df99dcbddc84c9d36c0bbffff01628139ecc8cbb6dbe558d9dce780aa921125ad82c3a38309d1780a90fe755ca5c753c2c896b2849fb8dad4d1fce7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h196b936626100df0d6a8019fbef7dd102ceb8fec4ba34c62eed114a62b93ee011cbeea994756ca669ebd1338fafc7f250531c6969bd6097bce2da88c6557dbf5f0d29616000ccaf12802f617f22cf4d2d241f766a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc4079e87600ae4800f398c5282640567fc01f5ba75e7de7dfb0f6f92c8621237acc7f9f73bdea67c1233375c93ae7b1ff115dc1f4270a1650c822d5672f805d37f6c2d5694e77802d8b15d1f126cb5ba390541bcc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f8e99b490ff38216b6148f5b960213dac42c2bdbc54b71c8bbc5002b80fd0b358716daaf320454b3e1099e66ec8501518fd6864395eecae237b278ac39dd339b7da2a712f30cfe68769e4f90ea278bafd5cc9c94;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h209cc4ea226cae60f11608f683baeaaf12d33a648abf16f0173f53adb013869d17f194bbdbc5f390193aff9f780805ddbb762f05677a4cef315487eb9bc2c241390113adaaa46c51f155b8e785d372e2a00e67c39;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdaadb7106ad65fac87961df88c0b954af6c90d3cd08e30d36a73e5cfff0eceeafd628439b9ec318ab1301c40397eff4c935d9ae970ea60a92b12b3692d176d22dca2463e3c37794d5bbf8cbb7139e4d4788c5bb09;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h484cca5b16d15046856df7eb9d5bb7d8fc0a6ff6937aec86584f0c056d901fb15fdff5d6e832003ec30eda91f00ddc9a7bc85a102d2d0250f6ac2bd566ecf62cb871e9ce03bf009f1c36188c4b0ae591e954e7136;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72e8079eba42caa6de244b7727af32e1e027dd7220e345c813c4ed05bc3b1f760557260a61ef318cfcf46cf40d20288f11da939255256f966227216693df1288b173e3525439910b0aa16184d9aa06c883c43ce16;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h966533fe94172073838825d591940ca9fb21a3db4c697b63352f2faefe52a669e3f1b27bcd70235927f63327ede2ecfebf78abf791f9bf15f518bff87bd7db5a6a0db9e9eae9d492939e70b204e13d3e40c76b8e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9146e4d1ce571730574e0b07bc370769efeea7072907ff1f2ea2ff6b9a5030cf9300f110be5890d8b9bd1f394fd9773520c65e437bd829a2f9578ae6b101aa4a3993458771ce666e67a587c2f64aafd1aa5354cef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h79679a44de7060064f89b0adda171a18ad72a2fe644e066db783176aae823d9468fad9f9a7b19e86482e29993f969f5385817cd93acb7926ac47388e2086facc5c62d588bb8bfa94aa605f797b21d6721d50c1946;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b52cbb86a9abcb1fbf8af8b01d124f551b6cc64bc693702917f3af922f6ce9a1bb5f43e0b7c4b425f0685aa62768e09733765d66dd6c214b159b7099b257fc2eb6f0f407c708c7648c3283c157972d33403cec5d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac8bb08efe3c888c8d285df55b7f1c3ee40b9fb8a4b9b15542c537ddbc2105b3bae43a0761eef3a17852c49ae7db0ee707a2c0ed12dc3ce09f2cfe992e81327b37dfa6d7a348e70133eb3d2e1d61197eb6d05de2b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd55a8957e546b7f7ec3fa6a1b651c24b1e3569bdb0abb2fedfc4b53f1cf08250399bd7367e2ead2325f2b25864ee553774110944393b73389b4e10254f78c2142094b25c9ce0cf4b219688db4b6fd570c8d015c9c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1e7a594096f90d667d7b4b9b3c72d24c90dc9183e18ffedcd6b7e34e465dedfbeb7e18a2cfc54744f178fb1d14f8b574c22b05d8444a8aaca77c27d83b267b035989d6b09c990b84927b0877f3b12ff8cabba870;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4726d681cf26e3368cc2943ae872a46a2d1c7c1f714bf92817d1a02106fc57607b5717f256b984355bb13385a6025cb97fa72a22f208b1a49350dcc742204c3a39aa5a892be7fccefa0f00d41c1d9657a69220c05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h800a4209032b2e4afad0cc626f1a4444640fc4ce31f63ec6cbbcfff4bebfc3414529258f7142d964103067f0a855f6169af51ef7db18a72943101529c9b489d077d361960d01d77c996b1db4de9d51a8f82d7e395;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b034efc9515bb122d7212a906386f0bfc43625b26b26a195a0de0cdf59a853a676c633af0bebb09533daa2524d7d49232a0fe12343ac6204ce3b00dfdde7da13161004ec3eb59d8616b1b454c64386ad22c8f612;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59720788af07881cfa02e23822a26ca173ef2cbb93d97d54d5c4fadf06897b1d546a93396bfc942d3ce575740343d964445655fe0dfae6f799aad6982daafa268f55155f51b280a5192c225f648c96f1d997321ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7c5a49f05cf22a245c9d71fb86869cc098c89d163b49e98b79df69f7042bef1807f6fcd49beb565305f457d99ca2b4e7013c6f7946eaae2467677c7fbb2462ff3be0e360d6dc0ba5d7b05b06405084bcd780495d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf853a315a1e9f1613bb4c535dcc606214ba00757376126a08111efe626b17d03c9b16905144a346c78fc3f37ab260d26b6908fcd07f1d1aea1b360e4096818d4154f46abe6973a174099cddec5a24bfbc4cd7043;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h757d7062a81daaebc280ee7a2c978dfffab86686eb91ce58055743cf800abf25c45f42903a0a4f4d752c61f38ab51d60f51d20249ce564573849bad9c859a631e612b169f6db8020cac543a43e68a879798e21b82;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbbeefaff28b415331dc2026339b8286db6dcc220e5b858ea145d663841aa15c9500bdf6142ef175aad7bfc6b0d94ffa0f7905013b251200f4bd9827c47ec1dde0506faf31707258f883ffe889d0ac43cef20e7812;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h499d1339a479fe29f8fca38597b8de90cd398e73c3e55dc9287ee1bb8888828378b2455b615193183f22b67aff75ee7d9b79fc999fe979933e0d273f63fca1f930db8f5743efaa51cb77a91b8ea948f5ca6d91bd0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd35720032c52ae11b7ab60f8cf549b2e35729d093631f16ced11c922791f4f962abf261c833d7a2f6db27389c793a7f3f34704d8ff90f08ae4343cb654e164ac4aea6bbd78d9bd7aa04216fd0876033b7d3634dc3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7f0ff695f93aecb435cc5180b8d2ad9bd442582c8fbc8358aa0c8ed7e8e0783456e9849bf2f5302cc705f232b224d4e1618a17cebe4dd8c7316dacf8bfe463d78b9be52ab8152e32c771e7a2fd6406d06fc65464;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h702b1270aa0a17ad27b83535e8de483195ac1a31bee1dff5895c4e8976d330ad91ac22d2cd969f27b5873aacec9138fb05d887491ee483f16df419f36fd26699caa7c08679248fd018b81ac3ad85bb1d71b932b42;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h528f21aa55112d35cfdf5e146016e873095d6eac0921c39e3d8be7cd90213146ae1d1247c702bb3cfd6363486c3f906de841b1fc09bc286f088a7d57b6fa2784c12fb8fd668144f3f074ce5d6800b7e18250e7054;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b4c3b01cfccb5039b4b8798edd6034bc3ec558ab454b134c4e55c23384ea72bfe3d1baa602ef54711b1d43a8db02c652f68d46fa4a48d0248b1e2066909ea5c40583d1120ff912997208f0ac6f2514d262baf30d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h956ffff28a54b710093ba0b4968cb6a257b89e89e1574e96a5768187cf46c97eb38bee5a698663fca3876543b40bb1deec86bd934d24b2f7b3a584b5f7af740f6b93aee0905c985d81a3afe2abc01d5b0b25a92f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h148724564818b39107b936179612729e352bc6a5bf1e445e5ea7ce10e63e94e3df617ce09c73f63b2c2a14326f085afd7d50ca2ea16b69b0876ae519a9dbd82a9c12231ea7f4b80964b055983795a5ff8ecf9146f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h40735f075436fb9b6009a4d774bd3ee02cdd6601e2978c7a21619c66f606563800b48cc7dd2a6fe384e17af136f0860647d5eb03a4a7e561287d451b311efb8cbbe419dafe019cf887444e36dae0c9d25cd186504;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hec7ed409d299582d56eec69ce5e20cc683e3ce5f0eda5d92041d1694744960260ae595c50dd17d7dc972537499284f1eee89ec53a045d35f2a1283b6245cff7d674c62f3e026445d5b418a723e8782a1baefde01d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h633afc79be5a5f000436bdb2945f98cbe3baacb42e431165674a464aa511b3b21aff5b5c503196134c9d74e1d64c8db1626e754e4a1208d859e53031b9cea654ebb273127b32b7665ee87845f8ee5870c417fdd8f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52e0e4c255da9fcff0e5ce70595293d6ad3657b69603924c32923e4622257e60335fe11f2440de68720f5f2b3ec274bf363fa74e11aad2e011fd136ba504d20d4794aa805932279bad746f4ad60ebe4db05789a4b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd8e2185d9bc1f4f7a5456cb718b8d02fb1c9de5ae92ab7608a7670e9c19776af92a40e5f3c9233ea95f71ebf612d36fa0def31f48cd78593e415a6311ddaaecb17973bc2fe62564fb7bf798dadfcc4e63b7bd2c33;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f1dca13fc77e1d515656ab7a1659c60b60208b8493b55df539611c9534948c2343ec80ccc0855f7f6c617309a701f750cfd349e5aa64d4609094385b876519acd39160510cdd720e2a2e3ab3a584060a7aad2e2c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd18c80c1fb17a02eb7e5586649d2cef63c3a3265c15d51f3b49fe5a4a75ce202c585fa1e1c009c95983b7d6109be3c927f2d97c0bf827aa52696531687b895ae8b396d4dda9cc7caab214aa100b06c5706c864ebd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbe22f0708652d4c2b0f661917e2eebe5700ade1cea650f93f29bca24559bdaa657f9cf0ec55bfc740e254de5611eb2406c27d7bc1c146c94187299711f52beb49336d4cdc13d2c36c138745f59340e579bc5a0f1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba2b0812f844c4809a34aa6dcf3faba0a5df680ad4c857eed086335490f3bf6681fd7d6517b17b97e6a92e92ba3b196034130f059b0d2fd112e655251e88c2de66fbdfffa287ce41c7ac95f44d5e72957bb151715;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h597a17e09bebd165df50097f076eb5e4b5e88be24612ff61517f114ee1cca832a586edf8ac241551c2b923a203a9bdb71e34a81a740c61ce6d0eabca38706b45f11ef57d17dee0db40f507b2924996e18b23ed412;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0c1d8d1f498685d173479245752f27fefcd2ee2aad36e6d5cf99ed4feecc4ffc0cffad566ddec3d34578f4d914fd547b684f9888a5e59dcbbee1a1e450e04c566862ed42d615af30feafb337b5a3d532639a7c2a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcd847af6568524c89bcad9607672ca80bc56671a0df65f7ff7553944b2e6d29ce4aa64439756456aefc83f24bc573bb180e1ed4e0f1c892cdb02aa2d1b37e5fe4c7361305402487f8bd53c19026d1c7485fc63ae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5ceab4597c380d25fef347415b311fea7fe941e9f4977e7055c6e314bfcd0bd7dc3c7dfc386c9fe135165017e4f248bc877e0d9f8d10b45489bf54e004e83bad612b1e928306c35a049b59960530f430c64e56404;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc467b2bf885ac409109885cc87b4f9bbf536436f72990f5306f3f548cb50f5e9f3249512a853954cfff61c164639d74029a731bd96e738d3b7bdb4492e5169b23e78d581353693c6ac1db18875c96ec66bd16567d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71d89de86ebba5ee489c90eda634d815d59498938e7afa1be5a7df456c975fd951109737708d8cdabc1a10c326598f9a85586c4797a39225a865f31b402c6537a8319edcc0696cc7581cf28f04dff64eabc7cc5bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb7bb80eb8a476b7688e215a078eb9814cb09d85d84482d2f12a8d83ee6355c2f6e54033102c138f5f31fb20df8b499e4176850b1d275a0ca623751e90b62597eb095a7dbe05348ba3f3351388f4a3a4c9355bd4e3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb95e95a395f2343bdbc278cc2c47a019e325bb078b99891d9dd900b82dd03da27b2a5fed8e43e28a5fb9814b4db35a8bee9dedc970152b82281152b3b039c1ef1419aa8576e5766f9d8b63ba949b38ba8cd5734a7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2574b6caaf88014556e78696a11df520556e12bbf0664e4f1077f5a34c6e609ec02518383d4948662d3216fe67751930b48823a56997b8decca635b90fe8edd117949ba0a204eab9b1f9b95a7744dd16265384e55;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h687d1588d73fd3d10bfeec320af3297be448f2f7917c822290d0b4afa0285f887eda5c289cdf8c994ab2fb14376dc4964746294493f1afd1ad45000a8cdd64c5d2145c2503cc743d8473613df33842d12420445b8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had9f16182dbc171da01722b5466637b73cde2b444b9816d8a9a19f784f038551b7806d1d2f86a5760c8b6ddd0a2719835ff948144d71d0e9b3d23b70dd6b6cdcd78d8051503b1c43211d1a23b5f93fb743ab39906;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8890f50db8be0554325a978139ce2186f02a4e268d9daf83a610dd958cabde893cf31ad98df95ba929ae3956ce2f703e12bea3ee594068e99fcb192dcd050d6c6f5fe559da57bf62c7e76d03d924e8aae75f973b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf9fc40d98dd8f83da64fd34ccafe0141b6348bae333920966d5e41c89e8dd54b388329c9a8ebce69f649f2dfc053ae69ed24ff12dfe7697784bcff15797023956a51d8077b33d025bed75e0b5201d076abcd9a487;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h249e91335b9c3d3a0050ac8c10e82c52f80a4039ed6726c11e42f7247ff7147ed1e2eba2e786f4eb3540d57fb27dac4ef303b4cdc8401decacc94bed091880daa45195dd56f8e3f0d4b582286a29af5f3777cf7d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d8ce6e3d6cae0dd836a0bab9167024e6debfd66788e231880c760f2227cb482d0491cf10f7072367a577c3a205d3e73fbf7fa84dde50404bb53ade523e530d4c804774594fdb14a5186fdf8637a4e1730c85a341;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1b7a096aefe941b036d374b06dba788d047ccdadf7e8b68795c39d5dce52d2046ab37487fadd967077c2053f49687a14a6d5c1bafd5ab9c9c762eb1a3274aa4dc2a4767a3b534cd24ab40d90fdf0fe5fe2102471;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd4e1ef783ef6639a9275d8b807686298bc145099f928bb94890274d6a2db58180b8675887412af775c24ad47420a4dceb018dd3e1f8dd350e6905543521286f5b1228818018bb2742e564a1a025fad74bca40c4a9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf08cac47327b8022adb293bba58348bee33ef04b23ec19f32a1d8646de4acd7466b0249802ffc87b98568363b3759a63025131dcd7396bef6891128421a30a06938957cf52aa17977052b5137fd5d4eaca9588cb3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a03860d05d3b9e139a47d74135e404264ecace7239c39ac841cd685f4b0de06284c192b06258b999722c107333f535af5e826247b2e87956a94fe9d03ec1e920393ae4bbd015ac40829264ec17c389b775143a73;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7da01ab702649efcd821576b37d588e3cfe4463176709973564b864e767fc12768c9f47213b4a27caec50e6d641bf41e0bc3b52e272bdcb5133a7ba67acda1eeaf3a3e8534a643d054f43d276d0f736fe9ea53f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h640b3ebfbeb5a77cbd6a5cd4ee37c67b3c36e3e64a517c865b27fe8cbc08921768be80e2e13a95b1aa38f0b7900a385c79d68ef9cc63ace94eb4b5a9da772add9dd3ad8b813b9af904840839985e60f1aa355abb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6146b7f9f3c4c013d5710a91edc850fb8ee29fae4eb6b70530c02b5dd9d22ac14bdf4ea19f156ed01b23c3d05cc019b2d946f9a696eef26dbef92f86cc22345ae33df9fe7b27a4dc155ed75be363fccd637792d37;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb65bfa6c8834095f0b517c93efa3bd61851f6bac6b844b8c1c1888f96d43bd26a9f4e304f8d3ce1871aa377d118b2b4b6591ab5f5bb4efe2adc4b219615d8eb2cbcc48ccdc535b143cb37cbdab8215b1b79efa4ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a0383d27605312ba9b30e841545d00f4f8cef87580c9b2f550aee61ecaef4068248609df12f1e27f9db4c91b26927dfedc0841ee573d8813b95084a02f927113047df8684862f178633323bd1d1de83fbc86fe63;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7f9b438ea6663834b77185c11817c0616ebeb1c47817b654d4cdbfcaea29be075f16de96e13bc74bbea502ab51b8bcb5f56c51df85c738d518adc80f07df8742c9c0d059da6b76926c08515f4b7a6279898d13399;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2924f19a2b8005d92605ab87ff056f4a873b121b923b2e44c6577a22a822d6a8e05c38a5f5f0dbdf2d1c3982f9d82106a7aa41f8de8afc2eec896f728505a97812ec698387da7149bce1c618dca36e8fa2b8ee003;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha27a7b57dceb54d32feabc42ce5da6ee864aea9e92bdd16edf521cb0345912e584171670ab9b92c5f04fd2c01002783c842bccb60e34e621e73ff2ebb4c038120ecfb99a77ce411c3fed04e56a2b6d3bb1e89f4aa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb9ddc02f7651165d36cb91fac72785976a0a63505b306bc5287e56ce07a679feea00ea330d73c1035375e1333a672ba57fa886b566f356c81bdbbfc9c4595e8c9298642f59260e8055b39472eb430d52058cbcb86;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35f596383d428ccc38baca22c397fc6f66f3873d1b3c917c1051e455c0318b9233b745d033f2d6d8adfc08b6403e4cb8863919ed8d8070702a216e8c50244c5b2c37e1279cbab4e32ff386392ad3a3836ecfedd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5f77197501accf962349ff23327973eaf209573af7b15343bead42a9eee04f62b881c60796ae03b5a6caa4e46eb76621fe1090e36592e2d63362686e29df4638432f8951e88ce3db504e721d6c5a3b311660e910;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h38ee9e9102e8bbcc7e8e54730966202ae9bf6f26ecf3c003bae0f71b0f52b101a26d15bf8c3bd94d17c59fd662313f6f980e8b61abd0499d8d78c7ace8af8554bf04611138c688f473a9c84ff0512f0aca12fc8f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c944d4096ca90344ee59221b314871904c2e995a934611313c836267f36a53168baf9236e55c6de7984f3fca3183b8c4976c51a6d85c32d3e18096c07195eae18dcb364796fad280221008a2163e4095c5bfb7d1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50cf0d91ddca939d9a4af5eb83a3c605c0d1d116bbe5f1c9a6632194bd2c60dc87205b703f1385201f9e95187b4634d60f807e8e3e44718352735d32010dcd9256cde5dfd66c41904b686a095ecada91de26b2d17;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hed3322c46ffb68d54836affe3af1a4f185d31e7bb94a8133a858ef2fd0219ef4fed5882eb966a646c4efe029552ee4edf074bbf64772690867c5f9013c6e169716f61346663325cb4cec081d9a70c18e82810aa4c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h754e6cb12c9c36f2d81c6cef52264d17162045d468febf3d1eb4b5cb845c3201ebe91a81988fed1b7de8c649a0db6842831f0165fd5dfbddbe92912c68ffa9369be340fceb15c5cb47ba8621ca3a4790fb2fd323b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3da0ae1d34d230b4d2449911ecd113e3af1a1deea1dd638d828d8d93174f153f35ea4f00900a2a2d63308c5e6c417bbd034dd1bb9e174768a7f549a69fc578dc2b3388893b9c8ab82a38e17d33404e862870966;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc7d374afdd6f08f46640a8bd4dc636a9ae186e8f1175244cb69851716b0acde35e459bb11e8804310f0766cb928936184063d8e924094c8bfee056893c2a7ed5c1f1c69fa9531338a72305ca1da7e3819fde66442;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7baac5c4272bdb6894d097f1b30a764c325c723b0b2b1a8e90c903d5e24377698322d124c68d6af5caae9903907ad9897b82d2eac9e1a142c3c8ee7faa0f7cce61256c552b9a842cca7e6775fc8e1f33eb737de64;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha497cf39e790f2878247877dec3f5357267a644ff0bd059f689792242afac046b8ca4ebc3cafffedc004dc512fce68cba5390f29e3a61e6cd593b0dab84374b2a533f8cdceae2f0609b4109af649708462808f4c5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'head66043696a8a7308cfff32971387f6fcfa6c04c715fd874086a0914bb81f76c6383e12a2692618c2ac1823409a537542cc3049b68f09850cea0947fb92356a1d403ec96b20471429fa13bc9d154ec25570be5fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h384aebf71af87543dc7b0514524e7cdb0f2d75b6b2dc0f0cac9f7d3a3d006d61913f01fb23ecd805eb64bff0fca1d247374ec5a229f15097a5d4f017a6b8b0be0efb9e29c91874f702b436a193aa06ec88f0d23bf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h819895d1301b0cf956a3acde26eab94ef77c54eb8cc252b08f56fb9cb89e5f3a9ea336915771081949c0a2a2431147a3e51f69d7dcf11fa3762f3c23305c0093d68ce5c3890a1f7652cc0e68e275f4e8df7a92628;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91f4fe20a0d1a34c2a9e41f0ee8c4111deed71e8dd5a4df3a6aace2bb9d1cf821c4be8f4a14dbd3bc9eb39c67423240b123a5fcc71439ac89b57c29c84a64695ef428602bcb138635586cced9309735bacc495fa5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce5073c9f241a2bdd97a3ab17f5c93c4adbf01ba85865231a2f6f2db0d4a9472e0f26ca23b1158a9e18e886d77a039462ca89ca8f9eaea72dcbe962c21e48245ed8ab0f4930474f834fd428fccf251f52cf2edf0f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h23d1a33c92db3eae1686ecde55ca52da946852d31a8cc610d5275e3d2378521b788b06cb6e5593950f1593e8ff6d04d1858b406ae88ded229dc84f93a5dbe9681b896aa13c030f5a0efc1746b62b09df55e1a7d63;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he0b616a8d40350bd0ea2f9c4f04c4f8e0262f5d050b305897e23502950e02bf4361cade24718f83a747a53424888c7372dc2243cfa628742e5f28387caa8dc8e6c247e46f8cb0f0526269759e7def1b118e92926f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99b768aa2f2be0fb7efa4f7ad2dc46ecf1aca03c448df702d8d5826e90bf5c3da8378d5d90a4312df30b015593c801295ca884fd0a7ccd391a2db29f02c795d2d0b6fe639d195128262d6b541100cc7d45ce15cae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcc9252e6b8d7cf48c25ecb0c16444aa393a3bf3354399654dc523b12e7384e0e9d6a7a68759cc274bc72941aaa2f2aa36d9b182e4fb8a9086642538ca2825d6006b778d99447ef6f0f3bde026a50bfba361a1f13;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d24153bd065a79e84d603f9dd07408ac24b668b9c09230fe7f78aa5d432998b64871c8423d8e7746b3fc75f3eb5c6c64b5015869f9a6787519101ca61a8441140bc43ebd40168c26a478b8dcee4ff187c20ec6d0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47d16793fa1636f2c09eabd657d3d0f372bfe67b67dbc17da0b4dba4a2546ec2f29e7a177bc76e3d6c106862bb367142b0909aae3e8f4adf20b9538c821c7ca94e761990cbce211e05d49a7fd4610a9bdef72b885;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b1a67cb02ce5a5605090b1f39cc324bb4d33be30be959de8edda83a51eda24a4a8e5cd246817846d2e4ea1953b479d55b3eb5a2939b8f09f3493b03c170d96f03842763c664e77ebdd94f295d71b6fbae8e5b834;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h978e21b825b7a40e5cac2a3c85d107e433f047be5c18a8a5ee860f17b88053ec83c3839c6040ab405cdf10437eab20d3ec8d3881834760ed1834c44f1b3b90db68e4d908cc7aa8c1964d950dd7fa722e3ad1aa180;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3d7f9a58c5a5ce1be0e1351f9f329b3e7f1c367b1d37bdbb3c08ee83a37aa949334c207d4935ce1730eafecbbe3cffd31cd58a35fa6f137dbeba0804089b6fe7e62cdd049f67d29986e7fabb7eefc6ab9fdddf57c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc282f9db8fc8c3d0653577053a93f57fe3f723368bfb31dedecc10577247719becdfb7043b3143f2c0d2cbb2f310aa46296668c4e79fbab94a828e97300ffa91c017a6e04ad66b601ec9b34f7f39b873f55360c3b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h75231d05a010f0b3113a374a2cd1474401dd4a4b608795ea96cdd769c05d78838b35620a2a78ba3c1f769e0875d10ba6196dc2c31774b52b99720ef82ec8323e726fbe2f56f4b55f4c38f7bec77c6c5b3c7f5a262;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bd84c96c02323c2ecec6747e8de0213e35c87791586c6a798cb09c09d87d7361f85ac1ca44ad9ceaec42f41dc913ddf218f8d6f02f57d320bf75dca29379dcafd668e70c872af499be0105ef69a8cb3b6337f01c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d5324e97e7a4a63dd8d58b4cc147a353773cad50827d3ac7029ec27d8f398efb4776f6b1c91c005fffee2b9c8601337894652b8a177791956e9bc195feb16b58b80527873df50fa3d91c8a858f36447af1fbe2d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfaae1cbe9d23144a915957108c190c1c99a1cc5a20fed641afed8f4966629ca515e401d69b8208f19877a6ad7f24340f645ebde36fb9e762c21b2d0ed6b75d529a26d5d6f635d4ab60ddf5537c22afcefdf591f06;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacc9cfc3d28157caba0208d79dbcac7d44c4d1f840b34f64f38dd2ea49f4ca126e92b6ac8b6ce830e473a58b8af0185c5823016c26d6d4221ef6951c1485e57f043d05088f22276f8a8feefc2d578c7bc8b4113de;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb097e780801ac1a3137e088734db0e090c282ea81f7107ed893d1616bdb72ee36e18086c19672cad8ffe15e49f23ff03e949b7005a9ad8492f778a42ab9e132c333a4e4c6ed3e8cfc9282d88d61b0a5b62d517c66;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hab996ffd8a112f21d52ff7c76bcb0265377d34c4cae9de9369ba44bca33fab89c362a6d54295662dd0ab96a111cb2121a9f21bec1fa6560e3fc7e30d92a075b7f3dc189fc49525b13a2600484965cca300f09ca58;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0b48b25914a4f894344ebb5c829beb268c98034fbe9e76dcbf32567b3ac6bc22694dcafe3cd0f0f277222aaa57307edc49e902a2b32d7f12168164b79ddf88fa0bc426c2ab01effb72e26138ebf5a9aff65ca5c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1dd8605216b849823df32b292ae6d51e4e68c7be00305d243a962e402badd40607c776c3de0e1ce99926685a962d119068577f4723092c363af86b9be66177b5c1415a2d1d0d7f68f342ba59a4ed91bd5a2325849;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9cf5ec3a6e8d458a67a3aec2837585861ebcc0ea033cd1426fa5fb1a50444566b2e9840385f1ee618ae51f9163b190ac505707145ed742392aa7011f56f8ea990b7ffdbd6127aa6afede11a1a02f28ffc21422fb1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9af1f785c641785327f1ebcab4ab60d274c71c7b8747da8b39ccbd988e9caad367f18a022b2d76c57d7e44ca4708681d0cba79bfb7f12d7526c665600c5b16e0dd61cf4d270172589f34b89d0520852cc1d38496c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee590262087d1d27e82dcaac9f3e7caf3126459530d11e601581bff4c4961803f339b26385b5cd3190ea44e47b64180912f1063b59452093766575b7834a775b8b272be970eb6dac3216267933d876702599fa50b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha7fa6ae23c8b6e5a105c48678b528f08f03f0531c61a942a5d5f1b3b76865c509b9ab1b6d82c336df79b1bfbe5efc70a9b8ca086e536c701aba0cdc6ea3a973a95cdbb278aa2f50bebfa033a5e53532001f9c01e7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5645ea9e43918e177d3d99cd9b11a51e2f80b4d6a7e364e7cce71da54a1ff299d6dfa0e504923be761de8640ac7efb36fcd2dbdf4257adec089faa78ca876799da1a7e68aed9b7727044d6ace7330b85482a4323;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc0c747e48dd11f451f623bf6220445366f54a705f302f5895f86a966c8a2596d2de0a749f00b5bf5c4d78ea5202e068e6607dcfe3876eb14e24a2a8de01387e40d63dedcb6ad84972b7356e0b1404efa786859dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0d4c42d0466c61a36b4aa2046aeea4307bb015f48e2f810bed85604ea464c5a7ca48bf3c38aa416b9eff4b6a2d1e926fa2d0f7ad87f55b73402433fca46fb48fc81b61f0de8a6872110a9a6a52e45a2fa4a4662a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfc08303dad0233a77b06cae46db9c938b758ea10349bda267392aa649595e18e97894aa40ed815ecd208561cb25f2ea7c5369f5ed52caca0ec38594c3d7acc37f837bfbb18a0aff0235d49fc6f819cc3fe0ba7bf9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h491248006f5fbbd6da290b3d89f329f174a446f9c1822b2299c6b1091978a3a172b77a575aa151e6799ac992e97868a45d9da6a4b7f5693e3dc0f6439651a67c7a09682574b90ddb2e53c9046037ab6598a34a8c8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8da505159c0aae00c684a0f4dbc22efafb3a543832489dc9cdc15bdb641497723c32603275e79ac1f449aa287057775826a1815e160d25b79c9a7d589dd2b9f2581c103f6363ce1cbb2f7c1b6f723341813d30092;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd6b2baae2fc13dcc830b63cd5dde574c64ecc56ad57bc3712b8dca2a6bb95a7f0932764585c2a7c8c551fbcd603eddea389fd673e2d159330d8ba57391710371cf37a40198e463e8dca78a09cdad247abdc501db;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb491fc3885e51f6c6c4147081261af9774d983c4fb3f2629c72032bdb9e42d0fe155d9dab2549f51526580fdb094dc8674477d3e98603a7acffddf9bac67fda41421fee5dee934f36f9e1613df08615e360b887b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd71dc3e90ab98d9f0ea16f6a4909b637b92caca6a764c2a862dc889eac7a89765f76e9904e5a5b13b4738dfbafe8f986e38c2effaa57a2f6909b54693d94a810fb2319ec253e6c120b79bb997531c127389c794d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5f50018e56795d54091effc92cda3c782477b00c3baa17ea9246683302bf26c9761c766617b341f1f3508ded357a0e7a3de7644abe8bdf5b2c44983147b08ff1a470385195644b4643f3c348381c3119cd34aa47;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he86e1281181882fd512915bd8450308e37e6bc8d00640bea6258907dd08b32609ffcb84632d3fde8007a1858fbd2ce8f096238631edb0a3ed2021766148521de0244fa6c718891f0403f112c5e6ef97f6ca89e4cc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9a15e5f74d3cdeffaa93705ba95b98d23c56d259cd9fa3264b3459fcbcc759e482a1610728e46b31feed01b768c1f89904253cd4287ec4e6b6a74aba78a534619a8da571241437507575ae96f3fddedf4b527005;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d77085bec408e5e45625805669688fb4b8bb8842be11ffa809b588721e86cccff903742cc1f6ce7498d3839bbcecf53e45a48a89f3ab92f673050906bb2cec2ae0daa28293a80f7bf41dabc864135afc3fa9dce2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8f37436db89a46980da2968fa5bf068118c62e7cbe722da8ad05105bc6e8439b2c3f056335ca88b0b04f2e6ae500d5ba29ab73d6b56fd1c7616745f9ca4fa88145fc299a7b1074545e22dca372e14518349e03c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fe60fdc3c11d2aec68441b2a12128baca91af984c38a3933c7617103f5a7cfa0f13de0988f3b60cd9f5b6a42cda8a3dcb50a9396acd761d88fbb03333bdbdd1ad3ff3799a703312c005d476b34c799b2e6180b01;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcabae2d3a75ccf52f09ffd15003b8713bed147cad59dd3c6465d49f83e856149e315504c2ec92f5fe6a95fcbee0a7d9ec38a4f59d735d779568a21b02aec14a1dabb0861a0b74daabc99a285462929de58cdd0580;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c4436c45f7c42d4fb5ddaa3c544765bb79c7cae195b0b5a6585453fda0587aee80aaacf36935a0fa6a24a780372fa2be11b10764fddea7154b3ebb9a9194c2a2008a873d20d9a422b8b56029a0a709617b16ff9d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h62adb5395eeeb9822aa178eca7ee0c213ba3fd82fcf70a2bad2a34ed8f3ee4075aab2b0075ad67a43f0202c85ae05a9f9cd58bc24b9dd80774d14e68eb5894314c8a81ed559c1ca63cad3db34eeeaae8a2205c5c8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d9a062a48892c9b515ccde75a225d17acd6b1405bf6e81ab193e7b2835ae188216586ecae62f00a90bb88411e222cb1276cae063cc1dbc4981e71516e1a77f1abbfc23e18838d78718196636e6d6c037b19636d4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h229d883945b6c0ffe787d730f73c16d154d1c703dcf2349d3530164338a2377ad6630d45601d2696ee9d739b584d16cc15e738726d770b32855409cc3d11e226e9e6f51ffd657556580b2b33e39a88893a16b7cd2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfae0496f81a0c8de0d07af308fcafb5dd19edebcbea45aa232ae192db8878096970c74680158cd5a6aa33cf5616e8ec4bf01dc8acf2f8c506474117cc695013af0a5d4c6a3c1d345098a262e7ff3d939c74aef11e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba55370cf974abfe115c0aa2e84ad176631475299d9641b21f1f59e1374d0ac6f1650431fb3a1746ebf0f412f05eb55e05ede9b7397208c2c34094078178ed343de6bd943aa3c3f69ba39be0486c1624a89b74c7e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb70e9b1cf282c345ce94bcf9b854da733dee44df12c8740319dba750634bdc92fe2a2ff85411be45f4af9893aa5a47df8e69848a4c01707e44f7782aaa744000adcf5bc82f60b1704846e875fc675799cc2eecc39;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbfe7bfff8ab3d13f585f983373b7bf1365b8de03b759825f8cc4c38062b0b1dd5aac59b63d96b35c388007b8eafd809b2371710a37db8b96e1979f5fc06eb53a0aff82c85ff1b65cc75bd05b0e5af2e13a212039c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68ae4c24a78351f89ee487266524718e64a53319b3a938fd8089b859eae0f82e674e188fddfb8c18345445fe5448b80884c1850c38c1b8d7ad38babed7b0a645d08ce081d24e5b24a4d8aefc27115561d97eefbcb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68abdfd39039b75c5a71912db6f432ccc547ac53016d1991ecda951a2c8d56f7f76f961d9374602536d35bc3b53c60339f07e35a01e0c8a47882816547261f722effaa387e9ded36ac2f1498880a96b58e5444dea;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hace5c21f02451655f3d5ee305394068a29a12cde9b8ca76d04795e643fe08c0984eeff3e849edfb94941aa32cbd1d6b6d33525d1959c99e1640263ed48bac0f0cd39c161c636c6c769fa4c13ae02ccd4458bc81f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ecff594287260ea44d1e14b8dd3a40f117c6d1d7a98f78ea65ceea887ec178ff8390e6628b401298e12262c76578772a883e8debd11529322173b335fe2caa83254ac412e1a426f0935de14ae4b24a41cb0e51ee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h399c1f320c7a9bdb8712eda338c4a05ea136a1ab6daea9666bfb81608f1f9be90d085d4737820908540ad2be5d9959d74f0b865b6801be3f4e8712e27e5cc07d4f0a96aaed163e790e62563bf71878712b182ba31;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf88969d97b2d5010e0d981728ec74ce2917e7ccee1c48209802059c9973994a360dea84114c0670baa7e07aedfd520c1c1dc64e4e35e70b7cbade4243619ffeb1a1b47f4e9ff2efcaab3ed6574741f54aea7f4d87;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4715bf61e7d46cc5aadfe3680bf81ea6d1c6eba8aa432facdd21684f8c1502acfc1d2938429d3356ed69b5556400de86f174c02cc478dd64c54e0f2f576610def697fc3ce1260f18e7f96b4e834e02db6cef962b7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4416e7a44ae1cbf1bdb28b62d11fd4ce971691eb216894ca593aed6e7aeabe01d12f3d1d5b3325d0705e589ea12735e70c53077c6bd73f669a1b4d9fd456570c370428dd91fa3e2c1b394b213f9a338b7ed452b08;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76b7a52be2b817a6ebf337ff3af94192d42b366816d7a59ff02d714472ca3353652c855e73c058773867aedd640590ba948c95a9099a226dd6ef4f29e07a57814029886ebdbbbffc96f1dfc8636aa88449937cb74;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0fd03e2df8ccbebc363218640c9b95345558924820a4b382b94ef8798d833c40768c1387bbb33d4be6142cf1326c09fa652ff8c7112e85bd7e93a732534c0657ea9277efe0e41b869c3d98853ab980bc1e7ec9ae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc50522bf31535cc8be84bb5662ae2335cb88a96cb15e02e0e8ca108986ee98b3bbfead80e6a241c7d1352fd6f35545a55fb402b2e5f0c4c1b960afe519c0d94c81b10e8a2a4964046569b0ede7fb126e37c6f7efb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1f869fcd99b38ad2376836e77494e3cfd36ea43d4ce8ea058b3cf5f6f5cc08a3c4a0723182f6a19980f4362bf60e22573c03d67eec4c59c3034e5f43dc2c86bb8b01e8df3697abb8f3273ddc4623baec1379dd322;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafdc53aedb8377b7c8cd3a700d336970490a5c60866e945f0afd606a5001f178d831b686a27344874b658d44a39dd0cb7501018be01404187e6e26ce7a28b1f33949bcca49f67d84e93e5fd20ce770e792de35bc3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h27b2e3a5e40ab2d2722da9315651fa374ff12b881fbcbfa6388193c4b2fc0a619be609af50ea0809fce0d0bfaa571969c92b0c041a36a33dd40257049b2f464957eaed780bfb8271b26ef7631b66b8466c2cdcbd2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc36fb967dbd6300ec650f06686b036197e3f39c9850590a122e00948cae719dc6ad61f1e64a681cf6967c70109f3841294f7bd4cddbe9f7a3e8d8c86f2421852b351dd86769723d5e51facc27cff531a28de448;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7af16327a14706091ad40a4c67fb1544ae3c780addcbfbbe8f5377eca084a2a0e0474fd8f08917ad3aabbb7e60a8f1582df6d5d65416287d5b711e44101cbf1e2183d420a0dafdfe720ff5445da4bb0f8dd96e87a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3527a66d09bc68e77885b8624b872fa87aafa04c1b3b93823dc30b48f7d869ef67740ef571d65335fc2aa4ab75592dd6bf3477c37ae4b60ca3375d8e7cf709f8926d096ba185999747623a86a97c7f03956f2ed54;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h897a61a384df726e55ba8ba0716284713dc375844085222788736e4d48143807ebc184c4b90a13c2582c29480544162c0c7ec87d9c6fdf052693c158dcd37baaf98371d8a50b1ce271056d1c320205cf3f29ec9e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7d0bb503bd939b9770c6def023b3a55e12638936373d3484dd85a5d0408446ce53a93835e9df7269b050de17c583a9eaf1fa71c5086764d30cb088e6f23d76359c6b7a175385f7aaf455d9ec1c0c995c80eac1a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c53553703b79c939826e2571994ef7d13d3184804adee41fca00074f024617274e5ef1a54738c3d3c3a985fdbae6288fa2a7780efca2caf2e67fe2e090b9f255baf42beba76033cedefc4855b383da1465d222c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e3435891cc80a2f8ba10e159f90ecdd08669d228cb98b3b58c35f05ae4f231a4c8e7d5d521928678647ab2e55fb1ad333dddeb0c9c4442007e3b198f918b0e846074a78da2cdbc8298218f7db04cc04d39e3f1fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf537c13231230088e39a25389428236be5731da17b83e6e10a27ceb442ad5992e99b7b1a692ac2bec3ef322a6ee83279c1bb840a214fbeebf996ddfab0302a30de815d46faa2a771a24148ebf82bc3304500971bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha9cb80b413dc01f9dc1ab344553726c3fd96bad3bccc3fd24cded4448c78484faf37d1284c3d6ce9a3dde876666d61280830b3720f81ee8c9b136b806afdd0c4ce6cc34954896b7c1e23202a7c9254819d7cb0e18;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8b5effab1cc9f68baec85b9ac27644243b44383eda83560e457c8421ae7deddcd1e169d7b501db2a5a57830397cb82df831ce293dc287e28510722fe642129c1644ecf70b01be3ed807483896ccf2941181d1def;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22485100812c87d87412455a77dd79b5241c848e77a630abb10136fd42f3f491d6c4f655eac89d100cbbb5cf64a6ca0cbc41f4166b5d756320cbb0d194049ea45727393032a7dffc170260a12adbbfd53345de838;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haaad1a246879a7bd5085f8cfbaed70eb052d45fa40b071548ca99a42902c0f2f2d26bf5ef7d8ea7f31a68aa1ddf8cd069c6403781a90d24ed60e37e4012c963a5dadef16060d93d45cde46a8d42cffba6fafdef9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9b9a23890f8c3a8aae00398e5fa6f5449ec05b7640260421757700b540e9328ebc26d13073774fee85e8b23a2db0cbc3112ee47f56d4b01320f29cabf4adf5c2187ea2520635c758b90513a6bea8daaf3555deb9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h329e90ba80106b436746da7e9a93c2c952bfb3bfd09e81db3034840569245e3bc63cff473d18199fc08cbc52aa0ec4dc0ccf2f36394b4086e0c50baf2e812dd26e591f2d759a4801b7536efcb6394f413427c461;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73aa16a214e77816b0112b76ced20c6f352cd4d7c54ca2e9a0b6939149621101361dbe6a2ecd40d904a515b43ef24a34ef0975ddd75480d44c3156ce3c6bcc91b61c722caa9fac7e57517eb8f3e5a2859cda1ac1b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48d7a1074748f99a3dc644e6056e9179e372ac7ef1c84d504a8178c6971fd135e6dc2b28977434f438efa0c95e23b83e0474566b99586d8406ca5a956adeaaad11455920fabcc91136506449624b4b537ecbc8f34;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50def24c423485b21dc132afd7a3a9580579a908ef364451e29675e53c5a3962bbab55067b9758417f57b6cba885b68c90bc36d11f0397edf00d26a24775c4730c54d2d27b7dca848c09d58732676fdd7458ee999;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h86de3112285b3028afc256269afe057159c93f32b5a5e2041a12abf7c2d6a58aba00f19b22ad75bbb949786a5524ebcbcc247f8d86e834366666badc01f37e977163e1857473b248933bb479f9659cf431ccef9b6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16138a07b528a8a53b3b327ccba1a19f948b065afe04a41125ce9c866c11880b1179503219ea185affec35edac16f6bab7c9401524e4a4935492b9164f628ca3a09e7a141e778d01521e070d06920b746ea55c604;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hefe1a38aa26f7a18f9de4b053581106125b3f628dbe9c244261938b97bd1f46043ccc7e5a35ee2d4f8acf9b0465b6d4d23b2b53ea8a9f5c900ba35ece6d9807f04e328d18b8ec96b873b55ee856f2ceca0a327912;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hef4cad2b4808eeb7fcb3a7dcc6bda04c933bb119826e71c95b61c6b7a3e41b0f706643bad685a01cefde39ddd1291a2fe4c34d61e31c7b01c0bb8c65464a3992c9a0d453a740ea6649ced05df679b66489dc12508;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf8a12dd838caec6c41e78dbb710cc87da43020c48dd0e6a8441dee72682f51f1c835c7a96dca211a04567de2e9c5cb5579148910d02f7075853b23983d4c040b9a61d150d96e2d254d0329149744c17157e4352ad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fbb1693984207289d3a104261803c7a18b4945f46ea7f29c097ceffcbcf40618f6b5f8b3ea04c97430b577f0f61bd21ebfaacecf34733d2bd18cd138e6c7adad585b55a57efabfb10b699aca8c3c93c0521a809;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h750964bdc5284b6adb5cb9bb87201add2a32ed1bdc3962608812c37e6f8c85e28062a8c41d0048b84a8af6907738bd2ea9c3165b667a352b8de92e900d4e2a17131edbdf7659d3810f0b3a1fac3f1bbfcbb4381a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9549751830823a8cc7d69959991a7010bf6f6ae4116b5c94b8acbc1983cb3ff0a02abf8991ad77b21358d93178dbba1c7279ee62d00a405cce72b2dc97d2afd34594c945d75268982a171a9c70a44614a36cffc98;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb48307668fe60dcdcd9ea70895a492f8a560e1f98344662365377996c2c9279c11f31453fcde212b5c3ba86a6389bf5e6537950fdb7bdfe068ceaf4ed8637e466b57a9831452e8f02f355483d2b999ff7c6214e0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2bb987d9a21fc3ad05716acf56a0b8d1d56fc8aa39e7e49bb1f67024889931e3bec19def32891197a84ca5dd130bc6c8878a58e4d5b5e1fa6c42e3b4d209cf37856f1f18ac27789bdc3f17558ece5f55e1f678f3c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f2b4089b74ea27bf05a12591a3be4b8d28654106d4cf6927a2dca88832f08cb0d5b573a4949da2c2300d9fd3d2d6fa0da38b82499cc9c6ff88b9569719125ec53651809a37cf5e573ac275dd14dc1d6250aff025;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69a1858928e59dc27e43cb3ef1739387cfdb6f44bc44d1b90ee5a7ee4b3a568fe7f16ee8661f487015db84ca359b02b6b3ded51973ca0ad5ca0db0efa8d279b502755338b0f13fee87c2774d93f2a70dc58b9570f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f4a17e3efa816c456c0f2ef21cb72f96ba10810b68b6ad737a866767b946b3e334824381970daa9d0832314191e6a4147b071b9e7f5911eb140fbd283d8b605415f4df973f472726c54d6bcac0426fda3038d864;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h157cb36c7550d09f9d5fedd9c7d6b33e4a6134f843a862cb2a90a3331151f737f5a36df440ab102cc28e99f90f4d4d9c93aeb3e2862e286d16f02f50cff0fb997c70ca73a7a6ba6e89640ffbb75747b9085baaae7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba4c3c2ffdb221b14a1efdd28b0011fd19d2dcb854774aed68f1b254c8b2c47fa4b5b46441c855dd2b88795f7b1ce9f7c0088cac6fa56a8e7d60e25e40eedb22c35b6831f3b6358ab1dc41620db886fe5cca0fcf8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h50a137dd869bb24a2b1992572f24dfe8b4419e901121577568176767ed0e454ac85d6583da91c6cd44cd5fc2bfb6171bc925e4df9f5bd0c2f20f106b989fee5b77fd8aca6e2b546d2583263e32f5315726e44740c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77b642be267f0c8d6043173c9a86df8f1b464aa2c7172112c8b82988ece9b1644fe22067f3abdfe586d84c30341ae66801d55284e7ddb212e47cc5cce08aebfb64439af9c3ffd5f5a9b3f3e0038c04d065db09991;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c71c19562f6e71d3a500d416109bd008b5502703839b496343402123a7932b5384170a5ffceda804713fef15c2dae5183928f22faf6546ac6e89f1e770675385c7a45bffb1abc2862418f657c4d1244f350b49cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h376cb351cc36789084c70ae8d828e57f170167d231dd88e29c10d394982739ec77b294da63baf34f84da18c6ae3a77af9848e9aac3ae68ced68a8e437b2ca354bd13318586109604b027c823cfdbe52bef77ba9ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h630a8fa35b80f5fe091e0a5c82c049da438158c89b1acd2cc344dfb6786ba585685d47dfbcf29ef3c9b88bfed68e4143dc2de1f9d48ad367e2c19fca4a5cc50b15d05d739dfaa779fee7879a95f7351b48ebaf171;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hadcc5f2f958f5a21d202970b60e5b67da068acee24a403816e1181526cafe9355473c612e1f44f4161214b456ba1e7466c0a0ee196d570b815abded63220171fb301a6c14b7a17600a74de275f4fa5b79df5d41ab;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa12310ae0d4cfb07582f29076fa37c09ccafb1d7976efb2e259335674dc11ad80855c1d75727965315062eeb4a4fe36c9c7d6dd7faec8db2ae6fc084ad3db61393cb3fe53a6021740d15ea1490446ff077c727bd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h88d05929d76d4148cafc521f57d48deb4acf87fda896d83c9ab8cdab24eb7a1a8f25c0ccc2ae86acdee3bc1f85c8bad1098142e793c2c8e8a687bbe04a620a9355feb5eeb9bde0e77b710d6edd8af602543d48e21;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h16a750f04360aa07392336af20f4aa83e9455779f68ccb891da1770d69d4c0d59145dd0f53c51ac8ba457be3254654e925faf104d7823912e8fd0381c8186e0bab2692b2c45fecca3c44bfce687f3b3b2a5006ad0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a22cf0db273595e9ba36d420dfc091c608c6ad3fa2e205ebcef930777468563764528611bb7ea827a0a92695d0d43ac20c55214f545281c3627c4723799f27499bc02e235b6f83ae0bf1949380b470b02396239;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f3ea5d84ddfed07e984be6c65a413ce56c3879df253b3235463b2432039121f83921bf65f4415c90193cf266fdd2ec8b4a0cea8f95134a9bc9b628cbf8ad2c3fc97ef38ed24b739a452eca3a23c149322112f8cc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55db3f642d030ca27932bebf9fb23a7df139d1fd1f62659849a941d371809b9d251acf3a519dfb22911937022b66939efc00d1ed8bfcdd6ff40f76e69420c9eb896ba82f1ec9125e37ec5ee12579f9cc0611b54fd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h46ac0955ca11b6ab2fe29d9118a8d4640c944da3db490a61204fcbfe626583ccfc653e0d774e08b2641f93b27c371462bbe52ed6637700f4fe1a1d93207a16ce8ae0c4732f122cd9d1a8d241a1d67e04add7ccd55;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h15aac7c2dc6ba3c870593366dd27029c2b75c1181fc1257d248cc29c4dcf09d9a07c08e23b421305a0e4a3332c4394e26a60a4245737da66db69c4963476f5a727c9584f60e37667f9d23e07f45c683a13ffe2238;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he58ee57198818e136e6c1fbce846a2b324cb8d4d4ff4ff805ee1e03ca3ad817f695a55e2a9f41fa4dc0cc4f306c57d67ce4091327c8f95b45ce4792e575bee5db915a2088773e1d9c6891412ae80c958f844a906e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3cd493aad50c22d5e51f877435b37fcf18a28eeaebabd478ef05aaf863d555827be57fc52b53615a901c7e3ed52fcc6747b702497d78c68b010c5ac29d811e3a66051c130693069b830cdf7dc0e94a96b967a4bc3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h437598ca2132913b20ade0f206ab634a3d0268574411ef7d2c384488e6e8c3fb933c7d2768f33c2d0c017b286442c7c70b361121e76954a5f6ee85f56ac3df4d318859f49269a057af9df5758f9544409fbc20511;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4f0fb7f48595ed25a96c93a581420544d100c098e305d5165e9d070e0b3ea425c7c7144bb6edcf057057e0b3c11e4213c0cd4a8e06506408753cf831f77c4f55d4cfc800b2124c02ed2fbaae13513036a31388b1b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e1afa72ff6713f0603c4871c81f4f186deb7068584cf7cc81f9828a10401a75754d6577dac4a34616a5ba6e56dd7d84eee866eae8f6b5b7f7dee5520fe4e9b28f780f43c9ff84c1077e9ee683494f840894157ce;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4995fa484e366973a7245fca9d20448882d1b9417117c2cc0486b15c2bac9c690e021b3dcf84c9149bdcd9f7500599e3bb97abe6d6ada440613a051f51478584620905b9f74955966b00210f39b3cbdff35e0b8c8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8452ef809cf7b61cc5f6dd058a95effb26848731968e881a0060a12579dd4a264dae7c01878283b2d0b0ef4bf17c59c0a5cf00463b63cd834d1535848c8c6ca53cd77392d9da0813f6c5b7027f13ce2f02ede82eb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd393016faa4f78a5cec01fd9f1de602682e87cc5398867b46e9569fee6ff73b916dc71895861c228d3e360030d92d208a1f99f168e4be2f7e4458f57176950513e3a5f85c4016cbe16b9a05a57746c2ea85dc3ac4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc7c7125e8f09f9c7e078f7dfda31b57ed42b667b9fa592990efa0b965cf539260300af5c7fa547b09bc0df618263904bec08951b14b10e2ebc429dcdcd0ad850135c8c4a58f4b027317cb74c86c0aa37c28814e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1992f9d63774722e968dc2117295f8729ae4fefa0ca76310737ef635b67efaac4cc9f57812b487807510eeae948c29d97dc93e96b10a60e715df5e4878e351c7cbdef9f8abbc886d88beb0c141e8a2448c36d8598;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he6f5e25489442cc4865c2bb8a844e2918276ef6abd971f487d9a4903f966b109d3ee02bbf229e2ff0a89e8caca6ca8e71a3e2e22a4743ce8a12d4c1a9044df115c09c0cf8661eb18d28818d42224202c82169c8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h686f49ba44af8b8ff535af47d971a02c1cde5277333434861d1ed6848a841bcee2ca11b60437dc34c179e8c2daf1308a542ac614750071a3edfdd0d5200f0abeb7bcde606e46aef1c85c5bb0bb995a2ad7f03c65f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h32c221edbd7de473a31d7de9b4115162d3ea3152a2bb911b33018c588e54461df999be27a9353b4c3d0a8fc5743600352567c46b366868571041420b4546beb7d326a546db5476b321d7e5b0ad4e967f18a73fbe2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h54a99a51ac1383808f06bccf41871daf0a4202e5d800a52c3f0b2c0de547253203ed24245f9f3c085511c46d88d935ccf224416b8fa4e425ddc6af5e6e87e8a4222b8be9703be994e321ac71f5ba0a811485515c4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h18cbd2da5ccbe23d53823fe17a1bbe0f8207be2a9b89ce29e7c66ff8000f32ef2aa3b2d1fb278ba5ee01552e01f0e0d0c4e517c5d1988ee1f2d46f8f79bddf750239cd8d090e7a2c005d79b5cda4e38c2dcd34a34;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc12bb6dab6a8744a3c356fcf0bea4cc012ab1283ff75d75e5f15a189aa45fdefee36c6641c1a3b6a7e8d7f8fa9644bbc9f51497f552baec5c630e60b9c916af869932673165e313f4d9819c9f343578a3c2ac22f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1918fd2cc1d4d77973a61b8bc0c3d33a2e1433a8854aaa3a15bd9a2419664b669c32cd3e0544a8af2455579ecf92a48e5233f5a900fe182fe79d8a8be12806ff0886dceff1a2a6bfc28e95b67aed673f3983e97;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0c2fc9555439c827bcca572f61251b8b080d6adfbdb3e2d2eca22823b7cc4fa532a8f627fa95f1bf6cbe2c89fd499c66f68887acb21425ed28895454f042f04d6fb9139ed8f8166b5656f0d232415cf8a7e15d14;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f29e636bf115653e176cc9a4f9f7d259b2c20065f7f6ba522fdb996bfd945e5013b8faf2cd99ea48145e8584643798499878652221e3140cbd96a493e4e1f5d48f7c1425f626b3b94bae39d45013b4dd8ee5e434;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d23c6e8079aea2b090e01c358357ecc2ef7a07a0ab8d2892f5f8330110c527eb0341c39f9f5e57722f7163e259134cd7177d334118e0e7bf9a26ee628f57daa595f442783cb583d9053ea7c85786442c43aa4d6c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43767e50ba64b8ee6f7ad646e30a6e1ede3ee8d7481d24d9b57bd9b2002a12584021af9f9a66a422c1ab9264a387ae2a89de0b17b5cadd7b7bd998b05b62787e946f5e500ebe68d7293579a02b3f96f185fa256cc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2d68fa1a657d3d207f0c40ceb82f38ac1a29710856dda57bcdfb917da4aa06925dd604542c10bdae4287685006ba7abdcd913567cfdbd9149a02ad823fa847ed684893c6618d7e82cb022430baf039b9c072dbbc0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haeb1be38613376642883cddb3dab8897e23884e0179bc2434a42d0d7af8957651f1f1f22229ff96794620416805bf07bc4037b17d6370ffbf5221218f6c9ea7cdc1a8d5f5fa0b061a74793b97c2f7ba63ddc3040d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3fc486d0923b718170a86de24e37f3709085d835c360677fce74dca4f184752295a83ddfa0ebdcb7b4928b445df14ed05a4f051721958158906fe2bea03a71aac3748756c29085ea22e93db1a1360124a132b7a60;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7bc754b66a36871c5e0870be552bd38870362cd405820c6257df2670a1dc70711c1f079e4dcd34ba9ba52da865659d48279cea02095b07e6b802620c8b63740617e3034831433e6ee9a5cea20610eb0a20e17c8a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80ac10d073e6f64ee3f41f0147a3a42b19d32a29a478c8d9513a78792945221f18ff55b7a1217398196af93deb9b56e6a583920ccaeb767a6e48b77a7971604b14d6f5be6239327e8098aacaf6d25b510776d101;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3a8fcb223292ee60841b9dd1315deb3569bfab48e7a1f16fdf7219a45bc6aebaf9f49ccaabde2ea88d636de3f09401b1f606ebee89602efcf41b298535c7ec556b1950b451f7b2e3751897c1da13a9cc6cf5c4448;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h499e1abaa5f5bd0b1f96849de17f49eb06c7ecaae736a7d28d8e847cd8d53046843e3f6d7e8e322fb32116f713d2c1f8180a50ec6eee56871c46028c7ad923b627c2b82aea8ac53993935891fda277d147fe23c7c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heeb72440f42514bd24df07ab1c85732bfd73ebe85a64ad90531d039e9c04f09fe5a5e7949b58edba4b66c66490ce05d9e4623dce0f54c2a4a1419ba82bc6a00e0642f03e99f019dd73317e9f2beef77dad973608f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h307118d72c7fb1daad3e911e5ff5bc0a75dd4a4f01340c941b685441639d878bb10ee0dc4f78274e53c6bc00b143c1b929afb5cc0bcede0ae33ba46afcbc047b55feec55d06d653d5457b098469ad03440a3e4385;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b0e78f68fec0459167aadd1f715e3b99b1c18a3d9d3b36b6df08e8dccdba231cede100c8f11c98e2f889ddc52ea90ba4c3594c2d1178720ddf25e11492bd289d2676e4080eac0fd94df5879f40f63cb70dc581e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haeeeff41690c743de6f222c02536880f2abebe645dd8ecb34fdeb7203240111fceea8eac83cefdce9d958c650a2b56f182ce73d6816b10529eed820311d012e903b7653a631f4aab6bf8feb1ef6a4aed38137046f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h105994b22321512ca16cf192fb377a8a30124d3d893bfe63d69cc6fdd07a58280f371cc2077792a01195b5a23108f69d672f38b3e1bdb38de95f52225775d87584ed6f4efd3b4a440916ffad49a6bc465c1adc38c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96242aad84706243d00fa17694013de585f4c55b006fade15be99a510df744a16b8a8370b3a16a112d3ae6c0d5399616f29deb8e1dec1a88b57fbf1c352f65acf930db45dbd715c2d12f7a0e6d8ea719057c20b21;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3ba18a3275e022cafd1547a7144edf696d01885852ef8f43022426fdcf57ae64b5428b3d881f0cdd6fa1076f43dca341bed3d0be05bf93198c701cdc5b0f8d6ff1934a70c2910455a8cd0f86316fd04c818277d05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h595f2b36600c320b0ff82245e8dd5738c28e3f0149a199ba7a64700216a7040880a360428761d0dc4998eb0a429fba36d346376a8e7797070e7bf87e402979bc8709fcc89abf702bc814860ff4b18a9c207c9bf62;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h44e1fee168669609f1666321086b76834b15d1722a92ca2d55807f2ce128eb6d87c14966d1885099873b9415f62d18eca37d6e72985094a23a5f151cfe403c4b7bd04851d59e45c3ac31ee81beb0f9fa43e96c103;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf400989699e206542a9aca5ece591949ff6f91eb352169e0bd5b999673ab5bb489f65e3e92c35a2320ae48563d8d8e315f3229be447eadc369d6e700dd2baf7c44149e85947d6ce30eabbb8048899ed26f9cbaa14;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5a4080cb568cde490e64358c53079ecdc72a6b2d2adeafa6c1f2ab9720bed00b87b32381676cf0c3b2f7333eb5dfdbc180de4975f698edad44fdfde35624b382f372cd900bed9bb00ad0e6ef1aeb5d4493c1daae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0552a914f900fcf68aa11e686b6af5249c4a411b3916134d42a7bea9ea7633bb7fb0594fa4604ccf0d238b6fa6c3e2711f3929709b50ca0d8c8a41001c4991bed5926f0642338e9d509669126966edf929a0b465;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd619876d255de71a98727e7ad4c220869a6df61a49217f45a648b75f60610d0f09816a3deb1eed1fcd3fb9f4b15a17e216b5ce89fc51b14f520b8060987737405f73dd93cceb3f455ba33008bf549d1e170363fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc307523f9d46fbd0457ef4a634a0bfd405178474cabb5bd2471120f5247c8d1149debbc4da374e571acecd80554aa33ca614a77d333e7a126b39d2e738301523a8703415d8d8ac4b770bd70d9063e8a717f1de346;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha488a1d9432f761314e40a45709399ccd98bc5b223a4e334f9000bd2bbd4811db74258707f2831f3b6cc1084154301e597b037ecdde870881117a05a25e2deea72345314fc7a9689d53a6d75191bc693db3d65001;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94d8a1de8cb87ebabb8e7ca5f859eac5521547c51accbeacf158ca38b2ad96667cf1a2f71797562b5fe2d01e26220cfbff09ef1573b4b54fedafc1ee00371f1a711c855eb4ef17f6bdd5954f5be1e84b12587e009;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84244a01c21b2b12539c520391196eae7fe02e6da7baa0993cd36be880104d46f72ffc303c2165994df940c7a089830587950fc3e1945e96120bc9c00938d67788f7a62421e00cc0f0ffebab0a73e820d43a02f68;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1e85e9e7ec0a568454ead591a937502ac013dd56155527118e3203791400cc8e2e5c9c8c71399499deec6a1220ef9da602a62ad6e1c58fbbbc3ee4b018a23b565c6a0d22b140ae45ddfd14c5ddad90a8f8eb54dcc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h67f25b0fa45de663cf16e20ad807b85160b269890a3e1d9a572c7186d892acf1bad79b11d971d79a39fe583884eac51a96e30f2adcc2089872bb01b2e34c5e6896f124b44c1a70a78b81bfc58094d779940e43704;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5df4de0acd3c0b8c1247252cbd169bdf0b2185a26bc45438bc2e906d735c53456a6aaaaa0510d5bed069567ef17684b2fc367195064e0c3baab72cee6d09ca7fc995ef96cf0e0f5940d10baa03a5a6a6a8fe13931;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a3cd9d8c2230617b9e478579f601b06e49ba7f3282d59926634164836436517675e93efed3f49369faff01713cd9e45e5c912e96f0226ac1c32bb354fee3d53195ca623b45485d18920f61378a5313d08057bc0f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6bef270f4cd12e418216d7f422351281f55de60e4e5e32f1ea32feedd1ad2c09063bd009bafc5b37e34e987d57455f6c2385a65ee8a14b4a3a582da9006cc04454b6a92137327a7639c75fdab4cb780ba419d39fb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1b320449d0a763ad5146a56b408b3af6e1a6bdcb25c9125f52fde3aaa8a60e9fba96adbe5a59a5f82ce2d127c31d12eb334304f0fd73d157d16e468e8b1bbc8d37ab1705e7c0747f4fe2d41da6f8db626e8fb5398;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fbd5012f768642e0a2c25627071c757f1d8a23eeb261a9b41f74a14a7542015d0ff8ba81f07b18d5cbc49d37fba2ebc3328d43559baac9c9bb44ad33351bbd9283899f4132892095f7854ef00db111dec5ee5105;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha873aed2c35518c885dbdca484d59e225dac93d35545604f1b06a76950fa7e4a02a7fbde83f685a5a8b89af225292212bef37cb183fbf56ed9c48502278edad5a3880e20043b69e4d58c573cdb83d7aac87d306d8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb1a66e4102994c87429a0c569c86b7f77afe99b0ffb82dbe9bf3ed6a037bc3093ae5684f1a7abd137e374579464b35a116894d953dfc45d4e9ee0b5cdddbbfb367abb5be0bc10bf793844f39cc16abb660daa323;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71ebf2ec0b17ab5448a5170be7b2788f2ffd071b0fba42cca94d595b7acc0ff78366af58256af94cc7512c858dd8393ef6fc2148b57818262ef4213044a229fb5eb6ea661ebc23b238f355344d85901a5aeff40c6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20e8c18c3dd21e2ecfff44f89acf80e9804fa85f531bf2776d46254963f4ef71784c51d085ccd0de1014c66b31057303de56fe1b47dae0cf39226d30546be8f522608cdf160875a8babcd6d6333674403f978fffe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h84905d96520620dfd44a5d54cdd260be3512dcc59ce0f598e0662cd87965d0755abcf016518066abae662bf571ec62ee20fe886dd789fd7dffcc982ef964d14d5809d695bd9183ca6c7ff3999440e60232e677acd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h535cf0cafd3304e3ca69a8b061828f53e515ce5dde7b187059f200814c2f8fc3ad6b5f93b06bd4d323b03f719e2f96b811eeb9b646e602e84c7bc7e3d4c848832454f515aeb50a1c873b1429e560c4b26cc91d684;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hccd76a1b2d676e28968ee482c8c83bd3c963abe95a9a5026de7fec78a95fefb24380d833b1b27fb8f7a54211f7f1bd86e3893538ae7c7149fd76c284c6b321e7c65d58cba3defe6bb78c99de46438e45f2617b275;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f502e461674744c8e10bb993b13004b8edc4d73ea23499aa913a9248089db1a7a986ba88c5c36a5184f623fed1d6ba4da7fc0085dc0b30b4b49afacb0918db5746749a9ba208a53c127d630aaed3ecaabf356472;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b294519c6ea11bf37d1d460857cdca71cb261eb1cf848f86568447679f845f178f40db1a36cccd9963b939e1307a4772200398d56d1aa55c147289907a205d93b6a4d4cc95a60b12638921a1c93fdf1cee03dfcc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a76e09f11a96059b77041301fcac579caec82360c3d2a9037a535ea2a9fe3a8a0fb67e3e0f2b97bf7155affd840fd5cab0c09775320803088e3791e97c8754c93297243a49b7e0e778aa2eaac9703a0d5b4da9dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc3b4eb06a4a37ddf0c7de40d33b6001110651f81685d61102d432f51b7a92a6f121c028508019defddb152ee1a0bbe8de571eb92b2c7cc4d74bc72a8e5ae966c7264d47134a7a304918247d6e5900b73efadad955;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59ad6ca2be208f5114b58901c2c19517a7272759912fa4ce4f1c591e5a566cd5f5e8e919d9291b2b99bb4656ec0224b885c8c46f8454b69d6c8087e67d2f553a22e5f28b74dcbada5970aab13ca3505f1835692ee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf858836c816d5b9a28488cfcf2bfb9324e8fd8b445737f13e5e472e6ef7777b26fc137964f2107abe7a4f315e43f44008f280047a99230a53273f84f44cdd3f96afff444d2d5fef84834f56b50b3b2d716ffe3db8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf0cce0326cace8f27e85b7c981a647e1e6d9a92a001c3a50fb46f909ca2b6a97e2abbba060e7e94c87c56404b1b6c52cf0c08ff405ff5bf911ef36d533709e01fe6f305cb585d3b3a5cea6ad133b3da85df373ba5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h185c354e9ffcccb2c79749e25b137512311ce0670ef011b2c001b45187c6cc3784614bc178d73554310e39ab1a23b380aa9117e2b9bdae79f5e75e911399cc04807f4247df2e8bc0ea88c2b2cb4837bdedb21fcf6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48ae688b58865ab74f811e9a5af0fa2408e482bc41057775b52a43d2df63e3f8bd443e7c5265438c927e0ed3eab337c85f8b61b96993f11b58f1753a38f42a4da355434b932c08fc0c22365cb2093bcab7b0726f5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68b9a729435a724a86d1d4b3dc0714ccc926911b0bc9d5a3af070482ad74246504483bea0d560b2e11b4f6783d600b72912dc43b442df112c64eeb729b55d4be61aad7f2fca578c59b97ec3fef76c73f25a4abad9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hafe9b2ff0d8d9d62d9d842b9b00919909155c0ea54486c4d10cb1167f7b90310e07938cb5961ae16d9e1eac04db008f58d055b93bed0912dac21581dd0c43dd105841844e4a2bd15a268297544ff70bd2b7d985fd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb998f8e52f088e244eee759e82d7d1c3a839f816788e5c718c1c3f409f9d2d2dc3e0a6554dd92c723afd96d7fc3d71d3c42465e86f08eb91422e7808cc68518a0de80046414a071deb365fcfc2214a304b0139453;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98b3946fef4dd294c33ae0803813e580672b5e5f24b410103f1ae1c685a8aa14d16be21bb01d88ad43433e84b0cde6f7529d7e6d9f92f3b1bec93199b4e65b150affbb83f60e44c654d3ace2c29171fa6ffe78ca2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e795f6168c844595aa46c4775f9078ab0b7a52974b987405b4020e956fcf25584c0f28c5d38bbd024fe665b3c7281a945e910fcd00ab8fc203cf44e33927034ae54a48748d7957e54daf3970fe86d2965fff0797;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0041f76b97139a150f256b7c8f811754254dcf592cb068a2d1976351d283b92ccd8b4fb61ff052698f144dbf70c0ab9f1170230eebd38549f22049242edfe88adddb6792192c98eef18f1b904c8a0df2c11af61d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99dca999791ba2b6d6269dbb8cab9896c1c8bfe69f4492e45669a9ffbd74ed22d363d1b791d06f151b998b145e6b3aef5423592343f5f198fd511362939b5648d5c18d57e3cd0d8af28341ca81a2a2c9f1b80aaa6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbde75f0698cc2aad2d52b9bd14b5f4f5a10315d55816051017e6380db485c8466e0dc1550abf0bde17aea1d022fa140ca596fa066b96eab20c04674d15a03397238747cb38fa3f882d77ea31ba3ab09f176112e81;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6cb69f3b344ee3a69ec0181594c55c256dec36a85d409099b9d7fb19ed49f859df5a3cc941d253fb92474e278cf5208ee29d23e2eff65adc34bb1efee31b818e8f063c386118d9c31cd36831ad84aaf4ec27a0174;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9731720dfc70c983ed4684459cf0012da7660bb620857f3e570858870f64337f515e9c2a1ed1249bd23691d4f5f653153363ecd02cd5e525264f53743ad1a758595b4e32101e378f8b88b67916381971816722b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff3561793e0210a436d1275d663be1794ff73d5b315425e2f6e4aec24cb275817a9e01f0a09eb5e47f80e6a0d9d1b86d48f9dfb89de4d84150540b5a473b48002d438c944d8a77c142e0a336909871b201aa645b1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9be6a201a7f286f4e88d8326dd572c44b05bebfe4391b5785a520262a146cea0735f7648c302ba18b4928a854ed36e0fcd72e159ee98146992b2c4bb3a8725be17dde57e6e5d12024bf057e020f60455929135967;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h21f1e565ef469fa31ff3467d23ea61bd6964a24c9489f84ad18dd2d36d6db78ebd7cc9febcb7cc3061a68da1678d37f5003c437175d9db2d061e8e75b3e4c1d2dd93d321396516edb974fbde84a20499ad063e925;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c034cc10ad40f6bbe99ed4d2df0a67a77c832fc9c42d123d0116551b99dd7948d0004404e244bcac3f44786bb8f348eddde52173a0f1c389df0a6985d68631154a9b48922b077ddb5b990f7be2af925e48a1967b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2de6d3bae81c6b088d94087e70b6e8ae3d0e330390a69c98549755871e1d4795d686a2bdeb5f8f0ae5fbf61ae3ec4ce272e03e5659fa465fafc1a32066685efcccef280f8cf5bf43aba0381df48468ad1d775fdc7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf37b1673065c30561d053f0ce3fbf1802a99dc5d8cb22b4bb18b9879cd31a21813b62447bd13678b8c374b2114b4c2510c60ff34553351386f6feec8256f369b8ef5c77ae734f2ab2cf2727a638590db8faa33588;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd416da6872e2cd5ba01087716df8cbc1c153e97eaf9085d56569d781a01b5129c93773f715cab82793df62d02df20589b8f43bf4c6c53fb9be7ea17f82b8675a1a5b77399b102e142f86c6028e110c380c52f575a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1996104703bbb161e09a98906dd3a3b8aa94573f91c8dbfd2172f50b0e4c64abc3bdff34992ef2901655712bb9f91cda502972b29eb6ac66b93fa93c2e77302e56fce7a9ee2029c66daf3988ac95d8b80a7c77ab5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8ba4a0afa5ed33c1bc10ac7905aa74c6d0bf1cfba05a2f43aee10d8cf65ae43d702df16c99e43fd5a8445dfff048da07f4ab8be5d69822dadee634edaf4e49630458232f32bdcb2294e504491d353b4da733fef96;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h461d0d0de86fcbdd8f21b044b60f0916a01b7f3da7ebfbdd19c36734ca1ee057daecfc946ec78c5700a581658f0989476a10399eec341f1fe329f645e6a817a54a3648d2afa7e2e9388ff011d3f699e6ded897c7f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bca74aa069d5bbe3f8668584633f576c813577463f4965104a18cc749a611afaf771a9e561ec525874b6b053de4a13c32386d2216ea150327d594fb980772491fd1f25d6aecad23ad5c2b578d77a6b0bd5ba2e22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d67ffe653f2f291182c1862dedbc4506416dc941dffc84ce21959e736c3241c8e4bf02bfd90e77a2216345cd4e672b204f469c5f99b6e4081de5500493520cf23d00384989cc53e3cf98579f612852039cbc08d7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1370f1e1211e26b571d405c16929cd40aee1c5a2c3867caa188eb4922f5a2b96e58a42491ab087622d0b75b2f472418c21a87b264b9021b0e4e991526ab0dd19a0fe7d9b249353ad15675462c8762a032e19706dd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea041cd6a6384c9e6336ea94f39764959ead0b3bbc49f53ee1e4dfa01f6d0b326d9be496e8dbce8c0b23cb0a5daf937688ededbf5f44f16302bc17cd1e4127c10236e9158b76805e96db340e20c54dab404a3519e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ef2d271e27404712984120297f68f8b189f1a5180b9596061f1535e3ff4be398ef652392c05a20d7b45e9196da775b32168552e02782f7895d86a7523e8fec4121a57bbeaa5b7acf01f1e37ea9aa6ff4513eb8cf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a92a067c7bee82a8c9dbb6777c879d7353e0df3eb6afb3c5a6cdffbf997a6549a43212b32f07e5d1639c1dab98f6343713bdc06b11195e4ffb2f922f356eaf9644d7d737cdcd47a92df5f8b5d2bf2bd9f499c495;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdc262d48217ff32f3f88ea41b0a815531463bc29c44e0c0bd3b500c45ae603faad792e417079e4bbc678ad974a80dd8ab5abb34e8744d1159e1c39b4e779bf0f886a2692a3b9e67a6d695516d06f8c142c3fd8bc2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6cc7f93cf6e7d466c58540e71e6a7316d913d316faaf2ff2671e722966819498b1b89b2300afc296fc6df005bf9e1834ed2b26124019f7d08feb2b341b242e4e498972857ee3725f6d3ec29ad4900697a39a814d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h35dda67489d330d3791595942da3f6d1eb4c968fa41123aa2173a3f4714793dbd61c739c1684933a2e738cb709d4272aecafa1723e4f97055a106bff468f57fd116cf69d18a83454f83d8c317b5500fe60736edec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb97cbbcefab33959b6980c9af188eb066a0c045dff0780196bcd604990a2a4d4cc5c3934e6f09e05dd2704f104e7e3f8f9f44f7ddfaf625b21d5b834452547f2b037455f92c7b5efae2e8a907817d0c5bd16e55d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7bd1e962d951a13584936ba2e92488f9da5fe674c0a13c978cad092aa0cf231739e5075e422fae3256c3f2644c60b0ec8d85d348db48fe1882b6dca3fa02fbdfd2ff4f0fb4fbefbcc2275fe4fa494d8719156267;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6582daff60d2d94ae578860adc04dd9bb76ef2a73e643ef109c66594b6b047a28842be88155cc1407a2d1ff4fa20b96d1c01979d1c518a790cf1603778f89e1ba38ded13cff4ad57992916b804efe986b3236e669;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2309303fc2fa52f8c33d11d34ec6f2b17f29cf9a067fbbf227990a2b8e708b41d122b1298aea1bd162a5c3e042f9b99db7871b9db292982007ebf2fbf2b28a8c7dc7531e3612008fb51948fc02c66bc18980718a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfb2f4984acc67b12b541360ae29e0cc33d715c805a8c7e05aad3152c842ee99985171378adc38e9e03a89e7c2a638475700aa7efd1f5018c43c0c6b2b2be0a5bb5cb1e1406d87bc5579c7d9825c4ae5f9733f1800;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h835cfe59438462d3a5f29b07d2de8baf323e8ab81dc452be8469beee6d38ab0dd1cec6f2b308ac181cc8b4ca52b8e767f7485afd2d5a92943563b6f0f461b5ebd3b8bf98beca89debb2f5967665fe3cc03265ac9f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2645d7f34eb4a313b6b58f8f098d9765a2a9a2ed33d8904295ea656f94bc457f1abfe6cf990cbfc6f5c624b42227ec65272aba9042252461134ff831a1e21495a039b99a9ccd65c0e2cf8d06e480f9c873001fe0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a57117390ed1faee9fb9f2ee29ae6359e1ac5ee06e2b56b10cef0b07cf56728b1494d4d592b75c16dccb3b478da90522cbfca046a926066c234e7c863f8867ca0786e2571a9dce21f2d1c71ebf5acc512eaa3817;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf2125b44961918fd524f4e14cce9ed32c68d526fbf6b623c01bcb9131725c58eacded12d0a512a69c154367d99d36776ff54dc7a98f4a547a485ad525f243c9593cd1ea75277a7fd66591f7b87127838c7089ff7a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb21e761a993b8de671ba112679f5ee796fcaa763a538203176de74d580f359b3a5acde9adf458e7e6e7392805e8d805afbef95d9e6705c1ed6b578c7f28c249b97ac6a0fdf71f2b110d7b559584a50177a28033e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha32bc1f9cd7435939ce03398f777e8ef2e49643b666f879925e5ba0720bff65120605b120141ec703598421384f7929adeedc46ff582648dcbce5b278792ad8643d68143b1f2b19591b19df26f6de613ed30cb69a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hce7263cdcc6f5651ba11d76bd030c5f10ad85d1e5bfb4ab5fb1a88d0b4e4a88b59d29da0dda8ae3dcae176deed62347c6005de4e2c32766249209316e252f8e91bb54b24ab8141e772c4fb8c45f0c11fef3f23463;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85090626757c0c7cc21d941f064ad25bcd344f9575189ecd7903035f6d748f6f1481347beeacc7b60c38d4e0f637b41d38d802fa3817ce44e09552256c0bcc0985747432badec1c3b9c099b994f88b443c0007ec5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f66dab0f0cb210d413ed6ad9e718b371a4b082fc7c8cd4b48ba8459475a1c01dda130a2efe70e73d3afb98fec1ccb4d6fdd5e595118debe212450afb3861e983a274185a9723ada7818bcd92149c5f3a239e6340;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h95a63121512790782078c88c8931f799411a15d06abf69a8340261d036ebb1ce638c556a124443229430835ccb85da5a971f8c438844932be61ea8f5522e8c83d51ff29a5fb65ee8fb9ff71df0ac651489c2f92eb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7cfc54068fc2d9cc83cd337312818e6bd011ad816b2acf9703b4d2685058f024692b7eaeb88eddf5aa73ff53f5f002858758352e2eb8a0a944e3da90601e87108d99680abb3e5da8084c8731e3fa7e892fdc822a6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h171fe7065fdcb607d0d20145c545a19815b613ce266fdc191347bce1ec3fde007cedac098dc0b29d3137b0289a864efd7d52f8259886d80a804bff8ad80bb2fbf76c839d32b2e68f892728906efd66045e6d96a38;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb15578ed8ee751871f189272ca872e55790400f7aa2dafcfc6c0c000fcaeb0d78abe8cd701540bfb93f61d16fdeffa679380319ca9f87d3090d78c2a95f517cd6b6d5e92d268354302ffcbbe56dfedc054e3db105;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc22fdb76a90e90926af4749932dc43f1a042e35e90d655e2fe5f3dec8d2b71537cec4e12d31d136438fc5a6ac48ffc3e2ac66163c8b2c126ed3a8593e53bfab2ab03c1ee767b74b91f3c28486212d3b932b7253d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2cce28405f28a52dad06c66b324e3eed9e923c721c18ef1e4ce4f0b602d1b8116c32fe7fa20972658e7125cc1f9a47f209a5b1c0c469b70326e3748f3771e3f732e574b1b45c3c6d8831e55cd0c832542f4200efd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f2c4901d4a8a12462b9faa012c4de17e2bb28ce687f7d575b833747c927505e01d308de040db56c9d97acbc9df95d0771ac0aea829f7cef83e2c9b987d5fb71059a932d49a3494889c9b4b8f2354eb7a69485fd6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3962d0e965cb92342ba15c3d90fea4026cac1dc52a7e38ce6b635b267f4db4d51047a34fdec44f36c2607dd4f4971126cb853796cf21eb12ea82618158323cad987e098dfcfbe6af482ef1c4c2a2c4cb8340345;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdbe1c92597aa57631a744e9b1322102cca23db87f58fe0bc0288fbfdbbddad010f32b371045057a261b3195ba23cf9af66c4bc2bd66eba890bc41771e38028eec413620e0fb20db4a615fa0b42f0fc709275747dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b5101ab1b7455878e59555c6ee5565bdc85ff1f73a2ae634d9a294baa1b8c14cbeeaefa4033e52d268769b652296fdf8bd46cdc55113bd65694b43a7b1f02a836b3ad0e0ef118ae66374cd25d612b8ed415000b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb0145c9b510b26dd603163091c1e6f6329b04c868e4a04d5566d887a5695e34df9fad8b22651e4e7202baffae9c7d7f7f43583f74829151a7ea99164a5ebbdeeb924a7bb63c0803d9c427a2927dc2f28a4338674;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ad0157c229af3fa31a7d7dca864b8c6f504b25d9e3c143f89954e4d2d839dacaeda0e1dd5da9e0b2c8ec73ad4aa278eb0aa8f5075be250782408215488ca3d135adde19576c4a02544ccb0f4e5c720cee3262aba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h98e4d3980438f971a6a8d985c42bf055b901dac36535cd23661d18ddc7c11cc9ced429714ceb57e2d1a050b63952cc63325c428f38126c4e52dc62657641cd02c482a3b2b0ee19a6b9a1aa1b8415850ff05dc12c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h747664ad16d699d7d9caf4f30c80dc6051f5ff7dfdd9d189fb7d29b00a6b4023c9ad917555f88bde3e326e40cc97bb92969361b7d337d6d8db959b25ed8d062ced312869d889d78769376ec9c9cef4da6b2cce3e0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h253f5f16814d2cc956f2c4d732a09cd62650b6b8e6b9d2ea2da78365679fa86e925c963c8eb925a3b2ba529946e11b587ba032caf308afd3aca5b4ab81a8dc4bea318998abdd9c78e8d71e558f171a6f47a538243;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6489bea35ccefec82007502b3019288ddc58301df610e2d53b1626e43d8a2b3ebe6946c4418617e585313b09ff2cfdfa0ccf697de742cf61bed3a9261766ee9c240fd37732b2937a498e3ae1eb15b858f33da3f55;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc0d8c0b17322073a5baa1010b05120c3d035cf8bca5a9a42b2fa1ac16a609f066c449312493da2463ada5023431ed230687043b2f561ef19d4503b0c87647741409d09f5dbe32091d27cffe7eeaa9533fed98f109;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8fe4ec54f541cecd455190ff1d102470019e06bc7a513ab61c65cf483fe543bee4aa32736c22f07c75c29995c0c6972e0993938e608100574cf819fc1df5a8634403e87a3c75290489a37ffd44ab1b2f3e8d4d0cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a694c4a9792fbd53b12ff17a4fe3156a8fd1cf77f9593d6ead6dca8de6aaae5c0ef526cc85bacdeb44d41696cda14eb1311ca69e989805f6a686f190e7b8ee5ef979e09f91444084a1f4c5afa908cc09946c04a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1cd162dc3cf1186a1a49d731738b6623b05762bc169413228ab4fcd8968df6f5dbf2ff4d7f159c72793d8ece4187725fabba586636940308f6941adab75be2a04dfb27fde5faf2f49524586c4c42f67a719b9fa34;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9f95b0ed6cea5227c6ed5e65aa593045db8e4e0f87c17d4b8d52451c46c16580d786dff68703f8cd71ce0d5153b8dd376612a60353370d50fd79bf2f5df00cd20d365e8b1753ce1f100f50155d4683c3dc9721a72;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb960c1c339723afbc50e7226adcc5dc96c6fd377845548d5670584bc9d72ec7c28a509cbc74fb78160a7921adad82979fb74e630f649f9648dccfd9a0d84f567874e38790f300bae67328376194b905865c8befe9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h917e53918093a95c6476dcf051c80f685220ddca5dfe2e2ecceb125ffc6bf33c3964a03feaf176a51a9da0fe1ee539e8a021a6637695f3da63f3fd4d1770b74cf4a223a8b25f832412e4b46443b257c1f75b1c299;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd88516f30e35741747dee74b2fb081bc5a92e991d1dcb92be5271258db3279c64947a9c831f33ed17eaa768438b6ca974159141e675c4ca5e6951c9f55d0c2d176addac6536e0d73f0a9aa4d46088063a8ef91e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h72d10577c17b4ccfd012667764240c1ecc86b972d32516f30f41d4a233035c9eba3204cf48e3109a9eca78a7256bf588855cdd9db6152755e94dc235f0545d4572f084708d10326fe33064e34bbfd76ca583573c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2e0ab22fe94416030b363195182ca6da7418c8cedf2b39b67be73fa9e28f6c80372f3080e2156044a691da68d40f4b12ab1e015b2d912f488cbcb3957800db55bd247479707e9cd6db0ad4cf693278df84198e3e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h61508cb3de774d1737260a327131d193f86c9c21cf6aea1b9103cbc9737c6536b36f3e9d22ddb4158df86da8ae8a1c2a9af0707308c410d85c98311817340a55c374e7e1b2a949842b4ae3cd3c309fbbe7b59f03d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2197d77f89554a0fa2b3071983e56f584e29c1fee55ffe97b04c574bbb5b684bec8227a18a5f1de2e7fe330cc64d430923796dc2f788a6f81ee7a1a24cd800566fafcf9789dfc16f6e9eda62a55ee7d20eb914ce6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70b950ec55001534e8d084cdfcf2a52ff8831072db1e1c9ea8d373cf5a394463981fb259603be5e663eca1dfed00455cada54f6ccf1ac4fd2795f36ecf0d5c0d0fcffbed2223d945c1f05b55b212e4b708e5d1b33;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he2bb0f700e85dbdd55c738b0579e2aa1e6569b1080198c15a4581ad128cf17b166aacb3910ed4c646faa0d61a782a355037e5c1607ae68b4b7f4dfa1daddd7f20082451dbf785bb51145fc275c2052dfbcb6285f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90b7be626b1100c0c66e8ec04790c4ea03470e1efde9c1c354e8846ab4e5aea6e9a1ee27fec6db381ea7520826ef16e78b575b2ffb127e4ed9b9332b9173b9b851743be1b152f08b4133d86f577f6a0ca164cd697;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h672ffc2be5bc099186a3b6d5a96c98911f744467d1f9294098bae93e50ade2591133935b92ff447c8f9e65d90a410d0e2cc8feb29f764ded5312744b3fec75385f210b7c5dae12b00aebf76f791477209d4ac627;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6fc722e362a78e27dec297cb55b26d66aa227915617c8665cd21c2aaaaf2438a04d92b645e2fe802d274861bcd1b30b08da20b20d35a948be66a2b7d7376c0f32d1c044548798ce49e2468335d44d54996dc284ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d3fcc847bc14f51188fc20eb9ef797b9514f759e414d8cc9c649aa50f098cc15edef313503b2f25228f7f5c6453379eb2ee5a96a6d88bdd546ec5210ca6894fe02bb871efa9d324e0b25622ff5118cfa1ecabeb4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17a2fbd74730798820237aaa532edcd52725ab92d40b5049338ea82f57f8422ebd7c07c1ae50f3d2ebfbb5790a330184c5117a770ccfe546c298cfa779877afb84ae2b951041060575944be41a9dd133d5ccb5c05;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h970cb2e95722c238383f68f50b8e8534c82a8fb0e1df3e5d8798620b8f6ca2ec650da6433ebfe0de280547ce64350783608c7fb3e12865f7fb7e467c8ec8000334995e34a6dd1c4092d1ed66e51d4710104bc2fcf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc8bf84daf90e552b7a5d7be7561700c08c16ff8de14c8c62cd8393595b10c9067b945a8583b58a9ce0c8589f32c2161d107b9b79e11fa1e34cbe80e5206073c427cf70bc1e1d9438dfb3b218a31e6306b44316ef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c21258631b05c01240edccce77f0fdb922559dbc156e7003c4390cb74db429ee92ee2fe1dcba844064799f3599a58470c8b20ebf6f8e440036443f3af5769a2b94fd1e8fa59c2a24f42588b6a8d5a1d2e081714f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h20bdc202d9ba3da5535f6a1a4c69cac673f66d99282c6351e036aea86f18e48361e0e76d620c7c582dcbd6564a4cf693fcb01de3faa7cf831adda7e3314a8e8a547b204ef26cf5db9015c7d1654fc8ed3ff78c35e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c409a131d2eec18f594db52b938fe61a0ddb3b8a625cfcdf70b147591001df8542feb1cd7a7fbe496fb1a8f88fa58519d28a5dd28989552ed8cebbb6efed15c6b2c9f7bd3f61b4ef5449b12c48c4a9f20108b3c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd1f9ada50c4c84a9ed588c7b563e0a0a83b252d2cdb8c1efbb407c5c60b3b5d7e4b503e8933aa7cff9599ed8db2940bdb849cc6cd1fe730320c107cc8848f0100e96249b36cb954ab5bd01703466ef00c754a1767;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h704ef85cb6a20016bf7db89e2254860f8bf4d5782eb97eeeb331982be52db49c5fd4a4134efa64154b701b986ed2e520721ec01f7abbc6303b6f0f46a9bf00f72370690547815ddfcb17c193b447e84cdeb5928c4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha735b379432e561b4ecdfc0f0a64b38c7da70d84913127ab60099c8346d3a3dc298cd42519e6db5a652ad43c8990acafe4523fbc90fab8741b9bcc4ce0f6c4ea516a5e30576c9e666e12f2f8977263f21b95f7e41;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb783cf20229337f6e5e50ec1d0c0141b74daba2e7d95fc6d836885f84534fae2cad911e62024708049c1906c37abe75713b17936bb09852d5c5eafad887d7743f85ed6b14b948bf574ba97e1d92b89e710a9a908b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f8a660b7890b3331bc1b1a97c53a9352e9d5ea0171a6f5afebd576c91bddc41630070f2ad516d30707ef17d641f4b9a40dd62bc801e3af7003d475d058827134794b0ababe3554721dc1fc1a57d7d2511a418d2a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c9757895d6bb000d85d66401e593431d65b3c570ed3147a10aa50f2708a7693a2564d9b9709c7faa43b10759214f5b02ed3e69f6845d22e9a304261f0ca62ad84e818bf0536b8e5dc94239c4920fee120763191a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4118da1fd8b432de6c7a3d0058bdbef6ce37457157646e305f28ce782a5f20ef2d95ffe3acd5e61168203359ae27a3eda131a1ef036545f87adc9a6d2d675fbd1fab40c8bf946a6673af69690935b3b8dcab7a016;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b83c94072c113c3bfdd9ad1bc52e7385e845463cc3e1745fcddaf9f2ce7f1047b6f714ba0d8a573f4c80bb4f6f9580037f69cb696f0d87dbc0dbae59f39c7ed7e96fc89677d7e19a99c2ddcb91f4d8e3593cbee6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h787ec4749e4356c2653cb6cb79a977d235c5824a0c164a1337a0f7c823e3f15218d4604352f14f9c182b6126fa38efb25d6283a687eb2b0870cab7e78adc07ef8e5dca7912458446c40e8ca765af8ecbfad86d92f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h720009ceaf108fd9363139695f65f89a5a0db90477dfb8c749afa03b459a5761a62ec8f892549de122170b4f0ae0bd6849198860108f78165891d43bf3b21ac84d4bbabf77a496c0727c2cfd3cb011ad5616c5460;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdbc6164f2021e6d68fad94fd53e2da4119e1b0d31a40ac290aa10d4c35694cd84d617d1a2b2fe62eed501edeabd624239eb8069c97c0ef8b6266877ea37f614cb06b98266947338e414522000f08176cb76e9473;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe20d12e996685ca38c408fc7a830720751b00aa4af12ef5127a2b3c1e876744993f99e123e76442ed33b923b44b60960dbccadba150b30e15356905e83f202ebdbe3fd70bb1d23c654d29260becf53255174ea2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdf85bc1ab77c9cad2f24269cd1d1bdc76c0d6a2ceaf8f2f86a60900c8f90f2ab1db773ca8fbce8f11d2dc972da7dd0219c18f97c21289280e6d9193ffcb4294c33288aa7224eeb1362d2124e6f1684270e9acb1b3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1884918307e126a962f34b1138319ee69ca9986c45d4c35d0c1c4eb60cd1f5c630a75b4eb0db4ba4d2b2c3fa5c671296c489a4d9eaa548eb41cd93506c52899ca5123608aae7fe3819a083d6352cb08f2b927df8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4124a7f2141d2be6bdb503790026ded2da47badc6b72a4ef52829dd0142281dba232dfea8df5edf520d1a661bb668207da58cf8bce0ab868187d0680e68ea9d8ea48adf5d31d51a87fb67b99f7716cb0a9ec59ec4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he90b3ba8330a4957240fbe083d45c078ecbf06b3fb7dfbfd24cde1f5b9c0d0854dedfb4fc9695370565bd3ccfa605edf262a25b07bebe1ce866a5021ece68abf8cdfa95f8b41e99e537c52301b4a535389eecdde;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h964215194d8c02f911506c23728e05824a8aa422a970d7315ae307ddac9cdf0d86c2be826eed9878022d1840a4183b456417452e8410f7ff248cd4de56696b7fb976031a0219022546268d6e8a85af86dcbee9da9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h42aab8aa218af7766377ac61b08bef3f7ac01072ffc172359c2adf643df0fea45ee2ad1f47840710a5e552eebc7f5fff4e088e01328d6843e56b82e958dd78b800f1ce864073ac8a0586bd43027f14ba81076fb14;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfe38cbbb4a9ca5db33909ae37ad0a33e1ebbec8a73a05bbd268cdf73d3c141f588ebe3f6d11b61d33162fc01a37c92c90ed68c4c0b97a4172f9b048fc6a2b48d3d1244edd9d85033eabf4eb050b96cca76e96aa2f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6028d4eb00f0be3de30cf4e70a8c8643fa6d996c13560c1627fc2e519e1095146aae52250f12671de558d2196b76c57bb1a951da9d25e778d0feacf82a3e576403bc0054dc292f7618cb9956ed0a47e6029d5b55b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64529773663967432a26aecae8ee553af031a69da57122800d0ac64cfc3d15042c356d44f554aa2909dea77778e2791ddb29b76d4cbdcf50299a07abc1747cfeb38ac4840518c47fbed17afa082e393b635e7ecfc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd5bee3fc5516a91b783d53b4b0e5a41c19b4ed5f8e5a5cb15fab244d1328ae2c82c5685e806299af1388988ff62f1ddce8d11147ca8f923c8f5c6d85843df600883923f912348cab81560b49595c8bcf8c5b0175;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8b9e60a0e6d5ff201dc3197b9abdabc61ecda2597cb7068840f1e445d99a01eab8a3b7a9efa5629418ec1f9b779c914dd5f536ff9bf18a9d7a48f136b9f37d4195d618d3ac3e3175f0fe6100301f6f662a7c379f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee75c1c913196545c5f763fafe54cdb5cb6cbf74dd82daa136cfddf2bbbcfe27982a1c287ad6ce3a7a16c94238602daf7db1dbec6ffe638c7e41a397edade20edcd010baa83ef10e96d10044f11ad6f83da93bbfe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h172e15f4234a25ffae2756f9b5cb1b15d7254e8076f23219955c7abde5e946869aa5e6c554263aa6231f527dccd565d4295d77c77e9c7bcda1486d42542ac80cf16728ea3dc3dc6e4353258e692b216da8f5faa4e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h87e3039b5269589b6a27d3435ebc643bc79576f67e15d5fb0990062b92da0404f2a060c9704f94d3eeae6a906c6b32bed350993b085e9b238935e9ebe8e38213f1233ecabbb0c9e209b874be9bd60aef91165fd0d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8afa51ede3ea451fe715ed0e25e17194f04707e78544a034e5a87b4e28a4de1f512d5fd60b50ebf02c1a20fb73b9362922c0eec3c4b914434d83bf99bc3019dccbd9c76b9509d32369465f0f08458d9d5a2a29f0c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1ef24bf48083a2494b3654d5e4f7a8d3fc86d7690c61c1095f0aca445422e5122539706cfde43f42da4b9e5151b8eff68f8c633db643fdb78f514ae30b841cb7722037dc7cf30b246126a2913399239b1a9982dde;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hea4be348d3d5392cbe5b2788e8773eb857f366c469a037468ad9dcafaf3a8aad157b5f5bc27a95c3833f06437e099f543cd1c0500af3172449ac1162cf5a1d82ab7d76963bb503204fd0804e8ea985f8e953ef730;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba60a97a26a6a26eb32948d7a6662b347958d3df88e359e334f72e8c6e16ea823f1d71fccfda6034e57359ad912cfcb87a9612e39704fd11a4575b99acb00074f883c2f8959e24855da32f0979d14141e83ee1235;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc00ca161a768abc0c5d3fa660b1f787437128bcba2eee76c87326864782830830da23bc0494738143338b88e044f8d1ecf804ae99e49297b5cb41565d0ad1e5ff9b8c5a3452b034d8683241ac273cbf6c9849daef;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9025308143b03b77e194d39e8bfa346e4476014dd65e5634160d6446d2f6f4d3593cd5637839372f52a23f8914e76f476954f40af35d4b3914c73918d4cccf91575b52d3348234a8cd3363e629e7ee509f7dba01d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1a744be42b7f3a72622754a8294e080675a050b091e302e5ab2ccc87de3931cd5b62ab6125a71a9b870dd95f1a252bf73d471993be6ec4fcca14dfee13d69030806d71eb25744a750249c14d98c6c7dc93cd6b569;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h850592d68ccb7431ee54ed26ee826c97095322c7c5f9efba0a95e863d179aec313d31162ffce8bf48e00bf860c09acf56ae221933398f10fd413179240d9ab4da1f25d94128ee439e16d9f85d2f497050de29305d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcbd6e608e4254073545f780088cb2aa9d7b6d86920611a3d6898382749633b6412cc342a63f873627fedc24b1f278d018733bbc68bbc11fb73c0bdd48c29b4b2c748212129030df5f420604aabeb39d427a5ab3f3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77ca35daa5c519f98a47a8ba602f3e108c9820027ff8c8d4c49b5e8b3cac9a93ca1bdad7d5e06c70e2609640bfd9827674f200fefe0b61b0ac5f34a2a2b074dcea1ec128b693e80d45139dbab138b854815bb13b7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h826a69094b213260f7b3daea56990d847d92c20ff7f7ea3d1cf6e824234f79b836180e41529db8e5f84465884652b54dcb4278753a1784d2864188fb711f6c07a002efde0b14ada57cc2a99f0e4510cdfa2044376;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f11400f1ce867419db5d3f938218cd3bd3d74c5b2c7827993855ccbf9c63ee75b0d257b9c0c81d5c52346f6c7e2c7eb4407cf4e8f807f07dd7eaf37582205e9d3e59d2a1ebb4b7fd433de321a3769eb88ee09d45;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he020068e2e0eca5289f173ee11dfc5fef8e91092317ab5a3462ef22a441cf76fce8593b5cd42df7dfdd8ac5522e5235a70e43809bd05327e2bc036ac022a8c17c08d9355fe45bd58d0d194d04d25351b710014ea5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7815aa4fb4444a1d8d540190b8aaa7dae32138d06b85fd7baeaf46e02762403227eaeead8ae84ac46372b266e5a648c8f3837192e497ef2139f04f9882bd777739d529c0e8aae1328b81713f537e53121a1783ef2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdbb0a7c7174e739f1575bbbbaf00465314d7de611e227629b1a2e24c96099bb2701dee453fd1cb2e7a68746a5aa2079c37a8009e80a169e6dc75de8d56410efc0faa69320b7682fa1ad74229f619520450a9330a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf25dbeb177592a6b72445fd22f58f5cfee003e9dc0f5b4f4b1238938e7d63e7fb1d88354d2acf09060c82c1a7ec76fcdad887cdca701a39da128df4c59c25484404152cc481899d9dc074ae5ed798bece1d615588;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h58b478a5daa25c7259c3dbdca8e48d454295c66eec77f5f0922e5989d56c3eee23c531f13ff1949abe7af1bb616cb45d90afbed77082089ec2d0ce0ee3b16d9cede0fad6a8d61b7949a487177dea4e635d43ae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb67514872c041e5af7a77dda0e137d140a880e017a925bcbf6a756efc57044bced4daaafc176ba77477ff7330e7c67208f241495921c583f5c3c779d90034db305165fc56a169bc7ac5a7a47a95f54405f134d44a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5534bf328c681383f6625ec8eeaa09f5b058a95cbc0eb094131494c291ef287dfb849bcc33eb45f87f6b602290d73df9a4212cd8395074703dfefeb4f600ac738d3b7d6bdeac24fdf61f261df6103c7cf106608f5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8cf62d4589973461a21d0bb2a545812024924cf9a5299d3b53f9db71de7bb8417649859b3e849b9b222b85978b6c2397bec713a24892d63a87a7ca7ff094091754568ac710e52cc53d9baef18e4b9fdeb0163df9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd76357fd90547bb1cc5156af1baa0e42ac70a0879648d2d36d07ca2f80cafe30c72300f52be828fcea63b1933849366b94962ddbbc84ef6f64e12206332c24bc66f458183ab84f0198e1cd60b84c843575704f350;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd0e07146a9eb3ad5a41f4a8708e225c3a294e9fe8771719e106de84602b2a0644acee754af43511aa75ac1cae5baf971dec7fd44fb2cdbeef483898c99bd7b59dd2c43e3d858d064de85a7b4437aabff432b7f12c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2772011cd7d91685bd08a1ce8fafa39fc566801d38a0954293e1899461dccb9e8fc75e90824134e4dc370aebdbf9f1d9f14cca61a5ea7becce1d1fcf2b3fe53ee25bee9b659a539c96952819368a34d680cc7d6f8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b6710b735ffa1658644f5945f282633970e4941f6024ac0370ce640c3652ad0bc896a4ce4e9d0f94ef48625112a6c26b0fafd6fc1081f75f62f2e7f82de0d2a2f815ad1f266cb50b9bbb0a58691dec0d109a754d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c5a5733b800b3010fd9cb544820a0036c6511ef489e1ffd663902ea1b022537b5807205a39e39fbfa4fbf5ad143d9c3857b9e4a831e946c884f0daf8f07921630a23151941944309cb0f017fdfee0fa1239e86cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd99687e1c35baeef8e72c1782979b9bf1f6b87133766bfafa4bd6cca16910aaf15b01b15b73b49cc5b2dd525bd3e2f7699e769b62ebf776cdd386c64e4fa5aeabe02125fe5e7785a8c8d6bb0436ee135ea399928;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcdf6215fee2d6e8785ec738d35d08f2e20d5a6b6fd9f43b3118695998fafca1ec354a32b0ee1927f5c48b8ad618bc37214ad706d3ee64badd109cd4fa5ca99de4595de6d4c98853c036a5c53998d476bf3478dda1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f307a5e88782b4375758dc3f259a1a16bb4d450eeba1d2d8295b63a9493cc983e9176a3dc51a5f25f6427bac710c823402421fe9067d78222f387f23224300981186d8029d6225d07f48f6609e0949734af0960c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6414c29169ba63adf655ab1a4a33d1bde4b6c2d003ed90cafcbb31f6522f7b55ef8207fc9d495a0ebb4eae796770bfa9b00e1961443eecbd11295948dbae3188d29cfd049ba025638521df7adaa724c3411435ff3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a857c235ea44d0fc1eba54aadcffde45ad6a658e865b4e734fa2cfe0e441719ab1f7efedfcc9fa3acf07589066f360342d1f9f7fd1e5072ce8f49a25b30d268012d72fb38237a564abede5af3775a79289c27087;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf20c5a59e6c2bfe61d1e0bf8c46dd31f66d60cae490e5e367a978d483945881b661ee0f0cb46433a539230525a5b2f8287bb559923413a17ec9d9e4329264b8a6d26f35a6de51e93ca2ee66ce5f7f2671c6ec8f2c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6361f02e6129dd647579df84683fe451e863b29476eb7292c6ac0be2d19d076af47e42797d77a5bd9c01631d8c423205576c90c3f9521ee828b3d79cdafa96f7236f26cea3e04dedfeb102e6539bf360c54cfd7d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e9ca6e3319af38a5ebe335c48fbeb474426f5dcccfd0918b723fb858561b013f83d5bd2242cbe61271d842846e6c56e1f6e685e7d006fc31818d4c864685e9b7364c63f3f8cc1a1faa0d8c548a4b5592cb891249;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha22f9172cea7333fdf1a82c4be2444bcbcee837f35fffcb1e51eb49eada99c130a6e8381f3f908b63b30bc4a22835cf1172f29bd45217d93794a58275f0bc7441496a62fb5ff146f4720bfbc5668239db2c77e794;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e262a05a92cb6e8bbad897cc9ca3d5f2eda2bcdef5e3c728b240423a5a5f1a6e6ea8f84b1ce579222742df532e05cede12beb759446458afe06d5c6cc15711c00006e58b0406ec16fa51c73477419d92e46340d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fa96181d0e97abe1b19f5354649dd756a8fdab7836d399c402a219c2141fb260981ee3e526553539220ff0eed2385b24e6f3963a4f89db75b3e576df20ab5c2177ad3d7090cb5a319d8b9d8e32f7de5d78063be5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb3469819ee250b6fba457533b060f8abd12634faa2a2243a799d939cf02fbdc262d108150a2dc4be8882f23bb2e5b05e2429985e83674c5121bc2994a9035b9d9bb7876dc2da02bf9023bda2fd4f01193e92ab21f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7d3f2ce3e619258012d6220022adb2b67883a421108df4be7b5b28bf842fdaa3627625d22add7d1ad0b4ff425801ba2d69712a7dc47ede9cf7b6b2bbbcf8c3e48f04e17f979c281cff86ed2fd347e7a70e14f0c1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb54699be30a8672bf33ff422f6a83f43825444d26957341ea312b9e69b4158270a006c59fcdf801ec722107611aec2bb5eb33f7ac68c4675fb51afa556e3a2da5863afc1da7db71301cf03522580304c4e9fbfa4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h631808a9772942fa220ade15e1cdd8a0931c032be74d686974ed4b6faf436f9b615d3e0096a1ea4106c9599d66526e73697488e566de72d9a63f9dcccca6f19638dc2174dcc47164f02d6a23c03e16161f5c7705c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4843a1a8fedc1879c132322b77bad91ffb78fce9ecca7fb0b8b9825a984abf814598e886373f217c15b3bc3983065d92f8618d81b96b3a1db040e7da965a9854c30c50bd56c15ff80ed33f3a0b0693dcc29e980c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf0a84bb18a740bdb694ec58eea65eceeaf3e3d58b401cd93c74ea434eb626eb495037ad837912d56fd94f53f9d12f1c6bf3b4ebf6c022aa02c56de23efae754b6f152542cf5182c3105bab73475fbd47437728f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdcfc25153ab5044b80982c2ebcf97ca587b32b04ef16172c718d8dec7f7b24910ccb09c83bfd5a511982b9c21a8f305db9cb86a3dc56824e029634c0464dfe91992dde614910c11eec5888356e0c6224582e13dbe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he550867ae3dce8d1c2bf34de988920f23ec954eeaf5dc434c210549fa0c69d1329955736f947c88739f026bb08eac626c321ff53b9b5a940ca08fa07be56ab86f4b2f52992932b3f34f29758c6efe0c06109316b7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e49519bada6c612282188de5df1eb30e3b10970b667a26cf0f742846a2593c66119f04ce6f97208856b11608b7ebc7bef973e2153c75fcdeec54001da7cb45bdac30d79d711cc865a413ef4c78b33abc7d76b5cd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9e8f47fd13713571f1476d5d360715b7ff753d29e6b4360f5ef1027bfd6806a668c9dec477d10229828b1c9e11da24370dfb7ad06e5644f23a2bb5aecc37cbb28a94962b5183355d8db7b1400f45b6f81ebcf770;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha96b6553e64f4ba622b3ec53ebbf1ca9a3168cfbc8eb97bf9a5e6008123133464c06ce756c398f818621500fcba5ea1012ea29ccefd26db1bc81cbf6eaebe60cef5be9f0779bdc02cd71320917658c930508452e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48485f842f42343bdcafca508dbb5a99f9b21ff2292eb4171381a4dbf874e37af1a82d7543d8f394a95eaaa10a516961ac6dab0aa0b3ecd975bf33a2abba743e18555ceab2e8ee40d7f034ede6185da42f81977ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3804cee8695fe88a520ad6062572bd845e2268eda16d705dfae7ae0fd2b6bfe897126dd9ad7c63c489f574578fcd5c4ce9cb11a284c474ae0dd361f060ad0ec56538071c88c2c0de960a4f62761e62b4564a1f818;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48b78efcb17794dab08d0a740afd3c866ac3bfa991243fc86151a8c3ab807208771b4c871512928aefa32fcf902908ec08d77bd3274ed0154e3ac12e4393fafb19a62d6ca2d791ca839ed4a37c2bfe468b5905554;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h76b062860ac5b3075d383f859cd6b72d0d47c16df3b5b463e50fbefc7295e2960624b8eee541e3ac0801d3a49cbad62ccd93d4910baaccf2d967bb33ebfad492fd2f890195a6aa1db71e318d89856e2cca49b6cae;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4fd3ec8f196aa027de6fe64945b56c322f23c7f6eb61046a7aef76f8bd2560e8ac60a748e3a84a4e249c309d432ca3f5a46479eab19c4492a1bb406f7bcb7f799eb7c2421ec653bc55fd84ba5e0d9f6cf38b7f2f0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a3e31a9c59d6e98b223d4bb2576ad562e1e3002e4fb4093fdee25de74ad64316190989287b09bd3e7e675d4f2065ca1793b8f1d12de0ac63db4beb2dacc602c3fe393efc20b034bc410ec0649ea8a6ce3e67fc02;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc84c09ec0a7bd7f9d513436feec731ed90665274e582fa02415d1871b03128ffe02702a165442d22083bebbefdac934dbf7a0beee7c55750f558cb746d27a0a5b9ddd403e00c4425ee011ed8af2e759807e699d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8afb5daedc4cf6c11ff78392206faee25783f801b622f259d79649982f7c8c8357dac5d71b051b46b68cdfee4df0a6778f2bae84d16a88f217bc746a51850b40c220805d487e0be22118c310aac49f40e421f1c18;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h41cb37cc673c7facde20ecb0b1423159debb5b8acf02a696ecb4589263d75e40c09ab6d8ac32cc742d33e94df1a8a3d0e0f70f22dd0fb16c656eb8894b021130288628deb00a95db8d29f2fbc1da73d58ad2d9234;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbd5ab51400453780d8b24f11fe01ef46a22c6b344be2270f0f9182e1d7f08c64a2decf7e81ccc83fbaaeed7aadb6f516fd0d83db9fe851a3026811f1db390b8952fb1e2a5f0b6f410c937b7ed37199e51f4e90642;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfccf15fd6e06b494f5adb7780c1f1dc96e49126b31198f7be56108e10352de3005a26ef1d0da4698f23136b9a84205f5eb3e9503fe8408e267226fb3f2c6d34fa60d68eb4fd575a91afa3f9ebf5677d6bb9cf7687;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h73009a0e18db5ef5c4aec8fb437be981c50b0863bfe6140ff6ae8d7b6b9c7812f698f7e68a9745d6ac54e9ab987fcab1d43a205ebbda5b7e5118d8f5ba12a651cc59d2a68c8a75b92464223d386c98d245bd1fe7b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f1a469f97ca865793696cec51469cc92a93a3a6f688fe9ff806f1ffb33ce31a8483b931c60bfd6b6df90b12ff199285d43bce1c6b238bcf5fd79cb96127d723178ef5c7f4395e732c054df4e358dd9bad16beeaa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbb4f99e11b4a8c2a2b8b4dd85c6b845582d7202aeb22d6294897d35a26ae7cfd62ccca931e11610d2bd348790ef15374be4139f81a62eda595cec3cb5bc9279d51c6c267f2db990dfe499c95f2661f8be23ef0c5a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9ee241e31dee46c70c9618d4db8b3e36313be9e7e90bcdf154c66c159b9aa97a11c94a2979ab2f3cb92c556d20521b99da94691b7e7493c352821efc69103e69c18139386f0921a436959c2b51fb9300a2e4a0328;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4547ab0cdfbf3c1187eb7080f9d3493b2136737f78b01e120360dec18af24de2495f0e62674137a972933e991b37e032f9b39163c3b93221155e32ca3ee8eb8e391985ba5b11818a9f39f502fc75b5355aa2a11d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac400d5e275aec2c605812f6447d033ebbf9ed2da570718493c244ff6eeebf655bb7cb293d9ebe7ca840a3b3b6a089ff3c17a3c3a17a0a58d974d787cf9884b58133b5def98e4caba354b017a6fc8c1e741ba062b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6596ad5d6b312156006a5843ec065fee095a046784eeed5cc1c433be2eeaa2986fda9a012d8f330863d4dc9a24d908fb34667e10f68249db282de74a3bf7ee10bc02230aacce0e31ac26610d619dbeb32ae4812f7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5370972e7bd13d9141b02eea176f8adc7a15fe9674d2c4042b05a24764d9e0e9ceeb0154e86f830d5ac1fbf028db7e9449db434b2d69f44aed0c59bcf1d530387e28c85031cc4590ffb845c82e48754a422dbe740;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3de063c06ff7ad90948d35111f697ec9a6380e68468bc586c581aaa3fe49fb9d6451d1a42974cdc722429d3c1a7def282f740f5dd205d658ed1959cf8422e268bd77e68c701cf0771a6729eb5bdbd7a494980ae22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h539abfea03150236f2cab177852295fd38b731c47e1f11d893e1eb4c5dd83f948914e1006bf8c7a7a66efe52d023d1bae69ec0f9507f15df600d5fe3c4a92f0c7eacc4af80e91854f5b1fe35519fe317a6af120df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h368a15ca5d8de66bf917d19615d7e85a6be6ec79a0d5c0230c3ed1a3c9f48f4d1f3b3f874a1dd23ec2bda109d88ffeb3dd9966a795da18f7271841673f0d69a994cb7fbc5a6329194064efb12f4824ff947127a01;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h147e0f7588f19c112b7c227fea8873e2d8529a17fc669724c481159f612364f00bb5169d94deafadd1b4819cc667055f5d09ed3175e6bb3f00ead3435f3d93a0f78db0cc5a1bd61759ed96445d3d573cc886a97df;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8fde470ab1aab1a0940bc17f3611613796f4fdb4618e76f33383d94a8a4fed99454a8243b021cd9de7fd8de099c443dc01215a5b4c0f8f5b635a6bf4327b80ceac16276b90c589979eaa463197c1859f2075b06b5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha98c26c1c45d6af7e8fe844253150ea3387d1bc60d006b5c329f338ba11247a36df7195eb7c4c49e08fb51986eff17a15dafcd788a652afac7990930b0adb9f51a1053522ad0c11ffd0f281f17ee72d0c89f0f43e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77d47c69ef31b9e89718c1ced531125b53012c11fbda96feb97e4defb6912212e2bc78575323f70110ea9845d5b444707c39ae2a725eac0e949ac470baddf3b086d8637ee2649b0b9508cd325353a4aa80858536f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he15f851051a5483ba70f79bd2ea34659ef0710b85277ba7d71781e0fe2af2f9fc889804919578ac7e68919a34c8b51f13f0bddbe8f39288ec6f58f68ea8a9eaae9265a8f273ebed31c2df4bddd72e458ddf024ea5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49362c1b9911571932da7b1fd6433fe094826c5cd82214b9dcaeeba741af1d1dfc429e6ceb077b3690b789408ee4dfefd89e085b7bbab81b3878a98232f51296601ab48969b416ba22162175c7ccf7bf786fa3b20;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3c7c63a140b7eee2865d6935efc1f6d05ac96657fb9223c5daae5111129f7621a8060b27bbf26cb081a68cf16ed5aa4cd997199ca6c48805e3e9e3a9ea2994d1c9b46e3df30bfeafad0b26f0a630bf5ddd22a09d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2734897e1b41489e50dc3f4d0c1332a84611207e8b4dc940740ee50b893dad3ee8f40e882344c68e2233b33be01fe0658b6f6d907445ee0a819d9aeb838709e03874e6ae14b1dc3292289eaa5563cad60d8ef7bcf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha567ab3a1bbc2de9663ffd0e6e76c88ef55160f227ac6ac825d898ae2849e03f2f9aaae79bd399d27d377bcc70ef50c3519afc365b89b5a4ef9dbc31d2b97bbf232212e83a417ad447547e46da6213d758fe7a2dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4be563b115ee82baaf904391e5552084ac0870036716d612ac04989a054db2b189e98c17d1d4e19f1e22068a22dc12dc3678e26171086fa8a5cafa0f7720a5ed51e4c65045001f2827be52bbe83b637f6a0e33c11;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6b08685883fbd09ba4721901bbb32337302c5e6f5dfef0d936b4051f944f870ed4f2b5ae6972360f962bce78e313195e454dfe1bf5482029e138821aeb84ef2520adf996fa0995dbb0821632bb90e574fc0b6fa9e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacc07c6e6bc8518a86d819c61a5b3b7e933a92730f0edd5da384c65f94f6a846312de039b7f96a2a684acc09b53e628111c7dfea3e8f0d920fe44e16acd3a5810bdb860a871c47eeaf0085c20ce7b66433fa95c82;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47a0fb0d1557f800f0fbe86821f39c9df39067599a0749bc0f7ade3498769e4b67830e9a40ff3a3a547c0966e60d20f70cb5daaf6cdc373a5505f7daf16d5c22caaa9a981477472b957fbfd38f2ce1b3b102cecfa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h17735c7543dc0ecb2262bc46f15c32a1721ebc76721d87e38e0aa5519568f18c9aa2a8a283c85d86cedca23ae620418bedce04bd5b447a12e845ac7adb3151b590744b2d4651c69aef7e1b796179bf6797cf8d9a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he5b186175af138be1480d07e631bc5222f25db682bd9d5a1a1325fa27c61956fad0d6c5c9df686a7539755b582becd8d17b3e8b81da2ae734d6415b87c42ccfcdf84db15bf41ce699cea9ac083b3b1e6b2950ccbd;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h34cde2db2fd226450af5263c7e931d0a2dda2c22cfff77c1aa1ff2f970fec36d49a212f0fea0d16c92322d6f87992d8c795fe42870baedad38e3b9407e0a70a28ff8d99987eb0b52f0ac549eacea099f313b103ec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c70053d80b290f03f162e8fc52a15f4d27bde7ae8e95f317a2a4e1f217d283234b754771d5e8113fd30573d5ef155f421bc180b76a104db75a626a8e775e954431ff0b4c7dd7b41b3186195d8c57003d3ad2f278;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fc0a5964d7beb84d72abbdbc921c918b19271cba4da3932ac7a40bbbf4988c498603474d941700ab9ed46767a14b78e050216955d852537895351c6308215d33f24840c3878298a628b384b7800bef1f7fc7135c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heebac1efe04ebd71acc998e468f9f9f65dbd833c2813edde8e77ea60fa071bd8fb5301931a71db87d52ec8d5bd6a27abbeb99cf54ff05357b083d22dc7b68671b40ecd9ec78f7cda148a15ea2d38b2ca0aa2860a4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h83386eb77eef337c22bb172b6463acf5f85c939ffc80b75b6d7e7cc01433c22fb85ebe454bae0cee8ac3ec1950e4cfa915a08fb582bed01321ec77b2b5f61aecd292b9f1cb8c88fd54f69461f96f85d4dbc64eaa8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fb4a9d6ad0395a245ccfc9e1c762cf7d59819a13928621a3f0a046cce86ef635bbf8dd5d174142692467a512c0669021d53025135258b1c24cb905c06bd013988c9437fa86c32150c5b8aff0d4058be79f022764;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h677537a0bb8de03c934d902c7664205b40eda4d61f85cf7dcea7296fbbf25f2804dd452e5e65669a4ddd944dfd823eab5a191df8a3a7205c3a05d300f1ebac416860e1eff9203df804bda67d2f55a24697b0a8572;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h37c3ba842e1bc4a35e2e4967c852895228e6d80a3e310999e175cb3764f537909cc3345f7df7861098d2284d1277eaaed4a2c30ef339d83335be498e0b03efcd211f22f188b8007d5ff9f23a2f18e187f31f8f3f5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf01de4eb29aa3cab4ba3a3627090d4680d84a95023551b61b12a45cf999bbffeec3c7acfe198f4d96f23a26763a34f6ca343fabd17e3ff1c860ff88ecb8d5dbbd7621bff395db807f2f9e3664f946b8b6479aadc6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1c41691db2ed853b84725861236eff6f56690ca330008a795d6bdf6d761879bd0e982e6ff52aabce5309ccaba2b1034b2324449b3163ac3207c296622b8349b553fb52a26c9360220d9d80b9ba4acecb4d82eeaee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59dbda840025e8a6c7ff6ef5f9fa3cbd583aa6ff6ae5babc5167ea45194e81cac7ac93d0ec2654defa3e6e6dd7d266f3b722621caedb4fd6c7914d81f0cefc3aad0e7eaa0e190462acc2badec5e03e502de5b5946;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb405c0bb0525ddc3d7e57195b54e551a7103243798090bbcaecd5087dfc451a6225c07477db01131085e2da9cbccf5b5b348ae17b90559e10052b7ac65664e7be22a17a26ccbad1f8de39c39439b25a09b037d2f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h939a030b26cfdf0441e8b581e8224ee868135eb7748e0b952d347c5ceaa6830e1f33d11c1c9be05d85c5e82208e03c363fcee20369b476eaaae5f24b8376bbfdd9a0537c5de7fd8059c9f5ec3f1094121a8d8178f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h377417c717f61c4bb418409190bef4945e8b661897067194b46d6a0f7f8821aedef1ec09d696909fcff363accda0cf671519e8c742047455e54e7e16c7e1ca5ff060e48f6647305cb828c21f929d72f01aa553af6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h995fc34380762949da0aeedcaf00670721e08fc5eba58a097509949e8b8c41dc529961a14d06941b44cbbb7a92e25ce2cb685d39911e86d2a4d8180eb442628d5b90cee44a515e25e0cd859934fc485e2a10581b9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he8edb3a2cf1dd5c61e2dacecaf7088e8f5b93e8f04b83bdcc229ba6606c8c2c6209891dbbdf4e0a764470b29afc609359a03445b45530b6c687cb2d2b01eecee48e24bc2287452806cd1992fac395dc3c60c60160;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfda3436de7819014f2a4781bcee031b97d5e3b88da3dd9f36efe96f4458c75492835dd5061496cfb7c0368c5763966296a298e1e4295b4c9cfae3e91fc9d76fa0c0f592a215cd4255e1b3d3e42ce71fff451d3cfe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9b342e1783c798e848c08706a33e0d635b967daf26e31ed219c9b5fd86052de10bab12d60105205acfb2598ed3423852aaaa95ae6a61bc8401535901d78828bf2aff9701daf1dff4ece1be133236c1c2c7a99a8a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9c2b0ba6125acd823fd421b6d3454bc4fba54c0cc4c6e476a8c72ec2e80c693dac9512081e3c59ae27b32e8212520eabdc1061e4ad99891f6febb6257369b946dd5393feaa464f383e84f81aeb40313c006a50e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7c7e62d0413db8979a02f7a66614aaa599fc007f011815c7e158cf8a668af2e7a709d52a36b20b26d0ca25385945e24afc5ab43a05360dab141f511b3bfcd226d2a7e98b217a041b19393680e04369f918334f3c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb04126b83c5e70683f3df121608eeddd84825b9401f3e562c67356ddf66552c56dd2d2d47df81d26b10dbac12f92a0b379e30e6bc47dbe4c2f50abeb3fb5ab08549f84a9ac2fdf15ea0d08daea07e1c1075909b0e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7a6781506ba2c47c3161a709b1e0b56b92f6ede317b15c5aaafa4c7011a5fb4689bc8b25a3396c46defd602d253ee78b3d06bdc023c4cef7dbf1025eac3cd1c684db3ecf56a98d1e7ca2408e8ffbe3eca56d3d9b4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8a9a614fc59b6b84ab163ea4d3f04e4f5bbf5653b10309a4993b173b9027891dcb3e01741ea74078951da707130e3abd15de356b6a573b86a20ae0bb9985ce9fe75bf889bac60205d2f4bb9ecdb961218616914e4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he7c77c35a929b95bf2039c6c46f75835a338f40c7698e841f742afee6b9cb71d91f9982a618ea3352dde9189510584945980286d00d0e0f223330f34f452caed1436a70c428ea7c4a1f7380111014e45d2b288e94;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha49a733289e6a3e3ce3c41151c42b88c1e80281d4eb9f45bb5f6c20a94713744266707eb437fae48669989fd741ab2be304474c6a6b4ecba80d1ce6f6b160a84cb7bcd67ed14b97514f82fda006d25ad428b23d12;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2553a1006897866e9785db05711d2181b00632f21f38e6212f9fc357f0e36ee01211554b8dd558afe14d2a1ba64d29d4b5132bf08cf46e96436dd73af5d06168e5dd3551f3facdc7658533e0cfb4fa38288db9e7c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfdf1808a1d1491e3c98388b61b38573c83bb6b557548642618c075cf141893b917bf33ccb2201353cf005037fc4eb4ced89b504474ac07ccb814f4a35aaa1e6aa78c8e84d62e553689627f6a019d85ce6c50be6ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h719ec3b3ba1b9ef096d19c56942921ab1dda4b439862a0e25f816393a865055abb128d2e20c5a7dee346cfdb0968d616e44c03945257553c2bc15aa5a28398630ed137f8b49c4f841e487c43d3c73f6fd0754ccb1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1516c4d1b981605e46c251c0f8ca6a3d06058b22f753038f702330a74588dde7cecd832f4246ae3d9853ea56990a7d94d51103f3f70c5b91153fa1d79c603a142575fe24dd758a3122c7a3b743420f1095be17c54;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4e9186297b12337608b28379d2fb7d4df619e7460561f14421c35cdd97dc6b458afbbe0185b1d6e1af76b2b4ba045cae604b778021ce3d6406ceadfa68b3b64d4534b6b0e7f45bf640ec7421b08d9efe91ffd62dc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h375e6672ef56681eb464b46bfa80dd7bcc3d6d23bd0e3bdfd3522f5ba8264bb40099cab253b1a9b9c8ca116fca7a0e056144b1ac2d502940eccf3c1e8435f3637e1a534a23d968cce1423e5fe516013480e593b3f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h80d0f141e56a076c09aa30c11291a66adec15f96a20b15dcc851f82091b6b88862711e79d71f06efc0e1a39d113aa74303c1093e448a748432cf873f435340b3cf64504b3fc217170a713400aba915d07f2e60360;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8fc5b1025cc697e447655f52b083ce6c36a003408b654702c73789b7450d4e922b1860e629d3c3d5a0ec682877cb53abe8574a85576c8d9e167f6c5d320c939a8a48faab4f19ceca6c0d9b45de44bf72e5aa92c9c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h911030506ff6c551dab7193f11a73ecd0d4e362ca6382f78f3c298557f71099f5453e74497037b19cd2ab108b6c543f4dd1f4372cbda561fed30e156293d40814f88ce9c3c449046f76200f8df38b2d5ec621ff0f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5048d5608f3de6521aa8c56d66b6fba41a3ee54d5d914f1074185edff767800a272f52b156c68eca3b7cd59780e744570c052d167a234f0e5e9e199cfca3e0ac3865c05e2b21a31b1b1f0cdbcca8232da427b05b0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36cb19f9d589ee62a3d82283fdd6fdf9d84375a04ab6f199364c5daac48f2fd5019938624a4ede5cb5b67f88bef17ed7edd8e0bb4bbf14de0a037adac7496f62e24f111f2d5a77ce1e3d291aab088fca23f777ad0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8d7f7caf968a747d64e238e491ee8c7f949c3621f2405d530bd61993afc6e7f002544aee5bdcfed43586caaab326c4722a4caa8c31f2f69174f60443f26e880c89b3bcacf0cc7dc569fddfe9fd3fc085bcd8e0fb6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5c06585de4fca14a0687ef3caa70cadf8823122f0717fef02dd65c530705ae469ff5481b90c54ba304e2f3316d72802bf975288f32cfa23b9dfdc79be059938a4f08c76608e35450780b667a4b63c997fe14ecb25;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5fe5d1ecb7ff02d205829ddb7b44d3c66be3b31fc34147656207a49a730dbead00a5899623c8b5fbcaa467ddd3b27f5a3c43772766d2ec23a9a8cea72b696c3e6abfff1d465662af39e25dcd17d945ae2236b73c2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6387127d041cca25ef705fc9999dd377ed2edc26698e3508e7ca6b33e27003185ae270194c7be1c53e88c43d9221410a50b13a8ebac294f1837ec569f4ec24e316bb02abf34daa6a61a9e6bbe102d027edaeb768f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7b137a0eff41db4d64f65362a409c27a63f84005b045e5b9dda7b5cb65b20a975bc5a5b88d58eba8882583e4c099dc63d4da3c254c7bfba498980a3696f382db950d2696cca72b65883f8126e436c43a294379a30;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b27612434236f4c9438fb0af7926ef750307465a5faa657bc1392baf49c6eb43488c076ed24f78a82bddc0efbf907fde0729b4d9adf485f3d170e12ce302a12905d04d7a58315206996e3126f258148eb568ffff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1bd6d80f1efaec7e839eececb8c9aadcd1e44893f41e5bbf341c238399dcf935f0950827405e81e0a95741dade70c4b4d0f43c598d7409ceb082c4d149a0e0d649db9257b0e78cdc034f29cd071d93182ce92fc5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3cd140b56b3c757818dc5a3afef96ec225fe59c99c7adf3f4a48428fd15a5a3753ab561e179c5fa65779b5e28d181fd1e7725f35edaa71f0c85cb5e9fcfebb87b8b333433cc23a08c0196c034b76069dcdaa88d3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h81eeeb0e7d0491f3896e08da7aaf5bd31aaefff57f7a511083aef13f72510844cf5a9df8071097f1e735df72b6d620f67537ec3851ccd64bf6369b6d2c6c45eb58b945eb4079b4ae03b5841cbca6d9403c582399;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8f8b6cf1498ceea93d09fb28c14b7f7bdba5066d889d79d3deaeb4b44146cabec5e72e709508f7caf4dba59dcab4ebf4c9637c4ba8ef2671644907dee0cbad09ab72da62e4019d6a48fc4601ea43c1a2e60ac90d6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6849f5c5bf9d82775b898eb446bb6842aa76ba4f8522ecd8b7ded27cbbc422ad545344bc6d41598516ff75d36280d475093cfd2cc0a1fe80e09e9e6e1bd54ebf80348a222a25b43ecc26f57c238e9ef24084da507;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hba5fac9e094b7e108202e5a1de327c872c8076b649c25bcbbe294970ca38c31f9431d225e52f71b5fb03a61112d2d0484d2738e453c6e49aa6c84f98865a80b975d7c9f1682b0b5d222a8878504c740e66b1c9ecb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h28cce2e5fb53bda2026868116298d49072ade203b17e67bed8e6a69f54803235d20b910a1cabb669eec76f58db02dc072b62d4e45f434525ec13a8c7132d5efc98cc460e543237252bee8b8d0b62d2bf71e58e0a5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22bc0aa933c27a9759b1554ce5f606fb64c26f997d4ea57579aa23adbbe54cffcc7e6490cdf39aeaa0d1c4e5f790db8b3ffe4c1a7572eeba0101d98884953e70986baa3da2cf68b6356296a9883105190f2f95dbf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haff7a801f5214c9a8ff1aee32f867b7bfa86ff43d26d98d2bb3fe9905e611c7f423ac482b716089241348479c802b59f08a49e46c208c17669a357363c7bd507e215794cdc42661924679d6cd48c475c3b46eb7a6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h341f752c5e30981370f72c6ba184d592198321ba64944cc0739352c087ffe31734c479ad22ae0be17283df0705fb2833d870220cf3fd3bce441ca84f6e1ae223dae4e748b1e7a4d80b72d8c954e3b3da93c584faf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha58cdbdb64eb615377c87079b0a859040f299b173b1f63403fe4033cd667ab1b6940d081487462071b115e9d6d84d22e93cc7f9592e7d4ff67364789f93f6d6ee67e7976c262a400b9696e6835c86fce8cc32369f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hacaba98172fef0f4d925631d1ce66efaddacbf7482f16a57977fae030b858a850ed481e19463b118a838a44bb8fba0b1a6d87d37c6d433e733287b341ce50eda4fa1bb2ec51218753d30b935f593ffe6216d87bf5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9d1b1762b065f03f611d514813351848c103df4012e4617561a02265c7e5bb439dee282b72e9ad82c95a2ef5cf8a829e4a287f83b2f87a6ddf0aae7f9619ac2c234a3d0bc1d86ac4b98688535293c2d8785df1213;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he3d8a2999a49a01e3c73ce40c5bc4f69d8647be2387b9a368453d93a2b184f121dc84899a480badf1890f0997f5ffeed2eb1d82e78211c64d1bdc421243ae3e6d5ec65f9b27ade8db65c4f960759e99c6478d96bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcb35ac8a9dee35bc88ddfcf5ee9186fd6c94cd6fea74a20e9f1ea9f92fa0d0d662a0f573462c417b5c0310b47b39ef15c51805944037bb9ebc0dddbd90296e10e37aa52a7fbbaceb0130236f2a07a6a0678c31643;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h932e989f04c898e7bdf2e4db5a435ace3f7daf855f3bd3650a43ddbef0681115447258d5a28fc7d0a2f46a6d16257897fe11ab8bc27c28139f986be042b95ab9ceec650eb9c2ae84172d5414ce5db74bb334381b8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd2d4c67d52cc7c8653aeb957cc0d095be60d1487f7410c00686610a13438db9e844e17a40b9a2516e26c2a922f5be6bab90822713bfda4340706fa1641e519cbeb0695ad6fd31935a727366b9b36d9a696762977d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbdecfa33d2de024f6dde72481f8f2000f843fd21c50f6d995275bb563d7ea535874904616c0f605f9bceb986b60006a2070f7e75a2a516306764e8b5a2ce95e251f4d60473530d92ec840dbba5db4711a0e779029;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha8098430ea7c2c9dc7321102872c0c9fba8d15ab158bcfebc165c5b0b09c8f8ae7529fdfddaab8622cd852c097d12216dc1f222e013ca942aed2516aeca1ce2aba60a6469d3eaee26f781b3a1db68db53efccded1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa20aa88be6a78da795bae3e9047fe3cfebd38ce06bf2c171e0ba6274f3d036868cd7f000460f27419a14f5d8335e9bd0321479f2708d3f30447e56bae945d1190e4e408f4921d28b980738d1c678524a5c705634;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6f67444c32734fc3941288a0865022bd27a6b196759e1134e93e2971826f7e4b69ed9178eaaa03c1ee161d69ed406aa4d27e3ef792d0d8f477737e082e41680047ce3c01c1eadcbf145ffd143140461ae841c3a3a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h53ae5e303002309243c442d8bda507a1ef303863499dd72a717d5e4b3bb6431651348ceca6512e353843e894c57dbb81fa7561e3d1977a1c7576a713cf3a16243891f94db5580aead0506985987ff794d403b39f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd175ec6ff4844a7cd9dddbab82d6c7233f5f02f30f7f1bb2b81c37c8b59607254bceb980ef6110c8297770a75d2806f50207b073fcbc6897ee50299229fcb24fd1409e859d312934aabbc725cb3e97e131a01d870;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h90f922c04df96a4510b182b237356daab1df683d09180f18c0bd04e0f17589b6dec751e6837d116408ac2679bb3c8913bfcfbe9cae0f6f55be636c565c40ee82540fa4dd47b9e18b4e850e2e7ba5c8f5d01f13c36;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf068bc0f7826ea25ac5b6b0b840bb62ffb04bfe1f95a2146593fe15b64a80669d45e8e0b2850e26c7749bd588ef16b586e6a5a00f65ea78da2c0910fc240b53739be65ca59edf8640115f2a37c28eeef9972a0101;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h268e9443f0e300070713f8f9362c939e2af389392f71fd38ea205027a9e24c29fef291722a6021afea1dabc9016c32a66ccafcb622b3f8622597682e67d7dfccf38ed9bc41187777a2c157acd1baedf7086b423e9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b6a58f7dfb00f4ea0386bdc94ffa270a05ff6039184019aae0a649fe09e188437c07541c0dcf8d8131f1daab8cb97ec122a746b1330e0ad11dc44e7e6123d370c084bd98a4f4a617552dd3cae0742a01539ae344;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h350f80d8fdb66fdcfad58b52806b47d22c03c20f0b0f8110001a9ebb92bd16e6ea358989b3d6d841635a40f16efbaf5f412b11ef17f91be06a55c1671565518c018b3e6d1466d3966ec0f3aca9f38e78f432fb1ed;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a5b2ca8a7d1fca16578da5e7fda1c3e542e262320117ce2ac3bf71310cd304a6fbdd5ee05b71f07b6069c790fbb4f0d086d5ae0aeab83ef6762ba0b86842e9d13ef3128a73b061bcba164bce0fa06d4bf377d94c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd80b62281fcf5210fbbc3e9482b33f2b4087a10f957e3da8820058bb08f2a3342b748b0a6fb2ce8eb6420d7075d15f7e1e26d2ffcce081a332a4def83d6127af95c4e0d1411e0175c4ce80948a359a6e7b9edd2f2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hbc2433e6fe4ba93120d56665bd5e24174e0326205899cdb776f277400373e770f0259d5c51454bc7fb965e1da11d321f434e19eb3f7985c847be3243fdc9d84a4e7531340abd2bf88f94463125980a4c4738c3333;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h252e75e38299ceec8349424cd192bbd663f170b30f07b4a61f178e8344b28e1ee0a40113ca07636bf5be74c98b4ff858c580e86e4f12ebe5e9bcbf84d21c059c8f549eec57bf1b701b785b0cef052f2585c0dccc0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h901b5e5dc656d8707ee2424d2bf317756f95560d6128989bac5cda521ce217e3ca9ce32fb6db6db5de88b6f588c7d4ac2ac0f76fac0a067a7be8ec6d8a3e48436e6657964c4c931c05a8df7136dd911cfdb647b74;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6aa2dc6dee6ad29533f9661f7c0813d09a57a45f54dfa74a2a96af6b490631e7c713c48d21cb5be31f4969cd9d5f28db4152b63196b628dbcd9ac554debbf27e8d0307a20563cd18a97b53182b85105242be6e9e8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf5f971a3f8e181d374fb92cb6b9280c8fead7b1b0e4f562d21c7722c965431fff619cb19403fdc6dd04ea82abfd278f088d6d601a952c7809339a0031016f7b8b3dbbc9e830b8a6f8a431c49364b9e1e6f89a5617;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf7c3f145604c128147ce6a2fb4ce172df7505ccf504624745dad11a05677d72a2a323a8faeecdf77ed7085457e815e96b62514d1759434e03ca7bf2590ce90e336bc0f35394128b81e8b1f14b8aeb6e44015efaf6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h91f42e037b690056c9a06b2e6c83aff7063c00a2411a5bbacf5e92074c58d11deefa2e97de23bb966e23f20d48bb688ce4e2e97abd38df46bd23607aa957a103f5746f909d6e6648d9b4fdf96787d12f4d849edca;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc1dbde5cd0e17e8f8e53884590f776be3212f256a5474de0381e3843dbc84e5c3354223b771132993e653de38d910fce0d92e00f86b0c9dd25a8cf18cbec5d03d142e3a23fc98744dce904de0acc424873319563f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hc6199dcde3260ad8f0c5c72be7e6c51dd0656c635ce64d58b5f79124c99e9dad28eecc913b5dfc3df268dfb07bc1c4da8609f4e0b64ef73af5e9238f94cbca85e1094c50573e63a743a15e3fed153b93e74c688b2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h69e9a611d5c4d432e078b09bb130db4e6d1b0a51e3a35adf23efa9d91b9b07938d5b0a0d213326625da940bf45b8deb0b55be96cf8b17f0307061c3bff3d76ca78473a18f807bf47b331e7cc1de217a5bac47aa28;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8cfa388764949dd9b273a0e9f097e6f6cff89099a01f78598d5656770da1ec0891beee7d42840830ebc4da6842a0bc6036897e2eca23ee97c2eb41f53e2e53048974d7a544404d4d0fa222f756c0fe3fdc78650d5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b60871ad31df4bf62e095ffa8a4b2c88c4a44d499c69a9c75c0bed2b7669aca6d567ec7659e2c46edc89f577063faf6fc7efbb64ff67fc33622d4bfd83a0438b1d0cf6bf516ba95e589964b1ac4b24b512139aad;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee8d21ae75e95214f7265e679c620fd29443e35a96cf08473c39c50b2a66b7e55090c1ae2aaa353673d733ff4371a30830e8d36538e1c2c59abf74e0754efb701855bea20abfbc5567dc99d829d541fcb344f9512;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8c2e97bc6454385a9e61990c0bc40b7a49a902f80deb2c44f7c6295ef419af8cb8c47258531a7919ad9419d6cd08fc8db5dff952c3e092d41c048636609a8464d8178fda6ed12023053c5c649f8cd158c37184deb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6a6154e43b1a9d902fd64af28017a7d368b3407bc2270da8f48aa71dc6d5b266e9413318af215c554dd846abacdafe43a6ebb205b508cfd728bf63a9efed4f97c42e8b3ab0eec2d0752c3e8999c87ce2951c36056;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h99d7476c3472ef9d69c173f96e6b726e13595ea6a96daf2a7507ca5ead8558591a11132883c1427f1b33bfa8498ed28c412d2d5cad1ba2c4288172ec5e353db6f44da3e9c6ef37f118bacd311d7963badc3cd1573;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h49e3b70df789fe5bd9879a59dad1545b9e9f421d5a23241e54a8ae9b539b1243cd59f97055b4f3c7af7cb30ce59f8991bc2e6ef9d073e1e0cb59d8b0e927b501cb4a9d158b0f7bd8b24a12ef5c6359c96a7e6a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hff0a3976360d8232f8692d0f965db1945ca06faeb3ee4d74e800eedfcb89386408e4e080ff252092ef5020dad8c86953db4056df6b5bb7e0be8bf1e2dd35bc9c506be27b8636077ae240432040ed5053418fe38f1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hae200fab6bd588de6fedff406e13fed549daad3c7aa0bb73b5c809c6e08b52d7b41bd93b1a1fe8c8896a5e85c89c3aab93e39824ca62d32fad68a12d1cce1c3a0e482324e0aa775fa43a08d00572cdc8900c9fc06;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h77f90f9a6795ca1d3bd4fdae7cb2920a2133cfb115c9f93d989b93cdca4be2612e5c94987c8f90fa5e4c8350eada67ce5e3cb2ccb2e78fd692f00c94e338978d70d92d64d6a15f1780c046cfaf6458526de6fa0e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h24e2a1acaff80778d2b8de4956285bcc92c07341cca0eefe15b8474d616c3093e26b3f5ec261b9eb215ff3a049b5bd2df6d2f9356b1816453ee8a7307206698496060d01958627483cc0d208edf193d06fd5b2dc7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h64c3892cd7f99a12f5fa41e5954946419a2fd084422520afb3e8cd07dab9ac9308b00f2355e820f4010691a99292b2c5e9d2e10abf3e0d2b68c607f778249819beb6118146441104a5217fb733f8817821d9cb17a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfcb68cd1e3d87a9f0547c3d511975fc377f8872bd25dd29822ffc3a6d18ba9b771cfebd377181f4a15055d20efed6a3512c0e866729c63f371b2301f9247d5419f1825c8381fc03a768dbbce54d900abb5b9fe1f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h705fa7d9b4b726321baddac1c2bc83d19bbb4493e29646a58843b08e98ad015e01745b651aa1d80d75c0b396e0612edbe0bfe39f5e1bb716be1e586a8a88cbcab0614354020c2492e558ffda144d4b4ca44fcca92;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5e6f1f55e250f3fd341d7a3754af29a5a174ddc8240f8a7de4ff4be406229f2ee4445d305f08ef686d8eee2a0c705a1a09f040f2327b778ee504a7313e80854cd0043b09a7d10833782a19b5ca575fcee82b07eec;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h36319f588e3f2453f7659ccf09fc3929d845112f970eb1ef7b35df7a18907169418969891a975f2c087c47d426b401c62d8f9d8a6ad0e18347612a9cf078ec182244031d17bfe3e38510ce1ac6e81721943a0e95d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h51bd302d06e21d5caea30f13573ec2c86f2c6548af3a0ac73a347c069f221db5ad6abe4377292144a042cfb71dbe409f65cb9ea00554035e647307a6b32c7f1e65e199d497bce4e9a7e4c3b58a797ddeb8e4605af;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h566d00bcc3c3dfef68016bc5c0df01f88486340158e4f3571ecf484dedf63e457fdeb2f0ff97959fa374b7d533fee70cd232f0585b9133050f62fa03bc29b167bd1abfb5920de562ddea5b7da6eb330880dfea72b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hada64afc86a1ed325b8c537deea00a508012b151794682b978923f03fffd0812d3b1537f414bcc9e0a95f15a590a39e604848cb8dc7cafa753d7baf865779215b8bcfbfa2fc7632d08eb46ef88306634e2149d1ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'heb0abc21324d42fd189af0357d46f7970718ed1cb4c5eadc469a4ec8290f09247e30d269d47f6194ba0e115b95e2f6e97698117b96255017a126681a0e9187ff98c054b81025d6c84c6890e22b60f5d062e55989;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he30f8caed2ecdebd4a0ee6a5959cfaa442d91d210a5385b444e0c91b5bc3eb6a3bc81f33f03ab832a931b799a8931d3d170fadcbfe80f904ffa917ac88666df508bd7934c698099feac69b7f151af12d8e66099a0;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'had5e55758a1a428cf1a923f2c3092a719edd953c664a658b0050be3eb7cd374267ca95c29942816c3b65a2cf476d7673dc475dc11821ff243999a7e4a24f1803fb9f8d2d8f35f2b245f6bb6281138a403aea4681;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h954cccdc1007f72f7580b70887b15b1fddd961b48f6032782cbb1781e4d7e48110b9e9f9dcbe4666e35d91ab0b6efb162dfd51b60d93e164af6aaf66d26b469d621fb1d9765ff3fcae0ac932dfb5d1fb835a0442c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h47e6ddb3d7eadb9c318402cb3f8f689eb9a6f02fb8e9d330bea077678d9254e6a2750079ca086a18d7e113c5d1c8d02ed00f56ea971f69fdefa3b42fb980f7934c6059136e06cf982afb73cf6905f3114678600cb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha0bc10ab060923110699473e796819ebe260af038b393e7654feee5b1e2224e81fc06cd691e3f5edc49d330239a2a514d558277cdde120f452601f7fb504a03404020d7dc30c704392365d24f04ae5bd1a1c6e71f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h553530a6ab340e17eee8f392adf9b730dfd6f384d1c68e47871aa1b579c8b0a5ba05df1ca52e22009945a0024ece03b4f8889d63f6582ac12c56042d980b2c56e986f83feffb85e27d3da4d04edc9ddc7bec0c2eb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hddaed1e58d36291bec5664c0d1c2d4e82ebec6fecff3689d962bc44ca0aded9e0e6892f905711caff08b09ef1a2f4b43270f6b3c03058cb52075852881f5ef81cafd15688888f0249b06bfc9d6141501547208ea9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf1359323c174ddf61a38375795213b4c03a6041ff8bda8651f2ea1bf1f3be123196dd2260fbe4fceb6bc891213bec65d1fd2b939d37cbb839f44235b19e006c1cf89a6da665e5617f8274f3823219d797752579;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2fbc67c3eb0857f6d27cbb137d057d001d5ea928f00cea45c2c4316d9eda97d8eae6a9bae383c860980ae845e21890d99b46fb47e70b4bb081e3b441586c255cef4a826c6a4ba949688482a780d6a1b8ce2a92f21;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfadc1934f26469e709bcd5e9ceabbbab2c64ca7795e94dcc9c405d36e369ada79d3516cd8c8ce9f482e09566f92db2c20e591a371ae2f0eaa0616b0b2879b2c4efe703103f451ad99bdcbf8b707c74e562b9b8c3a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf770ce4e062d28886db9286b95c4717dfeff663e31f67637153df9d04646f58ccb0bab6451522cebc744ec1f169b2e3cd254f7e7c15962ed88f403fc1a9e4b076cddaa9226bd1f8b8ad09eb8bc9d27a7061c97360;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h59dac546981324e11f6cd3890dda3d6ff55f920d98ba6b560d315512bc976fc2d0b816acf26077bff996d3e9b22c5d65ab8304e79adc826ddaa3c5b6e9f2039b392d412fa7f30d6822526515d20c7278766289144;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hda93e15777460fb9ac0024d21e604c07b7cc312cfbe1220c0d60f48fc7f345d52487313038cc5c64ecb9069527486031bde0e1567143bfcfc284d063b45c7a765567e5272b9c8f72037bce31cc3647a66b1304209;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcf15bc6b3fdcd8d840c96d19284b8172f9221d4dff86d6269f3c713d633d67c6231382242e9382d95f35b557bb0e3c6017c456f320562be5515cb28a4b85548cf11f37f2feeb7270643e666afbde3e0103168141f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h60de36779fa956f01d4f89a63fdcbcd77c03f74203135ce2bdcad0df92d19ac613d45fa7a1c22dc8916db16fc757f0b23f2e9fb277142fe173ec9111d408cf3adf63b14d837f3ff137a440e27c186e4668078848d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h93e473119a3d165494ae67a01b07869fd7825b549355e8a5e021335b7238dac6c6c3add6851112f7d013e4d812f42b6becc21de069bf4758768ff834f0dbb58ad74d544f4bcaa738f16c023ecb89e12ca10ab5907;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd7878b8e2551f695359a748a0fa4ab54c80f2540e45369f758228e20c684be772b3a312f543abeef50743eb0fde9caf781dc5a41c7fd93202482be4bf89515d61b44cf531febe43eab7d33982624f3a90c855350b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3f51066ab0caf4bda28ae1c7781b658a84c5c2466ff11784284bc52b770b8637d4677da9f3054dbf5f431547d08ee13f956b0c05cf655e827df5388a1b1f7d694fe0acaa5682a55c0d396ebf6258e9d4ca06de690;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha50a8bfcbf3be9990540520edaf7fdd63cbaa2c69ebdd40b7a3fa035c7d0598c7fa5d8ca60a9765f7f66edcb3030d8be740adbd6616cbae974e68923aa23de748713c80ba5f56b893aa3e06b035e990a846f1a222;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8367c870458be05d17d7540b99f90d6c8112682c2b900adf233e78f25ec41787763aaabe02b392e970a4019544ed4d3dec20bcf9f8fef9c91f62b638eaffa556e1c93b24b4f477d89e2aa6446c71d69a25a8a7269;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haf0eca64bdbf43e9cf489c87a5a78306162990d5991b2128f8f1816ac29fa5ac1fbe345eab1b712be23a81a1df20a94e6aaa1ca2177fb84a057eaf19775dcb66fd3395e9fd8aa1f4a3fb4bb5103081d6078de61ba;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5f8da335ca2176e5b9dfc1de7b47a61840301ddeb4667ff6c0315924b266c101f145bdb1f19e44de467261e06935b33dc8fefcbab1364046ade53ca42dc2a249dafe9a040b11f021e1ff64f4db5d27a19e1e60667;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd79542e1784a398ac5e456ad3e1835cd808add573843988ddf75bf7c9de456842332c5cdb01b33bf03a39fa7e45a839d661737a74c6f701533294a7318fffd1e11325b3d1d56224b3bcfbaf4c251550ba1da9f565;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h982ebe13c0428fdc4fd981993a180976a537fd9fe8d5975282f22452d77da093e078c8d6d3d0498a317de6028dfbe265a98130bdc24f4af8837a1a50091640e14b4d08f5a9f83128329f9b06d56412ee93300dcf2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h43639389cb7d41fbcba79fe35dce8f945ad10f5e970afc6a94c68d053c02122897cea61216e1106db885d3c1883c11bf975d23a9032efb9fd8e693c38bf301598c844cd26659f2e4d0b762703bc31896e0b0174bb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h71efb95f345d9bbe8b3cd60780f1b4f084d4d58d06bb84d4536837682fedff266e0b2fd6cdac7468f0319f0558eff1745dc7152e70e328acf0ce4af182d4a13c7afccb5b6d7036535d77ce9aa2d93b2d728f7b1bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hac714b75ea3bd16b6df83edf7878a6e08d0b1a3fd3422337bf14097e6f9d97e3e2193fc2cd2ce1dbffd5893db95fecdf8335ec342e86a382bb680e2694283eb08aa4ce78714236d45990230303e5d9eecf0f77020;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfd8d14b7c08111c08c637eae00de03a433cd1bbdd71f40b2a8fffb30ca44a97041c8d9767e1cc8f934cf1612bbe411c97f20d8af5a8456dfd15310a1640f3cf9b827d5db2232c0f57148d286c3a30e42a93785064;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd49d2ba50a4493c7daaa668b4b5aa04a80a5a269745f205ab11ccdf68eb3caeaa80b13ef545f18dadd2132fa6dc43a5016be77faaa2600b4e6b1e2923e5d98b53d742fe6b438069b9dd9dd13288519798cff0058;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h78c56c6f36b7088c0b2d4e1c51fd151dd0fa8bbd3235a09f5feeeb5938f983995ea4d1036f4d7c5e5dab4a793a66cc1e8c0ad77ce9ed3179d8463780003f7d383cfe924dfa08b65d1a7bddddfd41ce235f2e4df8b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h66260de0878d7fedef167559737d6707f84b5cd83fa0fccadc1c7c69e90a1023c43ce32f2a8a0e9ade74c240fde00a5279c62068e8157ba7d0f18d8d7caebf57cf8800b87f49affe27c06b038096921fee58145e2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h543f244bfe7b0d4e0e45fb3a03b14d615935c2ab11dfe82935270b815e0a4eb8ebba8556c8b10f4c730fd2389cb82e6e744dee5ef7846c0d815bb7d793ee71dfe6b68f7b34faf341d2f00a7fbe6db69edfef2d12f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6df99b0e5e08a3f9f2d45fa55628a34351d5a539dac4c8d4bd327ecb107adff47f5dc0d4102c82f6298d86278f78c23c4c2e74e127ed7dab056358a4cc8dc21f2652a4b6d04d76b6bd24d9fb35750e4297bc5eb0f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h92da925fbf31775b5b11c245bd02b6fac2cff3fceefb86767cb5d979fec2f3216c8c304b30f7b89f6a77aa062fe72bcf6b908c4505b8cf08f7d81dd7bc809238c43c0eab2358c0814c3e43acebd260ecaa8eaec7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9acb7066b08d7f282e34e3408defacfad0010b12856f07fceed897d544b428558abd7ae5d1d555783b0a5a828e3cf5224e7b468cec48a783248e5f05449a116805cd6ceb8600ad4753c65b66063f4d61fc3f8297;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he390a550602a4b0dce871b21263dcc945da33e43a6e11230a2a4f7ed459460f4bfb668e723b8a03b9c886454bf984a3bc9e3da866d4bb725eb4ccaf25960f5874ddea6a60213e635cd81f30aba14b646473586d70;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9dd2c78bdbd4dacf06f65ccdb0857e708a75a8411aa6df038886a36944a313fa8eb6daa6a61205c62dbec120c6662a10f4672b30524073920cf1fbd6e4ba993904f58c9c8a53272fd2e81651b334ebc5d83bb177e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd448a4038e984b5c555f5fe5dd1aa6dac0fe393ea3b668a8dd2bd82df66ea37118e9615ef349adc19be7c35097a98e1dffebd5e03358809d556293401efbc4b1304c3fe25435c2a9b203f5fb5349f6cb7edf59865;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h732c50fd38b0b127b47fd82729ff50825d3d5a28a89204749b5dc0542b34ab9989e68a4fac0bc943e86ba723e7d7f954678ce0f5a6eb86c26ae4c8c70e43a7d96190ef92e280ed95da72e8789dc9ae8e7062c17a2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he8e08965786605e381c290f69a3c0b4317ea16cf0128f2ff30be2cf646e1f42fe15493407a39b22a236af7aba061708593a3f6e38442ccf3b899b55662b939dc3688858b0c7205d92b983190c7edcacd775859edf;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2f2e1b51e55ced01df057f4ec71c0b5e36cbe5cd3818af92f769eb139d5118255cd0643eebf24fb9d5f9f7b9acc85a3de1c6d99c671e055c93db40b723b21916104dccf2b73003d00ad52901435a3064acab25c35;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he103d2231aa1a8c1e32d5e8b0da6d489ddfde9a8f66a45d6c242c77cd71cc41e5ee0f402efedb3e54e349d075725b4864684b4a3cd1f9e4a4631e1fa348a2e54c5504ece0a317ffffcff39bd09a9ca66d78b85bf6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf379d4662eca3f93ca5f79a8e3c18190e1d0635fb992e6715e013f0db666fe01000ab71659354cd58513eb6673b07bacb4a532c9e4be0fa66d5d29ab1be9b284afdf2854ee74c7fb2d929623d1c28ef27995e0341;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6d4b721e21e03560d2dd73c727ff1b70ca4ea93d98402a240d468bafe9be3eb07cc8ab2f1735d7e3c12da09c295225e72533e41ea2201cf014169f39b0851900a808f1e42261530a68bad8ce35938042527a88629;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb1c7ad562ce77a9166dc89aa06f3020b7dca1d254715da000d749513bb479cbec72e216c5f5c5d0e72d92afc2eb5f96afd2f18be3cfd90b68cdbe59b458c45b82d64c6fb552b5ba4baaa6218f2e7d9dc6442b594f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hee0b3a630923a87302ed6ad16950ede412b9bb382e3c025e2e3077bb84d1fc8fa9fad397519deb73d6d5418940a50d8745a9c3ba4d680effa3da84d8c727ffe2070e6fc10e7103ae9aefd05db8eaf66e9c45dda5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h68a0747ee4a29c4810fbc8f8aac05eeacb8e0a6ef05a1cbf99709b460bd75bc4daf347fa6533f3364be762b8a5a987952595664e92e539f63062771cbe8d1c07288254b2b045852673ccab316a712467a759d6f63;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6bc406cbd59064f6833198218c9abd4cf7dfdf081fc6b9cffb0b5eb7286cd6fac84e67c8b3510189d3ca04a9d04930f3eda430dec01af60b66bccd2653b8600cf2b77b99f193ff9d3ee75cb05750fb9132264b02f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h143b3aefdd34a320208611970e174e8f99424dc844c8ca6032e44be55433aae650b6c10751edc68b8955a07a5e09eb8d80aa60e856953e9a6b4a2b78d765977d497ac269118e7358cfb6dd00791d8690ed80bdffc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7859eb23bdc088883bc84be4b205b1d824e4f4babe4aea386a0bfdd07feec74be8d45ca4401ae677c09984b6db3215f05ec685fef520a0e590017cf06d9944bc9bdd850419522a5da5120bf8d4a1a2dc032942ccb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h1d854f7fa019fd40404f5bf64972ec0c78aaf99e30f106ccb4a5be6aec2ddca8dacc0414b95ccb62ed6dfc4bd56a30e952c798245fd99b35cde2f7a9cf9cba1f9dfb281dbaa7bf09b4d2563792968bb8c5bfd50f4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha1ee6d7f1226f487eb67374efaaec33eb508f08e4f24489558bf48a81c4cfaeda71abc1824f29f78fbb62c7b6ed7cf018b3e6d21b4f1e837a01ec8504eacc8fe0ee521bcfa00e1c546bb75da02be689227c79c04f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8e7957efd2f9a500df0013fc102137925d1bb3d81c1a3ecad00f4c2c5100f5380e81843e16a502f83dfe15cbaa6f61d4ccddc2a530390f169ed8f60c10fb6822df123bf74c665b026762e8d88ff98602be7cd5fe2;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h198806dbea4466673d6b39aeec93d0c889bd405e9887791047bc62e232d2a7c896884f6570476692b17d04c15553443fcd348cb22604e7d18ad4087f75cf42c8a6187af3696a4534b9a05d02d1f9863afc40d8f00;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd9aa7f2bce5f69e90d0ef428dd9d326fa9b36a4e0001ddf3b5a5327aaefda1df70374a6ccd1db629e540fc370ca28604fbda1817b6d30f94335a277ce83cd2d30aa0637056cc75919813e8b58960e77075ac5bf3e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hd5b873bb0b2ae881d8bbe80e3ee0bacca4d6cce30cb736f0ba886f75ac50719e0c599af84d0776c26cfc6c02aa03261da9ae1c29b4b35dc8f24fe26f6751ef51ac7cb471b597a7f3f7fac99d1893604c7dc05a441;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h7d02f8ab9e4407cb6c63221126fa38c85694c9a3fd814be06b548261151593364179da021b369c5503d5b4c76fa81751dbc819b77d7bdf8e94ff1ebc367d17913f169d3ce4d4d27d7424ee3ac2c3bcd3b33a1a21;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5b401ecbec8508e877576dcfc742e13e5987eca7109b2d839de81b46a15df612ed4163de0ca2261552297bf1754aaf925b3fed6373212a48d0ea151a852713d8ca8edbc2ae1ebdf74a668a8acf0b7aed7cc370715;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8245245da6a811aa92d036219127fbe48d719339cc24c182566c75c6bf12f92c98e0291e43135d80303638a2661e34249652ec7b55a2f94d11ebc5c1e9fee7e46850cf013952fd4b5cafc5a9149b8ba8282895023;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4c918ff36fc31a7ae94a860d13abb0eea621124ad51959ad1be008eb9036a21dde19a0d6c524f4e2421f7b1a74a4555bf5c4218635f9d2532f1b9201bd72da6e56c29adb5129f0650079128fb6ddf82209dd0118c;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hca8ab78a3ace1a9be7c7d496daaf472b332e6be63211fdc1a2cf6a7940d32cde03e2d70538d579470280464a29c94deee932ef6f44b87a829025cc2f6c3affbd2618dce2599dec663117c1b51c1df84e8de5a13fc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2810fd1d8b6f53c56269d31fc76db83b41156abf67dea5448a7bd7cd7e34b0f26b15fa9fb12c6e6a126e967640985265e556d1b77aca28ae90d7620a28162973211c531e6e0a7f6ec38ac3f7206db7480d4ecc355;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h995f20e8a43ab5288d4e77d06d902727361833eb8ba53e7123799f6da88a13d4e7360bf347f463ccac5c63cdcfe9ff738c1c743d4e2fd25b98040bb5a6b129be1c38bf0e379794ada4c3571b9fc3f858821c8bcf5;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h8296939855a1c8972298e071258f2ce14aab290676c582160727811b9d597f3e7b6e6df777421d77102f37d7c0d565e2fcb9c66356dcd8bf91ed0358936e230ec625cb20590905bdc8006cc8d0b419547cfe66fd4;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h63463b436bb5b54723e1eaf1bae9624b2d1540675b4a15b5a70da4e53f5b6080b4b60ba1e239eb5eaad32bf4a435ea88475c91187ba89571264bfe5b16dcef234da634d95e436be76ee0730e4cbc6a5e98a5870e7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h48aabb524042d5e38d49cbce577e787355c6d6643977d6656d46f40fd1debaf0f0f4b8e2f7618ccaaf0f181afe9e0001add0f8875e3ca3b3a75332d3ae1fc19715981897ab97b55800b953127bc734bd8ea5ee264;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcd78d7de02127ae0e1255d43f94b68361149675eef58fbd13937e4f444baad24ddfbeba86e1feeb4bce84335d488de188776b73bef56b6d45dce21b37baf058b2889bb3d9404813c5b850f1f488520e620fc8c096;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b49a8074fae58b46f8a9e9428bdb9605e0820f6b7942d045a0d8567d83e06e0838990cadc961fe2197452c2ec1e9774ace2f996213abf1f59e3c6b108afaadef55318cd9466ae63eb299bc2aefee657ca2686031;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2a977f5d715ca904c7883edff20f87da487534e32e6e06627c0ae4651f1580fa6d7fc3d41ca0ad7d4cb4a49e3ae193de056220311e7198a3fe76e9ea5a3c7beb5dd637371041e43eaaad99b842b28d24f3e7f3ad7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb58c3101615eedaf514d32b4d64468fa76a739aede46fc627efe7c7c7378de5ae464a2ef4bdd33bbbaa52d1b2c26f0bb5bff765ee8a79e5e8a144859588e7651da50d6433a82991e82ac41ed9acdacc5f688f62bc;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5bc814360941ad7a3d164916c735c16f81ac49e55ea4f23d1f19a1d1138a19fb6808723f75036d8a41132d64c097052c0afea5ec5a8146019640dfe2958d0bcdf993a2a9b992ba6e60e1b3e6e23d5bb02adc95029;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4a843c920a7e40bef9b7cb6c0da80c63d78f09a3e8d2a4a615d031cbed03bda243e99782f4ce79e06f670845188d2a0784b38d865a54bf00b278616a1cf66b73a31d96329ac0f4b810fa7b6e1aa01b27998fe35eb;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h22248cf9bc2a8fe61113cbd6c83611e379ee9aeff0867c554c483058e92efb5348a80694d3b7736aadd5dcd1b549880f0f2c4e96cf416e5eba2fae7672bb1f7d2c8a28ef499e8cf82e662b795d2fe5492db98c16e;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h4ac8b9bf582f9bce01c7df0d2d59a0a3e4e6c525ee0601b2b2023eeafa5f95ae3133fe8c9de650c848909bbd1d648cd397496f74ee832a41d8a162dc203c86b1f3b124d82625bf3da47dfe5311ebc2b844868b953;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he1bdf2494de90c5885f70dbc3fbd94ea5b60dd59bc341e9e73e94c533ae3315df97f49750b0a326dfb81ff0efec8833b924225137cd10c57775557b288d268c6bc3cf0fbe192e4ac2726fa7aa73dcf16b94dad02d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha6030096ed8677b4f3c32d08b9a0adf023bbb3d597ad10196f8a360e35c6fb2a2769f6f65f19ad550a3d24faa26b16d3d07fe9994df0fead327f6c58500aa2b907bb581e20801d130761e76931ba9915a3929789b;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h2b82fa35a29e696cf3e1948454a64df5133e2f613511b50aaac3371681f314f5f855f166e201172e1e5df3e9ea278cea780160e53a2de1f8f948aa53b0e0255f40a005fdc2d6cf0e51aeee4c44607c60a211067ff;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hdeb2da82fde2e1cab5141adb49472b88a097f6605482f42ef6d219e571a47fc9e31775a2d50c00decb5b626835bbb6215bf9e95da0ffbf66fa44c73e7a34f1d202bad750f648c376ec9ab0573111ab997a958f7fa;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcc512d7d249f9cbb0d11fc60e9ae6ce2274aa15eb8aba4064293687225b1b85636e23191b20857fd41218ac239213d6f2941a651a01f86cb4387efe4bda764f39e017654ebe0c90dce584a9f6b5666ea33a3248c3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h52a15d49f5e6ff838994d067def6556570f94c4ce6a7e2a1a8e2fb9506bead59dc9f9dc5ef6310aa35175b79f7cba4cec423416bf2bad94271d7e1b41fb70e118d134f2552f7ef4100f5c19f839584bfb2908b8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hcca97fa22f7b468abc48fa76682daa11e768b427c80988adb72a0ca2f2a9bf2f6d65ae37987e02dea4fc14feaeb13947e998244480671ef0b5813b4408cfedf25e8a73f28e3ac1d034e28e31927a2329cf6e09e60;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h94f37440d5599993f5f76ecf97dff29a0e29e81291a0cf08ef46046e47d689ba9e198788aba4784e36ff8d61569da63fea23acea9459009846daa4f8d398cd776882a15d952d586c9c04a08c3e75dc270df03d888;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa2e0c48f34d3b61ff1a5fc69dbff6e0dcdc0de0b9b8f217d04727a2dbdd4443cb77eb6e766d92e104a1741bcb81e9233b2ffc289f754f1dcf1b43d24cff518df2ad7ac219d3adae0168a50553eea8a3fd7b8395d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h85881e26905b3dc0b67c456f6eeca49252eaf0da5da812c8fd9d60a0172a61502681030e1876360497328db1549ed946a464633e37e9bacabeeb4e35334042e9115513cc2030ba372504ade3974c675d9f94ff9f9;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf1387d591d5c45e569e18dc3bc54a068da5068fa91e8ce9cb476e9859d4664d82008fd1444e06164f49e6d35fa6e653dee9cffa32ecac008dce389b56b227b2bf88dab09a2b9d3607e12a2fbfb756c2ddbe4e1050;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hf711ee6272b73205326e93f71394e5975a8a311f61e5e3692f115362d5d4f79de3345518e323fb23f3727b63b4e2fb675530b2aeaff2949ce5f95ef6d1ff972f748cca61b369a08108effc9c57e861f1f6486374;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hfa704bd58fb0ef5bacd1749bd8c783a877ffb85280ead3c338b6f562f373da246091c3eb6d79ee943a090776c19792b6769b6443f22ff05104a59e7dd8beb3a1b3d278c1cb61cf45e577d5220a120d633c2196cb1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'ha37a44c7c850241fc4fc25a4053244a565b412f8beda66d83b5c8acdef662b6389d19839ce8eb8b88fe4287b6fff9f08d0b7b822eb47a5d4742e1f1caff3e7823fbaad12e4f247efbf3cf0e1257de89edf54fa31a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h5a0c941a661c19116a008874040a15c8a6cb5691160f6e9acffe94d10ab524446983e5bc01b5655323fe26ca374bd59395e2f9084cc1315c5de0c1a310e3b1dc9ab544a52f65ff785c8c868c37fbd76aca110d9a1;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h96d6e1069b8ec0f68df9460ed54d22549600d33cb50e3b1c6dc7394e9e7fc60eed039f379f0630db9b35d6b8a54406a7ab581ec070b085b25891635e355c90d6c9f743c0d6f2c767551a38b0bba85ac57ba8a0ea8;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h19aac42221ddce125aca36271d2f54ab36aef3fede624586a176d9c18e9d951b11d15dc47d628f9e968a071a57cd7b90e8b8e27c8628b1d11a177d5d9f374ad66ef7a61ee47b1eb570e6ea145990f43cb8a4581fe;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h70224714b9856ad14b671ffc35d77a3a1351d374f39ce936006f4d7f9b1b3bde396cedf8d65cc67b88b912e60a37d371e74e0ab2bc8215746826db4606149075922cdf98b4ff63631c2cb9cd0c49305db64fbfb1f;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h82c4b2679735e11de35e531d33c5c6becd1ce205a829796661a4c4b7f7177b7c4f2ab7cf601e17fef68b5e1638121998e952eeaf3906789be6e8dba071a90116f212fc0f954a410bd45357b514d181540c0268cd3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h55bcc5383944c17ce1c0b813487173cce6722aa9f5652870a483dcdc7a5acf57e8b4ea74d476244818e7df55fd5bd5e07741326067e8517a576d240758649c69439c5e70bcde27c3acf2f3ad910aca923e353fa43;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h413d2c4b98d8d3d6f3bf90e9e639c6995a58ab1407df906e9236b3cb2f5037b19ca608a07863c165deea23e8747fb1601a9db71bdf6e596e64e87b9cb06c6358d0ed4648f2436aefc8ec23af08e0c1e6a6b785743;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3b0c4de087fbc18c9248f48aa96d49d7956aba8cb121e112b1f777cc0e3ffffeeb5ef90f5aea9150037662b14823604f1f8f489a619600b4ea2a58f6668990e3903deb6d7b6aae9a807ddd848359ba42939f00f55;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h39791f16ba82e50cbf251e0c4fc639c803958d388d85b8a6179eb6838d3ef5a0791478e1092adeb777667157c474f4394dc6baf564006fddccef3df10228e2d5d87aee411cd2b3ec52d6d525be597524b646213e6;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6146f1cd397b121c4fa1846249cc56c4f3e1a19c11048cabe9e15855ed3cc5332ba6fb4d8e8739ffbab37d1b2e14b06efbb181e0890d693e539e8278e2f932d7247b7632892d6cbc4cb0ee50980412a2626b2461d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h3e7e0a6eca5632c069c33d560e85c4c73607bcbd874acc3b429ba439ce969866e0f1e2e934d50a165bbed31f87c7ec68aee22a8795bca4587c578517cfd35c451fa047bca9c36050b97eb08a810a505daf6410bee;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'hb8831023362802fc7f572601d2c000a5be5555703cfaf79e92956405a7c02099555165d8c581e1bf343bfd43b72bc2470ee892728efe12ebfcc6ef66a7735e8b3638c1aff851d70ac8dc82b78aaf273b6ac7da6a3;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'he9652c2e4690424f4e4c44ed6790dd0674fcbe19ff4b1e6f19734e3c193c105bae537435b3c2b0c5b3790d77d71083260987a4a7e065ea69a34174c25d511b0b9ca6a706ed5660b1fa57963902cb82ec630112885;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h9703d706e1be48a7cfbce06b085ffda78e8d7fc5f4f9734b4ced140e462389007f7c693689fa63b85fdfa461e2a6521360086c635c0e4307daa9ecad4a8ac19d41f80c9a8907a8366c0735d9bc16ee7e9b926839d;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h6ebb8a92dfa89b40882599e38b6227425acb74e230f73d8fa0e6f82932446e6a3a0e8adefd2b70c5e937dac95804cc0c2282cbbb4f9c8545184df5b75afa0f74cf07479d839c75e319f2159f1a5759b26eeb138c7;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h695ce82591b5c4fa56e49b9ed2521380da59a2404d7ac11cf092212df3623a3337c6d96a4ef26c9b93f932c85597d35478c6a9de397c63f97e395cf800c700449c36eef065556d092b220c7276e35c4b19cedd22;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'haa76b84e387c729670ad168761e2bd0041766474d275a5ca2b2e80cb1cc1d59c0c4e546ed0a40de54309a58c45d4952c18dc6ec5d905000acca28606a4ac93aaa4322dabf9c2f758e6c0083fda6cd24cf8a4b884a;
        #1
        {src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 676'h146ec4d1d4b721ee6f48cb27fd4703f6485018fd1b1b12c99f6dfe53700103b71e6bc724f18ddc00ed32865474ba0e084feaf9c75b9da9626f5be2ed7e9bf8cffe74df172570bb37a2ad8d782582851fc0f001d1f;
        #1
        $finish();
    end
endmodule
