module testbench();
    reg [30:0] src0;
    reg [30:0] src1;
    reg [30:0] src2;
    reg [30:0] src3;
    reg [30:0] src4;
    reg [30:0] src5;
    reg [30:0] src6;
    reg [30:0] src7;
    reg [30:0] src8;
    reg [30:0] src9;
    reg [30:0] src10;
    reg [30:0] src11;
    reg [30:0] src12;
    reg [30:0] src13;
    reg [30:0] src14;
    reg [30:0] src15;
    reg [30:0] src16;
    reg [30:0] src17;
    reg [30:0] src18;
    reg [30:0] src19;
    reg [30:0] src20;
    reg [30:0] src21;
    reg [30:0] src22;
    reg [30:0] src23;
    reg [30:0] src24;
    reg [30:0] src25;
    reg [30:0] src26;
    reg [30:0] src27;
    reg [30:0] src28;
    reg [30:0] src29;
    reg [30:0] src30;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [35:0] srcsum;
    wire [35:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7d45e2a480283278c0ed19c0131f6462dc1178ffb61c56481b30ac51fe66c7df5a0516174f7a7f8a742ae0995bd583c861f595bd92d80b14bf63ecb8ccf096bc57e5a06400d4080d9f4f975f32cbc0013fc26321998052dad19b79a187d409d8c5f032ba0b5eed742d918f338e43576dfc839483a3f05535;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he66bd41fc3addc8d1fd82f15fc7fc617d32e8824543b2870cdd07e2151760ef83f2d3d9f6522946a312d56eab589d929f8ec898386bd3065e58ad5248bcde391182be3247c1462e47d882b66b23c80e218d5b93ee8174547c3eecd3114620e235656306276596dcd9735fd794cddc2fd4b3c54bb7ef6385d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c1d111b3cdbad5a21ccc5acb5ef9723bb566e56965215a432a24148c4f26c1f213b5c2e023ee51f1687b5372a6701419f23bfab8752420f56481488738f09fb2d0d164961d6e1db3f820d526629d6107cd43c9ecf4a8af17e56b6f956ba2cb60e48268d20f26459555927db92e47cad3c90122cd0aab3907;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd612b9a44c73247d99611b575248eed83bf197c789524f31d7fb84b77f80a2d4ce8583dc771b0304cc4d3b12fedce2d17c343d0c044d2acb4e7a6923969c2dd27959f5899fb7913c39e0bdd0b6b6f143d6ff9656c880d94f879959053b1b0bf4ce3bd8b342115e477d112e1af7c0ef91df5e0666cca6319b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h305e01d112c337641cf079b99b533954ab8399a383846b8e49de08a5ace640e0357770e8fe9f4f6bda2ebd9688307169fdb204a1ba635846e02651bb358606d0379ea4f97134581370c8b6e79752f199bb635b7ea9ec15ed11bffcc4b0b702a8240e62c54194e37f9ffe5baa16ffe000c403d7621455b2ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1580edc8d6cae3a44cde033020e99b93d09c20ec105cbb6034b0cea726d6f29e5a500741bee080fc93daeff06e66d06323b3d3aba96618bc7470f14b39a48f1833569488f9742ac17b48cde1f60d56ca8d6a74f071b3560f17af921882177bfe6eb091166f13a5b64f6de8a8d5cf9adebaa9947e2d97b1b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc42738619ab71da93b2f99843faea2a945cb90966e68ba5de512fbf7735ef30dd3e2cc1f5dd5dab44fb6f1bd4d7147f67a2b9b39350d996facc878cee39c5537dd5256bc36d92e2614f907c2717a5b5a1a87fdac900098651e82e358a56d1c691b2ec9d7a1055f7cee38b11297888916e2852c7de0062987;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d5becc107ff31914a2d455bd1df3b2093a67ca0ea6a2461783d1494dea4c40f24e67acf1bb6ac391b839827819c99841c81dc419f5db389d46b4355a645fc599dac59e19b8f3e03708648f2e18783b36a30c40498315f8b893051b25b2bbf36e06c9d3febe0845db7e3a1e179ac76692f4d515fd77b429d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h75a16b4cfbf2a4bb29878e2fe9f8ed3957103d3429b916f2124aaabc18226abb4cc182006e38fa6eb15dc823b8ee20e7b7cc016d608b558ee49c9c8ad8a57e1cccd0353f6a7a553787da331d94e7db856e9f34ed9a014b10b05971e75f40ad9cc8e15a01d5e468c7bee822922158dcdaa4155c092e5edf98;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44817e1927992c35cccae7ff81f944c9aae5a69515f73d0969ad3d668d87b406331f225662561198b52488c242d6ca1e644b676654058e9d6a81fa8ca47a7de0c0f3af4b1b3b4dff26f57d13abc2f69c0f66d56e9eec89c4ff6a40f6f45567fa527b92e5685a828200028877c6cc55eaffef5db6308a10d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17459a51a5f99c61da5cee61e4c54a9091f83e13b8129e28de98128efc729d49c8c9d28768a6777d06f9db6b10a089a163211563d632b31e7dffe72e6d71c623c6c8f43eabb1d43d26ab3f137c2a8280764909f36da87d68e916c55b77ab8a0dafeab82feefb634d59208aba8f9aebe71b3cb0880a86eb47e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e6afba980ec04ec89825e4ad866169f2ffcafbb6b1d6dd3458dd1be5ed260800bca8480becb0b3a2a0e4deec1d791117641abcf83696cc81fa22543e121e752cf17ecf22588326b46e29b9a9e675a15ac38fb7d3cd0284354a8db82729a88cce14eb0065f77308e45ba0ca2203dea7aa4bacee27b2dfa12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc02381f9d50ddea4cdb6ec5b48238f4c12ffbc5c9b6b79272f04af7cb8131b670d1b138c3c2203dfa45cca95f1adf0e0b5b2da57ee5fe85aed595458aee58f64acf032295a6ccfc7080c1147ee20b4fe7e07ba56986b60329f6c5bb8e40de5cc0d6b5002fb200bb9cafc23fa6e6cae37c8224acf08398e23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ca41dab436cc6f8368db1b70081bbb6c74af108cfb39d908d4558217274192330ca57134dfa62b32c3208a25f478636c5766327f858c096faa5bcffc92efc9f929d2e2f8c4e272d30fcb5db62306b70744d7c585a383fcce33934781a6e884ade3b2ad699a69c2d1de781287dca592ac98490053b4c385;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h358a894cabd5b3c6ba75d2463ca3460a97b1f599a2e84a7ebf47db9fb5270f3f25eaed5836c91923dee0635f427a45235f5710ee3688083fd40f6ec93e73bdb09e5c864a00edc3254e881b2fee9f6b225c0e211e1fdbc6061ad9191fb875fd4ef4f878047c305d1592ee23b5599e333b6abe8f94a6288e2c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1420ec034bf4425a137ff6bd4614f31ee540d8c475dd89c0d7e7fe4dcfc1440fb6cab2e17c97237054d47b83fa865733caaca3b6b1db934eda2c42d7a32f2d167ce9b01e5be8c16dd223829ff65dcc1ef95ba59a22fcebcd07246d114d71ec0376ea951a2d095f0ee331f70602250f2d0459bc4ad8c74e217;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h125a1859f7302f202a64e4e07113875dbd175983763aa9d11079012565bab093d4913a90948705832d72fee0f2ea2145c1e29be48eae407c332e4dcad79884d3247cdc4ce754d9735b738218c06f0b0ac3cc8a5dc29e1ca64fb8e800d37a5a0758ca64ec236a867b1c3532b4975757f82333532611667aef8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35e5ef34523fb4f5459458195aba911fcfdee7f578d4e3daa4aea61fb2d146081bf991bc524f608abc18f73f71c6d7d39bff192569677f06f85ed033622af3e36e4fc42896dd91cf0c771f777a110217f8744ead661e11f5ceea2267aecad851e584ab5e28bfcaa756d19352161f6070f9de2123f59ebbd1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c2684ba0993e561b2a22b156dd4137bd47f9b2f69e90c5a952467ca94ecca64993ae88659bb38083a1916bdaacdb575aa038dc89f8cfbf6b3b1ca43ba328e15139643b09a8eb3b6027424ef46ede172af954a4bbd38f65af465e15518851142746af6b5bb336473beba6361fabca8c635e6fb306f991bfe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c43ad348c64adad3263b823038c9c92560809460e54546f62ea14764204f95fed12c5041fdd4bf2b36d26982ad4cffe16543a69d50a8a8b1e8b6588bfa237ebc27a33cdab52d8a97f8902bdaccaf0694a01762a836b624371814bc0f422106de5cb9f0fd2cf3d4773def68e0a4a3302967efbeae08c9bf7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9326db1a35afad886b85585addad4a3dbd2802e6fc97b455cbb6ed0ea9aa5d41582928e14fcf33b8d593058813a1fc2023ff91946ebb4ec0fab41d2ff7d935c83d22b946bedc7075fe0e9a729a377b2b1be039f487ccf3e71fc877e531b7b1a5a9031f58e0cbcfa853b1322cb5088d64645710336419129e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd6e2db9734580d62d996a375121b4bdb29a59e3116d3540093af6f8372be0bd83890718d25561e00591e1a6708be1c4a4fc095fd2e83a2ad6aa8b4d030350f15bbc860ba8c1191bcc8117e88f649a42c2a345c448b3760be94e3fd1bfa2491faab849f27ebc6868e41eff94d743af4ecca95df89a07d6dbf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1821d30138b1c3b759192fcedce86cf79853fd2170bc534281cb2da32db21c3d6e8e6c78107f27c6ef5ad1e03c9628d10b669cea65cb3827b402887c0067dbc08b047f70736963098e4319c10276f96b02c437bc6e759b055f128b6efcf81c67af46a0af5c98e4baa8b55aa894250e8bb14dca6e6e39e38f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e699554aeb514aa38a9adeb429abd5168671151599f5bd75eb27cfdb0dbef3c39e243701180cc7b82beb70c8b85e687f098c287fe175e8dbf496b4c69a18280f34b0216141297c444a23efd14839a04718077f389c65632d94a7808ef54467a737efe2eca39621f26dc15d17fbfc933d3177fd6ec3eef2d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0be42285c142b7c52fd7f6aa13c223f3cf21b86d23b511c4643617cd3b27a6fff15a9f8059d9ed56ac948519b3b02dd30286e7a2c470a5aab0a267409c4ad497751f466fdce187ed36543a2d77aedfe9adfa1d96ff5813c697f275a6a04d7d8daa3990f8b7dc6f10a73ba307cfd871df81b67dfe4357486;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37b690481e2c6d2abd0dd4697626df63b09a8079bffc9abffb1622222357760f97dbfc9f7fbfd41716c6f32c84ed5efbd0d1097cad7663647a58ffb47c7c46964cc57c7446c3cd701bcc1db23a0816b9be421d48e8585c6fd15c112f757695dd037206f8333519f2e97d829b2b2ef2133f37fc5e28634d89;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14e0a26fae7dc27a10c9d85488946b5b235f62fbc94a789e91817130cc1876423220ef6d8693e6cac845d305048d28d22a8e4f7456f986472f510f9c4243e653ff3197cf26e371968bff45e298f3ba1fac19d3acbbe657d37dc05bacd904d720d0ff6d4226801a4e356669b1af5cb1e74712ed8d10c496bb2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h21d85462f2ede57d3a7a6bddf33037a6b557338a80605d9b3382d1461917bdcf081b71dde7ce61bcd8168876468284f73b542a6ff53fb1d72164aafdc0327105f8e4dd8a5a0554e3b66a68e6055b8b95b9e7a1b8b6a2dcae30e15a646bd363394d2f9cbf91bf061f6b76ff14ad81caf53bfb9e7b6f4aff52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd4234e84386983c879d15c6ee565b031c33818dd822946796db256cc635c16122c58712f67723b55a3b2d8a7ebde3d8d67fed90368fd08bd12a07ee4ddfd988280285a6db5c22ab5825d77da9f28ea72512f1e90e499a7246176ebd1399c9e97f2ac942e3b2301ca2009aefd797422f4dd5c021b8643430;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17a53e15c29516ec08319bcd2e743e949cef768b50d7abe16a0f3f4bdc90cea69afc7a937e98aedc4ec242395927f226d0f182326f717bcdc92fbc9bc95a91f42049d7e194a8ffdc0d9356881dbb0493cd227bae05f379305c66feb51967bdee40e1a35567d1f86b9fe346be404d29dd9fcbec17122675ff0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b518703d83b3bb373d114a036620c71054d2549586c7c0e1d0f243c2b7e44aa8e3d39797c3e4d6fd4ca15329df61d30b28c83ac3acfd457b7b76a20f948c57b8d88ad14e1feb8b807b458af8d672f0f04d7b204847f3a7a07e6b9f12b105b710d5c8f4931453ceb2db806c55329d57ad75c1341c8ba2a885;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h123f41c3d784b5a1cf487b604247a570b24961a83662922dea49832e8b3658ee1bc5635eb3f9a0e761c7c46f96cecb302da90ef64189cd39adb9b1bbac6e854a95f97a40b36f722a5621220dd794089d67b6fe73f3550ace67ddd0800523c0d4bffd75b22acc9cc0949342301921688ff86e0700e53a1b8b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f68d3c8673c9e81536aefd42061da5b10c924a820c68774956461e5b85b8fc51312976f5f05005efb91673741b5dae3f382d8a360ef53090514bab14cfd38e45928651e70d2ce97385649afef28b3a7f9c44ea74d2ea0c8a46d949907d202436f2a3b182e2bdb435b1f119a8064a32167bcd9ce124f1b0ec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d099b561c530ef547bdc34fb457bae8148d511cc7c75189c924260ffcfa33531a537e6b7083c54a4af80ca8ed796b59d5450908d8979598579a64fd8aea7eaaa762ce0d03dc0d0bc505643b50002037996f33813070aedd570a72f9b98e50eb68d47a2bbd59f33969ae3292fb10b4b18fb4e0aa88dd313eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha322472b4d85412236264c98089434347717ac2d5485d8631a2d3b3cf60a88456e787110b2a1c269ea35af6258229a0abc479a40303a13dd7818918f594aa23d3c4a7cbb721efa302fa47a363c652535dcf2ee6b04ff5274c27049940ea523238bb372b5cd35ca69a186525e34b8ec81e22f23fda7f062f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58d0f704ac1fe1a6e32a7cb70bdcd2c59bfbd60f64e94fa9ca06649a0b931e8bb9bb6b743c1eecaea69b9b25de80aac1d14b96165c4b277e20d58a37b26b366b91b9b7e343fc8ae5c99a1e27feeedb203cd8b7ccc2458fd5859180da1d781447bc49d9c3c82d31eb07c2a03e0de9ce21dade10fd20d84241;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h53a21c03a7b8dadb2038e700a437a500eb34f49f32c50fed363b780128a9744a1786523bbb943cc309ba40e03820817a7271bd9be519e32a161419e74b12c04857bca7dd436b956eefa1fdbda5ea626239b31650e91c99165f383aa33711f198b9f7fc94743c367127d12274be8517b4f5588733f73d3941;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1feb93424dccf32a665c19ad558a53dd20f76918e3382ae661b173a2b6829fca674092affb7d6d3a403549313568b5a3cd0a4b8552ee0ba778f0b34cbf1f44cc81fee548b94da04a75206c13644a9242b5e451150b0d803e376e9d12d68c2ae8160fc7919b1e6b7ebf0306093cc37b1e1cfe918c5fae6f18a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82dda2f87103427b2061dcce05e8229f6d2cbffd76230087a93e0f5121c7d40d73893afd7649f0f82e31f5306d11b99195a7d91190da1bf0923a06b8d64bf1c22f730afa3b779e1d1314225cde5ad11402889ff3879939725fb6de6f27dda7e22fabbca9e58dd8b495a1219224f6f5411bc1dccb49a668ce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbd7da9c66111d7712b8802ff011ec595cf67e677c91a0e485c7ec65921e3662dfe7e86427754dbeb7508c92e7d143a2ad516d4bac2a63f400d17e06100208c15015033ee068eb6254af65c957849b59e61ba2ccf7f0a59e5c0d5a5994e0f7999a3267fd7bbc5f30e17b9cce262f01b4e83b2499deb033f0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9e12bd590608deb19e0199bd3a4c6c6be55e8cf21cde0d2596b8df1c4b256fdae74dbfccd5c6aa0360cc761be581ce0ae128b5d884fed8eedce4293853a8ddb3305a2995e46e8567659642cb15e99e9977ad8279fe45660e916a481d33a203ecb073d8c9251968a8c000c1854d97be93ccc869cd6d27fb5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3eacbe847c0f191ed4a2657df1831cebc5357f7db2bc88fe21543836a2a28e3b7d243bd469c67debb33ce53fb23dde60f5eb31763c93003cb8cd65f057259926f6171a362c52f270e7d21163e8cc2008d0393b1ebfce2dd5ffd2d23f9c0c886e9fcadc64fb4b21fcff8c7c3907bab33dcd3eb4fe18b35ebf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9a46a2671de45c622cb04c4b7515f8a46d07bd828df3ba1d24db98b5f81442d27e27d3d7daa74e0fa1586aa0e90b0e1aa926e8755888476415454f8a5ee3712ca2e1cf224f70879ffa030432a4249a61ae1957a599692c0cb3c2f4a948db11cab567f8211937653881703fd6dc67aea59a5ce823c0089d41;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb54ef2591af1926fc0069b545145fbe5a9bcce3fb7ad5686390341a7f66bf636f03d0c048e10a34aa7d710e7831f11c4ddd23dcd7d02ae0e8d485be691b69946641e60dc30005c81a052f46bac459e3cc8cfe7d2a68bb4730fbd5752b385ef56a84c8bbf653e5b6083d5d0660246f7aae281356fa2773f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1661e9d8d599bb425c9a50c2b6f9ea4dfda678a4d076f17df3807b1a1ed054c912c261bf35a785bdbf7ef0073f72e0235bc9464f615aa3a728dbb5d211ca2cb196cd5d212beb292649ad30e70da10de662d7ca3b1bf6af0707deca6ad107dac929e89ba813f12b9c74002f4c0ac364eb9a2de6e003f44b541;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h125e14eb170fb7d6687750a473126dd7cd2183d6d23818547ba53857c8337d1a9e30208625851c35b78f63c44a3d45aa5a66aa81a5f658323ad90c7c761cca695c841513150e52f833c467d3a5e2b24d45dbf9c471ec5079120f77f585fef4d8deb0a3b0786e87c0d84ffd28f610eeb5ddeef5232e23277ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1abad8a98647a8c72e15e9cc3a9f8426952ef99ca56a4ba1e738b7bf063ad777d7e56f37b79eac1ed7a7d0d5b7cb2dc1d64e2838f4b9aa631ccaa566968bcbb20b5e79a78824c7ecff225d374305db2c6f311cfb387cfc22ee7b51d846a91aecf277347c31f5551cf231f6a3fd3272bfc3101243558819344;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1299dc6ea1332aafede877b33fad281b19effb7c1d968f8757a3af0a9b3e5fecb05f71597c83a448cc750f07681e53f5c4c097c4790d8c4cee182632105164c9846565845c4a024501249b9fca8322c001c0813795c7ab89f672499e49f78b24f82ece144e254231a3a16d09ab0507927deeeb334481afbe7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5db6f8099723b2dbbc62aea541e7024d73b0b4562f244a4cfea8e4549213add4f63f37a3507d4d33498e9cfba47e24a76ada0aa85f72cc2503368f535c0b574a20cb181cf4bee5a56bff03698b97b22323d272eed7a5db3e9af075738579628aaa4175859a808deacf3e0622d827665e513f70b99432495f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb449816b7effc289e73c81bb8c379520fbe837afeade849937a20f4617fc38ad2940b34a9a23c1182a6780eb0f134f0e88cb49fb1277c6e6c0701a5db3c01ab1eaf212fe54fc5a2f5d0f00f8a9d3b00f379f947523f907fac09a43bd617f844990b6f259fcada81bad8e1d589b89a95dbb9a9890bc26fb15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd173aa80e8df5da6bd5a396cd0472224d60a4e86d25e1567094021fc56195c0eaf018eaa2f91dd7bd07524fd38fad71f0409da78ec7ef4311fc7b00fe716d7b5fe25e66f097df9bc049b0917ac8ce69ca06370d4f61a5c6638afedc94943eba70c749e332791ccd97e57fc2dab6f5270a9d329f1f6f4c9f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a83fbe1c5fdfb3f42fee1aed0dfac9c65dc7bb96ca76b480799d5d8fd59fe88396d2cc6d37aa9de5288d1442ab0d2ba281b964367028432d03a54baa8862c1e15c871b0e01f1a8bfee8daaa7d692f406d9636f5315da42f2d4a39772f30633d61a8ab6771aa584633c7da1fb9a6d5f5c42d7725ee021b98c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h67777a5680c0029985273b03ce1cf9957c8464493e01a756826822b90715fbb9a74367ccbb801183b787915a0b78ac1f9f455b6965a624fc8673c6d81e4bc9e8ff8055a4cdbcde2ad41e24bbc04b45ee00608a745cd89468dcf7652d2fbbfe3c32a584e60bd4b807262705b3fb32c029844726546b220326;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5558c88609ff377caf6d442c455986dffbdd135af504577bbb69b021e139cd97f5458872f11376bf96bb607eee03dbd63c1eb8c59144b977285c065a26ff29cb9a2b4aa929aa2c1572510ebc44438a6daf0348f410ea3db8671377e2557bc1aa83b2b7902b0fe91988cbed103abe00d9a1b348b4353995e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f5d5b344603f5001200bd1ce06aaba3174ce3dbd0408bf2b2cbcdc3c81b72d22f277a26ce690a3014afcc0d061445f17dc8c06444af9a95630191d485a613beb8b300b2594167553fa4f5f1b46561fe87ceb1cd59a7a32c984dc86732685264b15e88d7a87ebe2e23b1b5b1bc19adb9ffee1577d09950cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h436047056b9d6e942e48e4ca1e39a29fce7a6c0f797dcce5050edd18bbbf4e8cb2518626bf2caa956a1fb0d3eed26de0eba1af930319ccd2900c2d4ff724c5789ce5867657929ba010b0b29d5c73d60ea6994077aa10197e24fa7dd7810565bd4ec6ae5b3ed5527bd6180ecdf1aa0db0f061ba0a6a888671;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc70b1db0a39f29e08f700daf260dfd595b2311d2a439be9fdbb1f55790f23ac10a18b65d0d2106757aa4887d8a98dc645bb2f1aee65953023739488a3ac4633a81ef16c027cb585176820e8c530817698902cbde31597ae0cdbf15ef426cd03dc8b557c3564b9a50d06d39247380c87a723f66a81b0ca3d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf636b70e4d7fc0a1dcd04d576875f71aebc0fcd7d1879f308cb189ecd7d089a9735bd0200dfd259594c25528edba26562227b4050785d75edd8f20811089f032eb37c99c60c94152e3e58d2992c9e6f00d64be30ad19f3c054c80269fb55265cdde5045858875382946b89203209e86785553e6adee6b62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7e66f271aaf6fca1edee264136b520475a4bb4371a4891b774a592fbfce5b1301f00a9e9dc7c9a251547be816e94bab46d6af96e928085ac8938e6c466439f6046aa313aa205efe9d35d0470e3bc8c6f253a0882ab506b6bb48fb39800674688fbbe4ccfe7735e3e5bb9e51d0642b0c0644b389ad761891a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e28e5a6c107f40ea169ae4f3a7fb494651ec521f0e393bf7c7291f68207ff7d9b932aa81f694437ceed4857c9b57ef7e68e35f7e35c0dd250dd2f7803564299efc43d48657afb3d40744a78bba80cb0bd333e3d2b49138955fbab2df25a3f1b68b08b78625a434bab4afeaf38fc9778925ea08fdf2b108b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef1154b86a1df7383753be3aaf36d8a5ea2f775bf14684b36e2edb9a7843df657ee43438348025b3500aaa2b34911e1e85e7717c2139c3c3c7b2305d6da52700ec377806081cc8975ad4a180d3990c3330a147dd2601d34751857bf5e8c2c81b0f1420d9350a352436d9d8e1a7628b4997bcef03eecd2d8b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe628efce9bd9ad3ebc33d229c3fbad8f75428c1844435c5fef458d7f22fbcf9bc60c2aa4d7fcd3ac0fee1e0b0b0e5c8628dc52c1f53754dbb8a72624cc776ce2e30c250ae419d1651d6de7a3a25961918de0a2e6783fe2cd55b1d45e9fa2895f695e20a6bdde8ff8de04405d48d68fad6a25a5b9c637436;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1782e0270e4cf4858ff99289bc186a231b44d5ce10fdba8c4b228e1a0f98168cb1dd8635612a1ab9fbb8c40edb9990c6c2ae445245371b0f7bc5b5428076f0673801d5df943d2a40ab0142d8f908e0ae7ae0d10bea13bd14ddf65a24eb9388cffb660f0fc7593fc71923235c3cd7a9eb9ffb48644431600cf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h53a580753e5d51aff638308de4ab89ec8625eba29ab7ceb0fb7ec61a76c639d850930716ab127e5c7eb38297075de5cd293b4d711ae5236f6c7b70991ae390c080a306f492799fb83427956d9b8f4ee0bac42e815b039b9687116c2dca7006e0ad6366416a2caffaba44fb106d11b0cde37aa19906fe75ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h965cc4993a101b4702733c658677bed7e93c4006bce0dd5936ff5f561abc81147950e75bc550c96f2a73710b3f94f4d79faa961064b5afff61495193ae48beeeff89b490b0159a2d3f80321fd3dee7f1156f8a8e25d9b6f9b3343ad60e699547a606fba4bf457a1908da84b54638cf55bb0dcb31daebaa15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cfa6dd27ff4779aa99acc2cf566684a9597bbfbe3de5aabcba7b8b645bc9b8cc07bb7fa0c2e63afceb9722859328e41d76da6126b6d858707e7f83a04e9d4393ff44b092abd6a233e7dacc8d2c0ba1b4694121e2ed627b82c6c0f00b5a361f932ef02d9779eae918a3e0ca663fd8a0e82a15845bc16945de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ad11307dd34a6ec1d428fa9931efaf244a88863b29cf5a44a4c102cf2ae478184a41b273ffe8d7fd6b9f2eb0bfb2a296a5ce6e54a6586a177e6302db26d22fa30340fc38382127840d4f9138282ef6d69840232279d19c56b581237cd3a796fb0dac7c5fefcfa0fd53701912206c7bd4c31230e1e544e63e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf7427c48f2085a1f6765b625b3faf70f1c8d16e584a1744e346036c47f1e2aea43b96c91469fca1d307721bd0d9ef7669655db8e8ffab730c9592b5daf3c59d3249755388e453cd13517cad19e342174be2049179a80fe20c6837d2541263792b24540554ba8a1a03238b036595f66b49c5b9998752d2d57;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h726a67ebc1462852f53f38496b23c58e10ba5f91ca23111281348dd6a14bc98ca1c7b1788a1ba6f3695f4a9629cf6ed6e3cc2d84a18cabcb27cb10937022c290252edb55a6c1232ea9f560fae1a190ba54f43f46bc813cbdc555230e0631633cd38469dded38c447c1240d7e73414ed4e60a85fa59f54117;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e28c38373b948ec748e54394fa100e383f19378382db49e72be2150f4ed9856f9d2c9d5b5c0acdbb8c8f90dbaee98c80a1ef269c27460e80db5937db3ca024b568a1753301660fda9c111b84a890951cf07ad6dcb3c4ea42dce6d1736584311bc3163789204d7b9c4c0e2636edfa1aaa4fc7cae9a2782d99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6075907992fd1adf9dfaaf1da3840f0ec4943e4cbbb485cfa9436c7e7a8b2f4e80583a1951180448558800c3455fe1c66862a870b566ca24991ef99765786d60de1f765433b6bc937d02d7508f3ce1c4ff39d5638bd2988b3f2b60f2b0cb714dab8a50bde6b16c62a34d4ad2644fdb3794e7dc5d8df6b70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2048445d8c3d25f483ba47a5652005a132c1b7411f8ae2fff677e057ace9549d66b3702cdcfdcc00d683b1c92071d7bc05e8373aed2c64c8337e93d04ecaf3fa5102778318afae6a756d36431db7ee0753d5ba4093c41637f54177804498f024c815c6112cb5a49b51d6744d42c7561b46161b5f23771af4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a36cad3a616d551ce1cfcc2cd179d4db05edcd5213faa1218983ffee9dc2ef6564182f3e1a38a9e3f96b5bea6c431ab9d103f6078a53ce74b222a61fd5cac42d77efcf1635bcc98093a076adc77fee6541072e0b2b1f432927fd65415a4f9b1d67b0d6e76ddca4bfde36e9969a5d6767d08ae70135685426;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a63139725a657df28951fb35baab013bb8e382924efdd892f613dc001f10f670219aab653e9f23e4e20ee391992631b4b7895fa295c78eaabde9c45fb7adfe1364a2309662f57174cf4d12af621a4a229e510d88eee584aab9578711e6ed2ce54fe037d6f365925e79609cfecee72cc4482c5260759c08b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16d539578f6a788f283cf97b93f29521f8d318e894a7e86449e2ead1acc07d727d965f1c59dd94c6a61c8d36475195ead07e0241751ca4d6320f849bfc11f7f567f16802531d74c3dc75de33023f9b9a5ed1b650dc67cf474e5b9c0adf371b00db410ac782c5497f5dd607e028252102237e5638741357c8a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f51e9ab2a6de1583a27e1cc82d789e04852042cb9577962014fc0238a45735cf2797dba48a19ebf5dffcfa4fd51865733c4cbf142975dff74c56f98a399711a8a3f3f715fe05588da9ed369f2aaa37cba1bbb8fa26457b4b925a9d5d2d8622ebf08a1962987893d4bb49e1e57ae7ebb967fb8e71609a741d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a5201d801edd2bf5bb861de16743e630c6c9309269e21e18353c683f4696d506e46d4d9dd212f164e448784d852f072a1d7a0522ea5a6db183f210f3f853621675f84a5a4fffd3f78b98af3842ec9a68a4952386b6183d7f1a5c0642889d34980038b2b5988c9a313d2e4ff775fc5bce51ec64a8e6772c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h95baa1b57f3812ab142f55886f1270a1a2d0f20ba949e3482de4e6c3d9c060ff865a781f1e2da300cc567cc27e428f79aaeda389f8264170c9689587838f58b43291200ca7514fa9fb6b5b5d31f65704a06db3ebf9ab905bcd9c9aee15395cf15c563c386871c8e1c883fca717062322b8d381834d1657ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e0c5cfeaf667228e6abce3127c06a148b342db1ea52f494aaa2839cae7838f5c2e5deb1d1342cbac1daaea39099b01df0e3a3b709d88415abcbfb1a2b3255be547729dcc814b6289c337bbf93cc6664b7fadcfdf0a30b64a6189ca26705b1d939f197c704abaaf72d3447e6add09933e45dcb7513ec3692;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3505eac9df42a16b04ac1fa0f05b16e8099240053918433beb6d155f30426d2ac5a20a778fea70edbf8726015c4140fb567f59de5e663cb857bcaf78e4f65a9f9ca4dbd454fce0c4eef418d412df7ebb7aa6de6c46ea9986d686762a2994fa0cdd29003d0847f36b61a92e1681cc0bb840281ea6d54eac7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1beb1d0d30e6770a901ada8482fee61cd7d5fbd38224348dd967892dfb37f95b60b78f858489d8df110088835fd8987d4c932850d28ebbfde6b8bc44fdd014c02305c0cf5b2e408660a7b311df499d190215b31f9d55c2475686839eaa8bb6d22a85ec2068814d6f3eb4aafd3ceef7effd3c49861fe787d3e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a3db891c477df49f728bacd92549c5eb37334721b80ce64df1fccb38a8b9e07c3ef2690dfbec753fb44bea7636d59be9364778d54719f10fa6fa60592da6fc3703e6f8f3c7c626b2c108117bd1c7b13c9271806b2358413c132dfb412eb5de0e443c4f1b4e312b12c1fb7b7b80ee9985524dd06862a02e68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19361d1d03e52a0c3fcf0f34cfa646dfaf575ae757a37ab2bf3561e2d2d7f75157292b08ad934ff5fd4e4bf916f66aee2b62176222c4e9dc1c76d0ac9f923bbca0c574de977981c412bfecb2bf50147c9095b46ae8aefa6f21b1f1b45ef98d93c8fdfef4aa79aa712d77af6ee74c60f35908ce89c509a9a32;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h138a6adeb7168ebcc9a39958d5c32dc74d4d25ae2fc64717e00375d76012b59db93ee1d805463e2acb06969469f214792d7baf16899ba3cb7fa3d5b27f660280e97cf373b20e2141651adbb51c93e45b1ac61b02e21f476463213a8c2747af334efef73cb5dd3e5c2b569775b6956063378f6acda1c04f849;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18fd5a416afa2bb2e3d981525df80267eec7426a7d4bca7d5804416c85b21e6aa554215ff694e239adbd1ccb056bd7622f722f49d2ee80d9d473756dad33cae54b5a4eb728df923d88e99abaff2458922e9df1edd78941b8156bcc03563012749a2d147d7b784fb1275af70d15457e70e026868413e1ad95c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc782e9e489b8afeb77a5b7419d6c17dd65506751414bc611589966ea7d24af08558eb7a17f6fce6aab25c7082671c0568f1a513d44dffb98adaea69751b65cc7a219a65adb318e0efb350007f68d9a2a7dd10990d00e47a36b312a1eaa421f95ad0f1e1e1494c84e7379e79142ca99e657f4cd4070288806;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb879cd314b9e9fa6a0e08f1aa51346ca1123d9ac96aec5e9aac1fc4c85dfe8ecee1e07631b388629ba4d915d5719c9ee5e2de56e314cfc8f52b3310fe77fcc6aed1d26561d30e41eee29220610a67c7ff0149556bd0bd778230c815ebb58cd3899ec90b51965702ed0e805c9a40e3d23d5de07e3c0b8fa8f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18a80aec9835abe710ee3018d0159d20f5c77ec9cb9894fe895cacd6fcafecf589dc0b01a7ad5cd1ca076edc883afed39125a59a1a53eb2ca4b973afc4cae85289a4930b965e99b706117bafa7c9a14909e5ebc8f904009cbbbe27f44f95fd2846dd28b7b2b004497a7ba453779323184d3aae442ea406cbd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha326a6f1b1c13d2babbc4a97e49d41bd5b7f1cd3409c09986da591d88385e35e51b36b454a691ca708931b475c0019b46becb5529d197ed828f4b08bbd89bfef47a62d18d1811005bbb811e435e3fe15690b719d1965654d6c6a6b7949de843297fc4c539e683268a776bb84afc884152ad92de833e99dc1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h109034d32bd78d51398313fb36dacdba7cac4184a4dadbe54e9ecb0863fe6601596de02440aca8f9b247472c71b0bd0e6ff4c06a9ec4896a20b8152ca94d52ce880bce5caca13504abf343f1819eb0fe6203c19fdd65d2b000a291ff5de30d44a96e8ef7e1ff676edd393a6eed5223d6ccc296421dc0e1d62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f9547d14315d328423e4a0e5d74cb383df1b165136b58dfa9ea55827c168394f5caff625a555de6092d096b45f943a2da9640f4ecb6ee9ecb76835f8ccb44e75a2986177ab64f7ea6b58d8a58e066418f5450788c1303b75081981ef2aa14010a979a56686148c88eb802a0f57ffe65f8c3bd38d1e8cd3b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc81f5509b713c47dc90f1963fea80dca887ff2f3ddfa77f15a668f6cceaacd3a17ca4c80d8251063149eee07ff95bdd3c0e05acdb660ff9902055c2647aedcc743c38ca6d46be72c3da150eac696c920e8cefe3c79d81d6c21f730561d01040fe931b7e032101c7945a76005ee3d0e292d9c92504ee0619;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5bde9ecd851e46e66a44701205c1730c91a4b4277ab542ae89b969eedb3128553b557bc9c55c32b127cb9ba082f83117350f9e083d1092f81914af9a472ce78d1f2e5759c4dc4ba14c70a6eaba161b915f776f2e5b175c9f7e2a551e216263ed0e6ec88d2db8de53e7ce84188b8976d835163505a80b4fb0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab530aeca2a5e351a67b26084e340fbe45724793365f94a5787289e1450f6520b85ad84feca563a6e37302d0042f698c11991bc30cb3570695fe72bff15a287bbd0d2b9dac908a690d096e10c1ec9d2cd8c88ef06e3f03ad1874c0d0dd699d63b312ce47263b6d35c39d3e956bc01512657e98e4ba78c979;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13689c7154fe27602130c892f35ae84b13b182faaf97c2e6382f58a243556c79c022f0ef0035457a3c6c818ebae89e86b9effdcc1d7438d50ee03924a1c1fa2e68521acf5ce49c31c1ddc7efaed251f38d0932715b4de0808e581af9e07e863c40f37432820d6c4a36749823805c4b8e56ff96b4db87346fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h551f9e849ca8c1e9c121cebe9c94a03d3455a81ecb3cfb3f562c2d8b607bb6c47abd9df08c7741398af1e4f268702adba720a6f4a7b2913a53b37735acfc29d7aec6a8da612e5999f10b485841f7bdc8f7e993b819d5f526ed25a01bfd211464dd0e3c0ba9c5d810713f8e5c84425ff7ff2d5219c6172253;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb2b063f9aebf56b24a163261103eb1e2711d80341c6c3d165e1650e6facc5e604fb179bc06e97a18427802754247f2932aa2dfbb140ceac867f206c400efcca3649a266409ff714ae35e3cadaf8e55b6e83622ff5fb14d83eaab782d5630c3486c3a5f0fa41234da964125725703bebcb8583bfd5e706bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c4a374847ff45698d6259a0d0d69e9e9dbdcb687e62c3dbf7ddba7af2904ea94e95fc0b31b0c8bd036b01efd44e15eabcc7d17d957d26d4f62039f703562b1fca8dc32104e152addc8f2b398b9a5c909ed8002e453e893d95189e89183b429688c70d48acca7ac321fe3997d07a106a23dbf08d12e01b1f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e8fbdd5e908ef1249caa3d83b466fd34c65a4165b845fc40cee843b9fda17cc6e418c63d57992ea3444370190462a976854c5916c71d382b6c11ed4b0a7dbabb8a2744a0174903bccb38f158102ca6321db857883ec6ee4c4bd967bc47b08c0a49e207e00166050ace9c6df2947150d7560dee07ac61edc1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h109f91f050baf8b57f9816a22a3a6f0fe4ad44aa7b820c469f277a800d48943ab4b6f60d449e670f458c7fc6d0033b3d03f31fab0e49d5cf30834387e83d45c6c27ac765534cb456927a8b56236483dddc4d726fde234d2a0bc22bdfb47f17985aaef70bdd583d1d1d09ea6d535b7834c0e7d0988ba3c9e45;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc967393225b03731fbf5200d9ef98070e03d78feb2d858b0dfe31bf2fae3455b6a7ccff13550b3e741bfb6948de0dfbb896bcbb62170d6d0d8a1f029cbb740e979c12530a30f93c3132a7da39880121e5b47f75dc617c84d31af8fd7d2d5b22a223790954db224657e928b6d1d247021bfc52636793ebf2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c8bc3ac46bede90a0ff6d8dddbfe4dedcb00610a16baefe23cf120ec3d2f14e61e4033782a4c54417bea035a491a352b6bf0c18be76869ec6b91386c801c38d781c0d02c49d5c8596b14af9f6da8efb5bf4bd7aeffd7606072fb7f00ba5ce745410f3feca411085d265c990665b39a608e9f6f14ad432926;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f80e5a0d9bb6ec2a162eb7b7c226fb2622bea04c8815c022ee139aea23ef7f026fc2d68256676d919e7bb494149f4a2afac94d6c3fc8ee7a6f609d49ab1b404ff6566755ee56c1cf1b7a3b9e1e9f6c0551e0e66e197a3c56fe8c4faa99e858e51b7f33de0159fd026ab8f29872b564c7efeaf3b6910b098f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151fc07cceba0b682eeb534def8d3c84423663de594ed7e60dfd8f7190b35053854a02aa3d8db1b37ee7297706a38d837120a29d5b763a7a80c5c16e962405735c7406285ca5002f19af24b1e113b1230ec7a949f8eb414bfb80511ea8dd8cfdbe7f5f5e57e31798a66053899586160247a0470df686f70e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8131d77d2592d27ee44378d6da66d0586abfa3b3a993fd30afb8bd17de2ff868bfefccc23651c63bc4f79761cbff393e72a986e54b0fa442e37e3a413dce04b27cdc87acee47bd4cfefddf9c204079965ac03b07a6cf4999c3c27c42060922840780f59b45dc14c20ee1cf9ce79e823b59aab164facb5db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haac36f7ba6be33002effc8ff7972475a01cb9eb7e764e6bf14f82b1f24113cfd9ce9ab01560519d7732b5ac423d645dd63591d9434c92717efea9eeeb89c597bab42a2a3556e85e2b49ab76b1277f6f65e319e90860fe54cd3dbec5d30a05d77d2e78f161120b057aaa5f055bce10603aca04688fac5003b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1243f33c579a13074008398c7f0ee09c28a735084b5656d48e91c07274b993862de77c6a410af05bbdecda6bc2666418210363bda7f766b7e55b9d01abb682d456d4688fbad5dfea54d4a318e4f981675995d9cb412335176bfa0506b74125163192102dd1b8e4e844065062ca2cbe108bb5fd8ff10443b88;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h761d8901f2c5c1f971517772264b2153a114987040a71b86456b26c198c0fb8457b4f44757bfa19ad3e6af04531fcb63a0ca614fb4736af67c9bab0762005b59a6cc5a1f5e23a843866464bc75607cf5c6226f7a95e99f51f8d49ede7c1671b78a1285c831ee5cd049ceaa7c7fef971e0e4c07abc11a2af5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f54d2c0d1244221e804d01af9b3f406b4f70fedf68b36dd5482af89226982c1b4ed74887438e4a2e7c4752781876444c9f3ea4b2e3791551f7f5fd97ef7e98ae392e44a76100467aded7f871849babb3f1b968e76b811718e80d1d24e2c7f9c0d24311c575db135c84929a840aaed4927e059f4e99de711d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha6d53e8691f12130f22c4047bb8cd94a0d19f6719dbed08e6d1a362d054d99fa9f3d847aba36c1be7f19f8ebe592ccc8c729e413056cd576680a4abb0b1b3f9fdc5b8bc1b0533313e0f346bbf58fa43f7864d2b52e572ffc38226d7132bef03b3b22c62bfb8fc42cf88fbebac277feefd3b887fd200e5836;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1619d435688197493ff155afbfc3962cd7f91a8cf17cea3470f864f7ef826f4453a0987f1bd919371aa71b7c2e5e3affb476d8fc8787ef1ebb73f388238c8761eb3fb4daa060def35ddd7d4daab275f8d866f82fde0b1131a20256b3c2f23410799cb55ddc5066cbae643aff5991a3254e69800767536f2ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190cfc6c763684b52c3b3c8fef3aa4da1ef309e322c106aa95313a9c83af302eebdefd5e1d16890c54f54bdf5c78eefc5a2ecb0380754d7002fc348aa20005686384fd9b3a0fd41e44110fef64382d60c52bd918c03cc3167f62222312a360b2be3968d9ab155219d459e1884779ef70a1aa8f6bc22f92535;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha24e50970d4485bf6ad2a5f1c5d488099a6fcf6b9b1e64f74fed7467feb9a46bc7807e144150ad6c94667aa0d54cf3342ad918256a18f4d3cabda419246d54526e9e6b0d8b99a6bdefd440fa7017429a92011bc7c4f21c3ded150a8a0a8abf6870e990e0ca2750e3662a16056c9e8bbae9d7069d255b5e20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1144440a9a6490f790a2daf30f627cafcf26b8ea529e301d19aafa06fe96645ab4830234372aac5cf818fa55a00f2090d5ea429009671cfb647c69dd22cda6e1f8c1cefbbebfa3c450b35dfcdc2b719fe529393d50203dda92ca5c99744945e3c4a91bc015855dd559ca95c92b8626c910dd48629cc93ca7d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h73529d8dcf9013b3a0c5001908bc208d3ad4f805580cdd8142e5be911607579ae28fe29f87183fbec344c7f9d04f5ded5731d9197f38612e01ece2efac07329246ee5fed5f26ba3dcbad3eaa4180e1ab3f482f8a2bf6916498c6920718b96bf5d259d3f22e0b92a7df99965c14b2307eb410573077509c10;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h962e418b1ae909c162998b2fa89e4ce4ace30c80a2df6aa2d352e9848647936b241b2c6fa1269162268bba006f9aa291c1853319b03daee9ab1630c73d391c15c5e67a4d87009c1032af287f28e728c3ea765d604de6def6a53b7425938a2e0ece280d110fec88cbbd7b7723bdb45249772e9e5755e06e88;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8fcdaa4025cbf477e0d1f8b72069f211c11106491e6268b377b3dd3678ea33027bf68f96a6473ad320536b6ed19ca6a026ab1b9f68f03e5fec7e1a8b15d4be32563a0e84f80611575674f8ecb04d747bc42bfe6ca4afe4d83df2c42c167f0d6a6667852e6e9b9c1b23644e865b1f8c23c9feae7d3cc27e56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc9f9dacc7f4155f483412c0860fbd4a87ea2a0377d0a918d55d526b17b671ceae79fb991eb0529806f1c4fdbac26565d3edc62d40f9e5cf11506985ed2a033fc33b3eb2c06badeec6ea59f12321a5373d44409b6e464d6b323bd0f27ac0484bad0749ff9a565db162e7961b3cfe078d2a6383287a9a85c74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h21086c9f267508260a8f4a3e132be9d33b135812e998b72905927eb3403114bf65cfc0b603eb6e532794ce657b173ae61e8822d2caca7e3c3dbb7e734d1bae0dcc39d4bd5e56e776e872431cb96505d5981fa4770af1c00e774d26cb3d0a04a32f13a1a59febb3988ce7731cc8e523591a3ca06f5eb8ef03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1320c3b010ab21bc868a2000e07f3895e2aeec62a4234ceca111b7d414174bd333da3ad6eec9a956b8faf9f63878ccb757f0f3704fec5658be96c5eacabdfea15826dd439154b6b8f993f854f955dc35b3092e20e57f29603fb08eb4967469977fbc8c162d56118bd13f01baea28c864ad1eacb842ecf96c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dafa1adf61d949b97146e9d880635537001f7e0d50614e4600d9f2535730312795c3dd69ebf88b215bf40e9cabbacae13df1e9d4074b15517a2e74e887e4e5efce396092a6fb195e800846fcdf0269bcd6a3f6b6d4a24e937c00cc64c69090d3a012c03af437714ad20546371eff44311e4f5932dc11b8ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc260b82c583450179b4b351dc9361114aa5c21e233a342964ed90a3a889e7f4b7a50fa7e92fefd94db5ac715d5cec3c0a6dd0d05ee656b8519b1a80ee74f75c18e16a91e4ed6a6678ba89ffea2d10306ca33336319388d6348dc39081a068989ac23d9b82ef006a17f976721037df3469e34f9402246ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fccabc96ed670ada976549b5cd850dccf1e11c7cface7c83b4ba49b7a59b6d23b24a898f923e6fff4b8ab1da34d02528c29a36f8d84dcf70a03cfce29a858713609606ba26c27055295c3df0a27a87f0e263fc5ec0b55901ac0247a40beb5c0ee9abbb33b005fd5dedf919ed5806de761b51e3be68f19ca5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h39252fedbbde3e57c23661dc437000296bdbeca8d071f87a590b602668c32bfd129c147d4469bb9750b25165d55096cfac63f05008e9014c9ac8390f78a76815872fb1a6143dd4febf39adfa59e71dd77c78bd868ca1b5c32d72294a6a35db6817e0519e6c3a305396867eebb503a20400f1c55723f67f32;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8ba278ebc2aa630d1f1a274b2e6b75229c7cae8baf980808acf71b0a12a1f00ae1a3dca4b89fd6ae0ec2bafa29d110ff701df68cf8bee4dd4f42038e8166156e1c807efb9d05abffc1a4fe483e8ce11e4e1ea02e29dda590c42e5b16c225e832e0633303a39800cfb898902ae078873b4cf5402f8faf4f3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b9a3dee3d410e9c774c1d6fa7414c34d18fe44e2e75b244ae66032f5fa2e3cfb222482bf2e95669623293199cf3be17a93ef128b0ae21712a52572c47d32b5d9ee7cf9656764bb1faafa490004719e13c67c6e741c1e6bd42c4881f435e192776ad7df9b92fabf5274d40e17a0b050e4e334951203893831;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18454a4c04a6752bb19ead29ec4493579b72522868ae9a998825176b328a6d115a10e11c2e628373868b5925a19d4ae91f9caeb0cf3f1e7b790d3f7a4fb9627f7e47df527403695d12cf9aac242b0c5a13572fdfaa7177f67e1b31e3c452f6da4e41c78f41da2fb3fde93f7d3983dee336386412dab616324;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151efbbb3d4d0e0f92acc63d6316d3e4b632da54c7944f6dd3c855a537c96bc959db757affb3f4b4ac1993c8dc2a9b40243732c6bc5e3bf6ae053d967808ec69776bd0450c631993a7b1287ca1ede4dcb93a8aca7cce1474957ac59075d854d008880c1bd354b8812a827d00f82921c088f510637ff5b0c29;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h65cf5b21fb64be508e15ada8c6489ae46315106287228d56cb713379380d792049ed9d1cf3b273d086e3e1a9f83353987cbf58110d26ae6144718144b7d1d1d5fb2465ed1192449cf25aed7b04b256a0ef53e34b3611c3e930ef6458aacb031701896b89f76aff2170afe6e2b24e5e324b5fe2a3bad01055;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2945f6d01679c089ec5f6bca49dd8c9050ce9892e4c2978aec6f67d0dfce5924201291d8161191179482b04d0736398b858d056eb9617e065699f582387dc380e07613d3c58977e60137e0843a95e23f3da4b52ae791ed83974266d31e8694f709732cd29cf2dc1f5e334323116114aab1def4125cfe1bc1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a735f06d9ab9a6cf8cc5025591678c047cd31eae7288e691baf13767aa44b659dfad76acb2fcdd1cca7d6343815d2971ea86d0040e06d51adc621b6dbcebea87c16eb88740f7d2277d22da17f5e76cbcaf212342462fafdce3333345c070a555714b89edd796a29bd08ee3265836fe781742f4ef37bcc930;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h154a0ff4ed647cf37a73102c4d7b8dafcd0a4a9f3dfd170246808cd557d7bf4fd6fef923b5cd576704a2985d085b171b1dc8000ecbacfcbfb3ad642c119fd1ee1ef4099ae6e3fba139fb528f4ea7f92b1dbbca3b01c64f93954c1ff5f6cb8fc9a9a8efc716308e2809a83da205082da6c0e82ef82e019a2b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3642bb375b206211924978b046e1ff01e2644e6adff5e39b4959b03b3e6718dcd405124425477400fa9167636c6ec5417d1a56e51bb3c7c620237739c48c01d3875853d1594dad43e088e5ba69fae33f519d34aa26ffee1c3ce7dbd27e3581b35998a620fcb5ba67cff0c9b39da2418c5b2e0275f448a19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha18c7ac9e8ff327bd1aa3c321ce4a45f82fcc2a53c563bec70427a760b5b87cfadf0a69f15be2f4fe6b8d75664e2f4ee5c2c2bbc56788feecfc0f4ce577149e12e959639e8d0d1fe579256d0254cb03ea1fc2d8836d94ad4f3adaab901b623fa6c4607dba8c70726d3be21bd2d400713806f1a652f87e118;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h994c4c2f526e986893325d75be922b3372ea91da183b67fd9428a477e3589047abddea09665e1c6a0fd2b93e3d2ff8e9eb6ed7fb47b965b6376a06d219f298d8fa7bbf59ea0a3f16bf312858df30a097158f6d08542887ce254f20013d0c1bcb4320e8b29a504cafb7006bcf13cda8194cae56c2a7a80735;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd0f80db7876d46d79b277a251f92e21623e8e5476c395ede17f86eaae09c7c9f04cb0dc00558e78a8a225c74232546c9d652158bf6054aa68f9040db6326a2e3f6cd06a6956fe8ea8efea3d98edc71cd914b37eca7e5203567f0eb589d85e033ac0eb744439ab5f7c49508a41bda2849fd4b8f6473e63a15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fbcdb9b0011031297ef9d89d50d0b10c33f41625a293cfb0dd1ac54f600c338dbbeec06f49a207771ba6143bb17b127481852c8518f042b14a57469a21d3fa2a265f5f11accaadcfd0426c8f48d43d330181d89bc42d6c848a47c93438b65e44f3e2a9c9940fc708c6dc0d1cc7a1b92ce2ffe5d02b8602ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19070342cb27ce0a89e58aba70c99ccc7c2668655b88f63ada07d469891474afcee638791e774e6befe4cc50b45d2e8317fc82d1fd4869981dd4874adcb6e4041734b18fc8229cffef0ad76a2aab9bef1d14861eddbabd6efeff9904cae175d6204a7a70fa5b0c08799d14fefd35ed8382ae9f0eb2617d49;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147215fef3cad91509921493e1c632bc921bf4bf74e0992f8634396836fd0b83bba0b1a7bc2f79d97f884988bbe3fa4efb607cf5aae49e8f38c4e146a3bccd70c0b42cb72a3b862e5fc1223bfad23ca274a4602a22f0cba1146cc3e30e67e47c480e38a8b03fabbe5c0b958db3320b7e5bbaba74623217817;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16d72430b0c1d814d4174c82702cf33cc26ff6008c5ab5aa2a425c8153ba581d3d302ab6bb2319e7e0b44f8898be10d6700d9b48249714e7fccced9c9171c9f4f2fd52aff3a748437e527722344afbe26a0294215e369b0bda2a23cedb74ab73d6fa39845c2ff9444851eca0cce5cd15bbd9d6b66da4e5286;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c2ad8a282e6be572795d674189fbd50ba46dc52dc61db775a95887a9998ebe7eb63b465c43ad8dab393a527fc2799d09d679aebdeebcc1d095747480b538c45d9defa6302a5021f6b54e9c25934c1abb358d75e2d5b0d2f163d70ef29c161ecee6ee88d910bee2a638e3818cfd49f8db1e98105cf242ac9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc47d0bfecd743d14929dc319f972d80030b07fbc1fdab02fc181a238132ca2b185cba8b27d550687540098a2f2c0775cd3d313253d2c4a5d8ac287c6624b6f904fc5b4319608ac0f249183c2f353004abfa5f87483fb5a1ebcc130722f12aace37c39791e4f14e8220cac29c48684ea5ab53d544ad85faa7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10dafd2ccab38e0f6685545a586843a9a5a84342b4c5a8cb105a0f9e6a38ef09173e514ffd9430568f0ac42ccd6d8251e9ad9cfebe319f65aaf558b69c38c2f6c2eb428d6ba3620c8949fef4ec024c59346868ebda9575d36ef25dd5d7b63dec35edff45ba94826c474a023f3dad9e03618710ba67ce0fd36;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee4ee96ecc902b5039f89cd7fc9f7371472361f4d1a261ddb5eef7a04b9672f7499520ee7e442f695845335c788dab214a59238a33f710c38b00e9fae2485b3d4f67db99d9dd501a539bfdd1922559cd478ce627cd8a41d645ca42ef3b71e3d86e27d2df98742bb1beabf91158997120faaf2cfce39b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1352607d3a2d1a34bcf0dca474e17cd7f68310899b6d75d2465af8b38455b182b0555721ea41a497f32e3ed76fed676212b06036a81074bd5fe774c7350ffd54642993ea124f9afcce0e29be919d712dae573b69d0a4ceba1f8328d6d0a78ef88022f9ff7a5bd7f6c42a6408d767d44b1cb73bf53fcf9df5b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h199dc124c005c3375b6379c383d5040f30d1fd145e6a6bdaccc4e58cda1f1cc023e2452e4a0ed382368bb628a8a892746a47307be26ab1671f269800ad2c95227846f63b7d9e373a477c5fb85603233a4a68fc68dd334aeb4b2114c72e5b6b07118ef1547c92278ecac575abcf56f59ef85b7bfbdf1304564;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157c83bc0db7d2bb4bd455e31c347061262704dbdf4210b75b26d55f75747f81afe24386ee9a7788ffc5dd85de1e3aab3528b0a449e78ac1db051e475dacab9db51c31187e2f79cbf14eb9f85874f809feeb1a38ca41a65f68cc62c806bb2ab36a17e87b6c728aab1f905c8d808207e6a011f2f6ce0ecd550;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d3ee6638e756a98c15a87a944c94892cc4db788874c3fdb475867eb8f9a7cafc71c3392af1959846c71c6616fba03bdd4b787c30379b2e3800a470e0b310b3460e3f9db0429e804e570e535b269f154819e1c9437300d86410e99d97d78c197252ca5383c6c43fdd47a26ee12b6baa4e4d03c7141fc196c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8340e421a3e62f0a2af60f27d9ecbb1165c2e09ed0806f3e9b15713f9159d3d45861d0694a082ef52c4f4f6412f071478fa15db1808c9b86e7d229786e5ddcb9417e9646e9d56fd67faeb7da302648289c6b63acba3f0f2b69ed45318abb60f9bc4266ca33732e64582961fd1298dee6d2970ad058835e83;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2524f3c5c06d257a681ba899766324e35a5f7f695a60f6315ef6cb04856eca1bfaef90367de5d17c1d8b71bce587c4e492a075616d4a4b569f7931675b528ba473b831798798618b9ffa400eb83c0026aa54ee6bc0fa646bdd8535660bcb9d9bc73b4bb50e1843f72d1425ef144294b6522d156aa30fa76c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4be196915fc51b3136866e4ebee89f96ae7d6893393c6bcaca3326dc6cac73433c0720e12314fb023bb21c690c89e8e4b79211c3819c539f165eab824a1b1c766e9203192debbd48dca80e99e936265e64686ecbfac39e854e2bf9fdf6c2bd322e876ec3f658ee2004815d46ea671f5792a605c0f642ebd2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1491c527121578a17f6e4bfd3b3a1dc54ba4cb83f27746de76e9480ec9fe699d8d3846079e279f4f24d4d34b3b6bc23b6f6d56c23776585ccc2b2eb81c735acf93effa2f95a2191706207c34228dbc6c641fd6fa7236314b6a0dd494fe67182de760d0e1f5c51edb9fc4bb8d34d103c607a66985581443550;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h256fdb869e6c67eb24b1f5bb3b50ad5831503420eb45d2bfd0d304cff5e071c3e81ffccad7e7eb6785f8addf6224310855f1bae2f25765a104ad74fe9847503aefc8aba2cc0b6c105604224544f98fd6122ad20f5c25c1b967ea25db97f8769b3ccac66efd08430d18431ca309b4c9560f71787e23c4559;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ddcfc679c13da7ed95f92ebe9685cd3e828653b79bdb8e8e9359174308f77d1c67a101001fc56bff7a01e553524f69f0e8772a3c849d3a53fda96e3be68f1d197e83c8bad5f5f993a5760d9b9a9b9e8dacb826f391e324f3d41f22dc76030c820505c22deb2cc7fe2bd1555463a43cd8ee34414f257bad9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd9728e6ee2a22831746520ba1d925b52cdfb87e72e3044b1e022ac20722b25f73a65b4d6be860745fd711459b4d8fd8f7bfa4a6425237c9d2b378b59dfdba7a1bdde359a831646d634eda43e107b4ed5864d9911cae4b2c08a2f3593e5fd4e9e4807f0a7713db3e991ed8977d421895b54d5fe11d562309;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f661080aa846c1c5f57b94d83c3480ae49fd6fa94a1c5d88fe92c4076a437c712f20c75367216694e6ccc82b55b76230a1f737b318390e25243bfcc2c6599b9e54e0653fe70dc2c578ff9ca0db777c86393617d3202c78b72d696b9fa8e93f681e71d98f0fcfe8f27fe965f1c3bd4a069af0a89c14d5020c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h487365e0f173c27a7d787fe7ae8521386e3fe61da04182f9ae4d802a847f9fa1c76211fff37f4427bfaf28f95aac815d91d724962ccd74a561a790a895e9b9598f0ad3a2231407972c0a8246a9cd8d24dcde8836deae59a3f460f7795fb04aa9815d3655d0b41d920ddeeee9160f7481edace4cf4b21a59d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2bc2c3c8d69060e0ce50b40da4681946b6d1b776c52de40da7bad5a675bd5053aecf2c34968caf6d894ab968b3703984ea45fbd0271654282f500559c3662312a68793b3927d9c3f80d0957f68908d1ae09979fd1bb76eced2bc3d7d1f570e3e0f633cbbb38851caf9d7cded8ae52f217233058a43ae78b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18da4ba3cc56e1f72f10898e4a73e7ad0a8c38013c97249b272a89cec659225c568007483e6ca76d7e973dca63088bf6615d6323d3244a14df8efc0aec27c5030536852cf341efa6136b0575a128b3637a3d88f46297f772552e8c70995c7075323387a4962aed800dcdc9ac48a4b7b267780b5ee9fdd436f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5cd6923a0bcdc79588cd5e34ba6f7142dfb4a221677ad56d46dc885e4f9734be4043162f7b460283a44ba912efe77a9cbf7459516f5c757034660522c6e934ca0cdb2fb7523596ce280a3f9fde0aa0f481fca9f68ac2e0a342125f4a357eb8dc0678fcc49d337adc984ad9cd08b4c9382f94c06214578ffb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e97802895fc2a407e302cef6d13f01e1709a3baac0e3da5ec587833e5ae5bd00e807fbbb7cd8ba9eb7ed0ac6bae7a1cb24bfbe9b89e7c2060c305502425ea186df79260ec4c7ce8acfbcd298651572c788d094658995ee3b10fb03647a0a9a4ce9022ab66ef5bc91bf688e5d9bd3ec5969ec3eaa847a7e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he35a20bf8bb1d4aafee73edec0654278546cfa46eaec0dfe4c5bd85e0d4f23c8249317a189c9090170ba105caabe9bd147bf15afcf0f1633e1b65e1f3ed8e5ede639b83aae47352096fcd2b70d34d40465bbca4d6eaafb469802a72711e36609b5670b74e755921d4e9cfcfa50673090b38bf14e69b8ba1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117b9674bbb30a84766795d54dbd10500613c1fa7eac5b5ee65b3775aff6ec0bfd7b7eb784091156239ad396e8478fb67ac5b43ddcabec4dad3be44b8cf03763ba891ad1ef0dcdf62965c70c36f27b7aa95740aebe3908a8d8514cec591a9acee29b52be1dd9e60e652c87d6cee953e5cdb92e2334de0c9a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1418c778e830f2c92d896e3262c4bb37ca9278cee893963d90293d86e1e85d6c87db156624572b7e15d07735e4328a8dcf3d216fc65a7bf8cc770043f30fa509227696134ff1a61dcf69bd377dcaf59dadc9030cb7a00be523355d6ea1f32e583102adcce9969fe1f7ac00f9eab6e51021f52c101b54f20f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h150f0286e8971eb4f80d467f7eccafa5ddb9f378c80c85cb8baf76e2e421bf825a0b8af359034ee512a397b05a74ee35a755dfba9f6071e9a458a9f1d06cc0689bce64e77be12f5a34e02f20ee025644fd7d36948f9c690eb0317cf1786cc16dcd2f8ec8cdc76370801c31ea486892ef248dadfac862350c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18450cc6b5a37c65877e12f2580a114f62f0bd84bedcc7e176e895b63cce797c00a9d59c4cddc26e8745fb160d09fda454c0e9daceb9c3877bbe9d12ba5f4fd4ad3faca97916e0241db8fa7f1b43697034e4ea1e2ca91c215e8747659ccb3b5c2337d060295d601bc2fb42240ee460b42cd1124d3ccfb8ca3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1552bb231c167fa5e93e5c831acd2ac3a6ed65556719e0d1fde433e34c040c50c6b0fedfa332e26efc8d7a385c532655043288097affc14a2b657688170bb841a46395b72381f050e64fd6b25916b74f1be75655917fb593e73f7237c05c9a3f69768387ba3fcd2ca9cb509ff3b9116f64e11f654bf311759;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc25e0da2cb8e9c607e44d051b94bbcd18f83004522852878c5d18cd33b60c8383d01cb31474ce92b5ee85a5dd58b317b71c36c2bc38ee7b2a491c5b60b7ce6133827118c05bf431bf923397961cdbbb04a781166510e1d35765966bd3db5c79e9158c815f5bb326943a252fcd91dcf20695d8bc4b204495;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h984a158f0d719ae98471dc16b8f6188a0a6f7a621c411cd15005cce2da3b8369e10848129bcbd58ba623bfe880255b6acd5c45ff17931a102d5322bfe6d74b9675bfaaaf1f07e73f9dec6cfc7eb8ff212f36be2209150694fcf69ebb0cfc4ec4e2dfed4b52ab950fd302de06fb4d7172879ba42014dc2301;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hefab2c2dcab30e73bb883855973a2ee635fe4f2449b71e0fb90c76e1a3f20b378a61209bcfee17e6db445de39bf536245980c90db1a38745bec57caf4bb616a93f96267f5a5bba8cf741dc56fb184c5130208c8d64282c30fef3bea460fc32a2c3eef65affff2dd30fdab9d692fae9d7e0bb7800ca280518;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfb15a7a74823ec30a649e6ae817c696a7607c00f491c47cd8a74009f34411db26bf678c3c2616d0ed0e5c73109e3a8b1bccc76613b2db6b7960d05a51381b17fbcb7dd7ed2bc46e40d93ec8acb3c880312a9ba643e4fe49efdc4ff7c556c3be9d2b4436a33d970ddd8a7e08bc6371a720d5ef145aaf60425;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc830c66c2231c397f2b42b7f757b7be82dd6dee4373a655e3daed68a3b63fa3210ebd2e2ddef46ec07ede57c627d1fdd8f3a28ee4350fd5bbef45ff6a6c7115f893cebbd572b1a57dc0b93ea984646bb493cc050cdbb6b8ce4844bb6f65895bf250d2ee0af498763c230ba2fdf6f3e31ea1f84345c969d2e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb06ee7b95f86e038c75cf822a1d832096620ecc7fb9d36f869f4ebb49954af209b033a462dd71f6f7be605a28f3241bc0ccf30068000608dbd82a46c1cb4249883eb5726459d13b5b75afaf9b1883e195fb46cfebad219e0353a2234db8bcaad1761f8689a7fba5cd72b91f7d83350c1ad2d0ef3d0f9600;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d9503d7d43435948fe3a7a94730b3c280dda304e2d602a1526ae970621f5b2ec978c602984387ca48cad5310ed6fb254eb912179abc90e2d0d2c8f5ae79784486bcd3c050c144e990e1b8bc225a794fd561845e6c6c1089ba43a96f1f88f92e5281a5f436f3a0799170b6e456be2f4a8a3e97b5b04e68268;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f82896550afde61bd69153cbe205840f3302a6f7fa22be26e35b9405082fabc232d658f9e73400fd1727eeb9d6f8519cab261abddbc454c90221c6dfbbb1aa3ddacf33a87dbb6a8b170ddd26a72389867f24eed99dc488872798d0076cf74e79eff78a4e1c4e3eb9d8307bdb16266dbd9d63b80add018a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h184209b5be1c58b0e454073dfbb8ba290e5ee16bc5f221f1d975e5cb5e2a9595f459927bc4eb204ef5abb9b83d56df55aabb732c42a7c9c8c6480761e7f23889ce7b52a22ca407749d1f8b3063af5755bb266ab9e70f3981a4a0a3107417322e40bbf5add2ddc91bc4c656f2a3af7d8b9a30561bc4370a0b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf4d3913e6aeaeeb309018c5f855bd6920331cb65e1e5064177e69328e826af888101b96567d665883ff535cf492b1df36caae89163201af3e676351cb757b3ab533950178df51c468b3f179955c23f4bc4d31fbb46e004d3da041792037d4befe951011ff7aacd70bdb53d89935580ab4ab7f1494f141f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda2b9fc19362e7a98721e8f984a19926b7dcbddb35c92247dc36d7d1a7e076d9b5481588f8032117149b7b8158d02bd0c7b550ed69dbd9c0744d5ea0ecef03a4f8bdcdb29f15fd1e2b32f50641ade6d96eed0a41297195350733cd4625a0df9860e1db3dbf409c16cc1ee3353588df6e1fd61e2777b684b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15d6834fab6fb7ff7aec48203bb2f25510ab1c0c18740c49aea3a15148dfde62ae71705f53957db684096dc6cd6cb8d5556b4c7e7911d98fd6c5ad43cd81ee4e88817a2b245ec256a90a4f4de7cc42ce8b15a1b6fa8b6d6ee468b27ce9d6ce63ddd9ae6d45a756afba30a6c54cdcacc2b7e71a05fa51fe2b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h87ab47f55c113bbbffeeeabe6a53ddf265fc6f2cebb26ddfb0b7b1db2edbb3f7a49270221567e8733325c0b06103040b1196576d3f5b08d5260326894149c3f72357e0c724c0d041e786d6a5d2c7f3e78a64a5e4e5bd95f6b54fef4c2cdf4ac6a31d600645bfac42bfe1c21b50a1945a1395c47a6da7a361;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10cb5e1194010a2a7b9c4d07d4f3614b32e15e8e7ef56ea9c967dc80027c0bfe6ab41103e359d83fc88c327bd2f3e0d35f3b66f681480cb70636807735b4a2b63bc939370e88f06c851c54c2ccd7deb46c484addde52382a8db2d72fab84f33ef97e3e60fc782a6f3c5fe92cc2eea452474d9cb9e1457adeb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5deb43ce012b9a7cac6cafad8fba823ef9c9bb3133c773ea3e5cb31681e6ceca87c174add6c80053b67bf4acc36e30dc5672e8a453e451ab0940ad60ae1cf6e4911a3e601d9449a312048c6b3984eddf3383f23deff906360116e861836414e6e72d27d7a00520b2dfbbd3b35991042c68270352f4ac01e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7f9fd2ef82ce191ec1909acb2e62cf3238ec882554053e38cd9834a225835ccee3c35f5af8b11afe00a906427c26907a25c573d887375172f00c97e58cabb75f74fccbd3762604888fda896269981b28421b36d692354600dda3f8c7ab1023de39fa5c9bca34af0d31355566da0ad586714de908f8e25391;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hecea9ace7502fe831958099cddf305163020dd586048ccc331da8044b6ce6733f4097b9dec27bfdb6aedd153f7229cf1270ead6afc9a1034b7e4e6c85a49a77feca473edc112c87f804657d6cea763b33983263ec1dde2341e510fe7606d641873651b45a69351ae57861dccf8655eb3006e2e01a0a63eee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173e3c1799d0fe085bc085b3bc8ccba9891535ce55a92bfbe5ca2485d0973d942d6a3a347a0774bc2a67e3171ef6fc5ecb2f4b75e4df3f0fbabd35435161ec7b11b9f2871f30479b3e7fdcf19bccef3cc4758399df414e9a760f0dbea7a4e93a7a96ef72609358a897b4f9e8191c145959497d873dda7ab62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e07f3262ff227f11f917a9a379f5b41c7401ef135065530c8b85309de161ab653c5b970bd93c4a02c6c6c28451a300decc19e99db1f4e9a637606dcaeecd66555670a71542207c5524d6c1478ff3db80994298232c3d18c007b570f7ed0da996ca0ecaae4d71bcf11f72301a90e2744d86061a8be9a04382;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18cd4e9895336ccc3bfaa6fdb96aa9e7569fcf2741a5d7d5028a770771c2cf50aa518157a3814916b703695ddd3aafa650d6cc9542f28b903b6cfcd07ab4a7831049eb1dabad15b4bd341669bbab8f76d3c2d4ca97836858761bf5f194d466f28c440953a25e7073dafba38cb28ddad9c60a6c7d62dde95e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1569cfa0fa95e620305cca086438f08788b2d482f3a9e2a2c4cc8e9515c7ffb03e0ef997712f766e91448a6ce8b92b9d78a4d50c0b341f4d018c14c5ccd940b5e54c854abbd5ecbafab0125e7da0e1ee7b5a1a6b138144bd6d57e0a66ef370e8f1f11f38dabb6cb5ec7f80eb97ce8de549d67610ba0c087f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1547597024e58c13be1f9e7e6e696398130ac62ff273fc06b087477b3458acd01585eee24ae3646ca4ed5c473f1d3bd1a0190f524784f8f7635f4f1d8a56dd1bb66dfcf4297e6276eae9e46962d701ed3979e6560bcea18e88cc333599933b8bd30b3466573643e58cb5d9b8a98f5b4e9a3e5bafff9aebc8c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h243baba9b5a298765dd816876826b90bf547c5156f8e73909a40b6953fd3856779b975e80b759c3c5ede93e74a489aefe951be7b6c2dba2ae44950c33c003735dc8ebf9f130801f9d7c4ee283d8a6eb59043ea24849e4a58c0ac1e5237936c222e761c47656a35afc7462a89bdabc1682c50f8f46af64782;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173c957d95f670a6deef0a01ff7bb6f19ade7ba47040b58cc7518dfa5b8fd825fbfc0776be904df8627efa9c80b1d94e266b070e098e761027dfd33c112acbf8ff2b2c2104b89dba91b68e569f6641f5e758be3e3a7ba74ada0f6c7984bfb025e4731f1610cd1d6a588beb25a0ac528bb90afc7141f84db98;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17d8906c7ac9b3575411497c513b590fbeead9eccb0299a651517cbd0cef8a560b1a5125c3260534bcd9a5c17afd41d88ffbaf515db1183af848208faa6fdf4a97fe29bdac8cb559ba5fa50a8f2dd7747f59381e1f2903164d7803b27afa3c16ee22862dee09e82dcec1a2314842fe93212695115a15bce02;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c577f88734cdf63952b1829a6c3e834d914411ba8d83f84ba981985873002577be789014b92b282edf58a026ae9ae25436127195880a7c279a2840ae6e842454b6b991a0decd30c88b0463b0d1a1fe1698b9d4d90e9ff571643e2fa16e040dc8329540e6c7b662cec6ce5f60fe63f9774b5351576d8f029;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46e37877cb0c9b593e42b261008187dcf0b404abad5302d7c41753b9ce879c3923e58fd44e225bd64c05c567266fd16f3b525fa7409797119f0adf75144beeb93a54309e2ed5cd09af8cc900a685acd9c17635018692eea4ba93b8c51a92676eece6ec0e02b58958694815828031768b1ea08c79b3ed89a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfb91d5cefbfab96a94db33098aa130f2180156f8a30da8bcbdcf19da13b4dbaaed975e5983d928a5393623387b0d8278ac86708368ce8b7ca9aff800d885e93f3b4776eb44acc1d73d1ffbe230b495dd3b0bb1d17556fe23c73454b6c95343fdc2a2ec353b33859764d1d9ddf9a1dda76749a1c9672fb312;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h642359d6a8752ce34ddb2ab34fa4fc0b658ff8984805b610f8b02215772f6da57ede5a63c89d1c1c91b200236d6fdbae7f2feed0a739bd7081884245be232e4fe2742f66e82f39029de434ecd67f705b8064846277875b035260571b81f3b5db7075112f336851d021cb64727e9da577bc4218603d30ea9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c8fcae8cd4eb7e087c4eb7bca2fd0820d2b5da04de4a076c2ae74712e3816568f961e7c2a95d1a3b4c10a3c70ec7e0c28ee497eb7ae52d05b56796ae76583160b2cd724465b8c8c15f832c378578ff5874e6fa03e484b4c7604cf563f8f3c70a317ffd5903def9c4ee1b50a0ac927f8c3968aa9bc40ab328;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h133b66fa7500fbab7de512f67f9a2bdde65b6967312623fcf7bfd1f1172fb7190ca20840ae848ac1a5bdc3e1334f4e7bb8789040a6b234b111005088233f6b3978356672c1ad6d7e77b2be80a3c28eb7334547a2dd96cb95a3c08cf54961ab52162db079fe94d115862e92b9a3ab82279bc6df34e8921f0f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h553b32e987b7a77c19cd29bff8298ba5dd37301a3bba106f0cb0433803b0fdeb6851a7cde752f63c7bcd21c17172b739be6cd51cea15a2316a99182f9f9c04e526e3b232dccc5ac8d28d338beeebf9c24a72a185dc4be71d7e0c0af9e87fdb6e444dd4bce2c1cefa13f8908dca19a110b8fda5e85ca2600b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18e3d435668df08602bca7105254593ac1d8e10eca1ae8dda2e24899fff56727b531f209a014cbbff3d6375e602f32aa9bf9262c074d358d88893a0c782be63061fabb21129e315d3712b0d784ac7cbecb0a075014535af31b34935d0fd934338cc553435ca57ea21f7bff9e5052e9227bf4739b51f8f4cfb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37b3b28d102253aa1fcc5777f0788c574ddaf5da3ca768af750756774a7351ede090decae9822e3039adec830f4171d7081730879ea4413cc62bcc889df897c410bf4fe00d2d2fa9e732810c46e94bfc579163e1c8712e3be11d9dc9807c6140021aa1f8439e9e09ba4183d1400ae21d8ebcaa4e048a02ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c8edb9b2aff3d0cfd08213c0dcc9d637a2cde40a54021e8f7338846794cfb411aaad1a981737775a66cd65f75755ab4ca7e6fd58dfa984c59beb7730ebb624f7d33c755603d9b92916ead00cb64a6423bda9c640f0bbc9ee816f5218d1122f16591d829467795036d7eb703b4540c598659436d2fc5c445b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5dc98422a435ebf5a606c020258723964bae5229473d4ef3be5c02b38a05a7bf0dc0b7bc15345fd02cf2ea6b182f2714648a39baa15c9016b1f333a51da50e08e60eb235afb8f99bb354e4953bb9c1cb224c0d6c1affaafd8a9244f1699f7aa29907797dbe50fe0153d28ad7f8217b62489ec39dfc2bcba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e27482967cccd7ce77d7d3e66a3071062b9657150064f90b4a4fa33e03fd24dea346584fe8e6f5282442a15dd229e1d827af8f3c4d7f41523010c4a53d6086bb4272d5f462a565ca7cfe1b07392d72b77627109546ee539f310bc0c567db52d24212bb58614476a84600d00c57e8c13a9494e7e523030a41;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'habec05c691e20c69f31db7180bb14ff2b25b505f1ca1cebfde76b34da95ae2aa97772eacad670a8d9c6a203de4b3ad8ab4d1004aeeacdda28a70c46d4a5e045ca0f821a624b41b3ca8f2c16b673681cefb46482fa7948ab19b3c51de0111d8a4b5d0ef3bb614369f404103dceea6e0c409347d2cc28cac89;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b5b9522bb6fa1e8ced7b216a707c3cd73592ee0517ae4acf769233cbb1216b50356da24ff04023071f0f48a1f8d926ad06b7db659201d54256d634fc9288595e9c0dbabab67164ca6f7d6b4cedcba39bf3a3d1b8304793a01fea5e7be772bc9b8ef981177e67686ff52613d689adec5d3a950f45c6eb3009;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d6d964e9f98a3c7621d633805cf0bc4661be2fd9fcbf184419e15d5db5e7a821445094a6f1467f106a02eb30201919ea9912edf6605bf9c79c1265b862ce686375a747d05d496147b4871d68e5724e767576965ba05c3946a2b6cfb6b55c8ed186a19a3f4a05ec2061b4e47fcd89b6767f9f51f8f3b0909f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b9d662fb649780c3f3db1cb2bee4dd8d7e227549aa0640df47ec0d04be5c0e0571974b8dccff47d60f1a71d0776d9bf8b1419f0532c366c573171b1533fa3318bbabe14c9ef3b2f243562f69ab26e5438c8596b680646985ba3dd1162f65eabf724e63cd121b2b0fe80ef543026cf32ef64eb955de9fb3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h585aca6387081a7b345f0d960244d459a86d141142a6e7f9abb97deaf3d1a6bbdae0bf90aaa6cec394b6292792233a3dfb6c365b204ee55857e1dd6c3729b1a873701a369528d6b05551dd7391a173e6c5f85b48470440a25d6d01a6e29dc581a27f1c834662fd7ab4a762a63c52f3f91ab8fdb9c7cf5ec3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha846013d574939524d55829245080a38647111d29ce3630f8f412775b6489d1f6802c536f4a7f81fc14740fec06dbf29d78cdb62bf6771c40a37698488a1dc3aab65728bf6d3768e0628f70f016aa6b1658520b221111367b7293d688bcc13d6b6e089cf49b398fdf9a1b3643c1564c868ffc6f501bea4d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116944efb659fbf1d9df410f723b77c75d92c0ec51e778fe7503673c179eec1d619d110d767224908ba90489d4a26ab787a8288d8bdec5bb526241030c9c84552e9d74fceca6d6cd32a574f529e32dc573f316a6318cb0292cfa26729b2de1945781bbab5b62a6dbaa822f895139427148183fd47a90ed6bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2cfd1c473c5e9ed99bccc207a730ec9c7fd6fd278c31e3f0ed52a20bf6c0a2b6523f1c8e5110a50b7d40a19b6a7434de584b253f8f3c7c42bf637892ec534c78732283037ceb75fbff86583fda27d2ffb191a6b999ee4310eae81b7ae9565c5208e3bf740137ade2dcfa8bb0b415d009b176f4550a81d3e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h54f388f4905bd0bf5f198e083147704750f989f255bcc89db51e9726225d544f77f50ed6a955ca827fca10da331185c217e7cdc02f3f9265c5d48c4679d2f5cddc3c1018e06badabfcfa9b8002b8e67f4da9ce67e6733539ca6d927fa829e6034b1e80d13d4c812b969f5d2bf55dac77faddc466d71735ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h23ea3b86f14bd75b16c6abc08cdd13267ac2bd59048e6bcc059da25d3660e3ff3d3ff4a1942008785d07faa8bd4e92aabe50676482c0fabf7d037d8220469374b19b7d85f5970853ddfa1702c8c7fc076cf33cfbbfecbd841c362ac434605f270f6b940ab4d24ae93a7ce4e0267734d461b3f9071e7f0f3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfecc2e197b38de0ef614c2f55c5c98879b439793e77f2a18f634d19b8d2af3b5e3ef441c978dac9b28f0a89c762d65ac19fe4a8f2048f3f7c95ff98289129dbc58aed9222407502eeff876d49ca5a4bc37d00cf1851d3afe654c236d52eddbd7a9474a3f2db47413c2cc2b15893be5e369316d6dbca840b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f9edbd60c00ece3b03c1d349b28e435bc21218468b80f465922f2a25059e18279f0098d3ad4f1afdb50c7aac6fc2277468fd2522b6cc323aade8f8ad76208a077f38b83f588b0aa9b3af9219ed521f1055b1689a3224d1a37f132ca386570c1c96450a169b105550c7cd28ac562dfef9af1aa1a148db1fb7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h95c62a213ecdeac83aeb40df4cf3a57ef98ab3679fd776c65e77bb8ef9fe8c290fbf56cff1149980a6b1413c3375b587d93a8e0f56e488bbc29d25c3cc62f4f9d0656571bf570acb20dcdefbd4058c4a84b83a577f3984e4d119f2b85df60b0232922e6cb2bf398d9e6dec5fc7efd51536493e9a0577feb9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hadfd81be4efbd7947ce02b0fc961cb5ee41b6c5b873c7df65abba78f946d7109ec1cb40763d81c7ad3a9da8bef3c2fdae217fd19df46e0fb3d71e74e351155c932ebff72b742cd8d1cb4b5e0457498a177c1bdf53c925cc9ca791a2bff4f89daf01ee5665c5d44d95d1525879c1013f61e8b98d1da350d4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ec685ddfd630480346f29e784b9af2eb55b71cbfd0e73a5e163403e59e2e70fa3f56b63868a58b38d8819b4c0451fe6eeb39cc742253906e8cacdfd4a5e112f1a1b69ddd40cbc4eb5ce919c2c754699cac02ae7a4c01a4e3829e62d0cd2502e0839dc76e9ecdc5e265271d1ad6ac5d918cc761d532eb4b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3c41d0360a32ec14419e643a06d99f2d5c8bdfdb73090a3ce7783df8e3a043a58f8d5e76494b7a7d65a3b6a2bf2e1483534421b66c135ef7db6dbd20926c6f9f019fccf347a754375d087e62ffb3c0505aae571747d2b32cb6dcdb23e2c2052cc3e92758e5f072d773b7cd8c32148ac4dedcc3c1f48c76f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a77d5b128cd8376d2582cf7fdc5770994ef3342260eaa5c91cbfcd9495b9b375d1b05c3784d5ea04bec9d8c2c96736168478a614584bcc8b4278f14a75497f1ed68b67bfe614fd56fd04b859dd12b68135ad83283fcbd1c4535140852c95f9525432ff11917b41e839b00b8faff9cb6b8074fdde71057c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fb77b1a1f2b211729ed2ff6cdf34df9d779276a1eef8b0e3b04f3b9f5f96a9ee642fa3957a80c71e057272a604d5728c536a157f489a944f04299498036bb5a6eddf30f768cc752e9919e58da9d56a20d8830136467c5d6dadf7e2b546135cea23acca5c0fe01b759cb9181efd4ce618604df6e84cf9f874;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b28907e8b8415a88c1f95af0e6bb2d85b7249d930724cdbe190675cc3f4335d0ef99b901362fe12fc364298308b6ea71d62198a8c19fcee1d30712d0db0ffa193a7af64eb2655c70a66a921da6665c94abcddc604347253b1cf26dd98e97dfd29f0a9a51ec52eb094d0a2fa08c0ec26ebe623c312598a2d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1016e629017107969e5bc03adabe3558cf1b0682fb4927e78ef02cc0b4a653c2dd8a2c531c6737d01fd2f66f64e8c7d15407ba1c72bfb943de1b572301712ef1e44e06c72f9c6818153657fbf8a196a2495ca721aef295ac6ffb1be73b993683b05691a25a3cfa6e53fcc155b4037936f90dd927470689f4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf10df8c81c655bbcab9ed0951d680424a4f502c9c1aab507913e58398e9e21dded1d813d282f2990291e9927d1ca40f3cd643c1b5b595249e37b45b3d01665a79f24d1fcb3404da22ef8993e82d77b8b54bc4023143038438f87b215f56b911a3d2084d8cd3e28de6a4212a077e3ffa148ea21d35a728044;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h65af3b0f804742d65a30726da298437364c763183993ff035c3a5c3861ab6c4b5fb5ac67dd9336efb52c8b70502b90b4c0bb89bb24319674fb8e07292f5dcb0803a608c234ac1f6e99620622b67c3a3f3e8c33d3a5cc52824a68b40829d05cc8069b44b510f0f5f55f7d51c3c3b42695f1340f3210b0bc8a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h134cfed6127f826ba27fb816fe96e3cbca88480f987392f782a8ebf9db3e2ac1b8f4ef9acb20925fd3fae5021b5e2ac48de77232d64cdfa1f7915785875ef994098013a1e1a9792ebf33154eb921c7cb537d596a4c42992a6e4ed5ed8cdf11524ca59a3a7993733bf38eed836c36e555418669d93340d76de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19719777e3c3c74fd062aaea0f87527e85ae709a0e519d71763eb8ebfab63afc6cebd8829de359dedad0af3d8fa57771cabfca14573a81647e8635ad6a7d296f5e221368d71c2a24897f142ec66c6394e9a15c04ec5d7124dcecbdb81e45576db169d7cd2e4fb2fd3a9c02649a4bbe7135ecff0e2ae7584fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h73215b9dd1fa7d0a28547f9564a1a06b7030cfb3a75d219d496b6cb221b027d4ffb9dca523362c0fc8d26b5d6166aae71d8f6805472e72699a903f9daba0fe9876b4ab602a75f803f7b4dbf2a936a2af4e6de59e394648c87113e91c43b5e7ee7d5d65e203c1533878d50d495f5bdbc2d8ea27b9e7663642;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he169e4361409e5b6b5b8de28263c2ffba9d6c17b4fd0ab8fc6295c5965744e8be96371451f189c3ee072fb2e04fcda2040faf5cd00861b090e73b9b829d536c200594794ce0e86873329cb9509c6e515833afe184c4df94219866e48635463f8dcdfaeb31c7dd360250e4e3ef635a7af3e08729ea5a0540c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cac586c39c3908be36d7abd3115b3e9db19210d548ca16a23b6d5e38a11712ebdd2fdd0a984a4f8e98621a26dee7b3260dfbc830d01ba1d787ae511e8ddc9509c7f3656b451ceb9dae8689a8d1cf5106f5c5837c3e9efeedb0c0fc1b404acdb0ce384c5589a3f1a90c34a403e6a6d0f703b9b7c2405b1496;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19ee629498dd6351b2279f9091ee13c39fe4177f931aff73f4d79e709b6249e7b2251ecf7cb6eaeea6324d69878adc8ccf7c20f7c21d29b4dd436b2fd7b1d9f9d712a9b7fae4f13a8d294a5e7a42bbe24e9e792372a6cb88f1b8111c844c526438362e863e7ed70b62a488125d8c1805d4efeeae13f2d88e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h161ab950d12f008b2541fb9cafde4283c6b5cd18a0c2d5cef4c396acaaacf7bbc85188bc5bc94a8b8c1b5a0007bd15253314b7f7097499a38f0b8997c21d2a219a546371c051d4cfe3ee05abf5676e846978e1e93f034d062ea23ab11e4bb44b463726e401886e7d32517bfa48cb2cb0087276af15d32e1d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10e5e44bb3edb779474f2edb2f6eda8b9bc65d172cb57406d67e8b155fe5a63536e384fe98a38b4a141c52f58e0cc62e3496d1ad075c43a9dccf7f47a4d211e48c8a8fb634742153dc2875d50a6235ab8010dcffba545fcec202b205ff87b1dd4bf0300e5ee38578eaf71119a4eeb04903a602cb6eb440263;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf2ece9e738d1921ba4d45dadd11b073fd184fc6958c7911a371e7c14b6b0f760df31d08f82eb7986d32269493774343fe929cee7aac12314164e38abe2568396032887eb3ea62d5b35e2b65127a2dae3bd3e742b2751f9bc95b9124e3d2b4172741d2f49e1ab2d30d63db3673082cfce4058573809ec7d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1db51bf8b10adc456bc2701e0688d6534279706d5a01c66b69cf472f5f44182b7684f98cfa644d03f66a709993441875a7e479d4d6e88f6892dc6f32dee7f597b97d3179026223eddc076488115bd40423972cae55a4563759e9ae02c59709276331793babf0718a4e350ff6792d226f71122cb5c1f7b3b28;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hefa8ccb064a09545d9b10faa6c22905d0c12d54d1a57c9e8fca11bb87e39cc0eee16353062e0d10711c78ef75b712ed88598858fe973d0ca9165fc70ea88192ee9077b95b5b5c0b8dbd396c11aa19fbadb6285ec2cad90bf19a99d3dfee0cd5e9737db3512e64adcb616caa0f051c21da5038950d281bd8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h48ffdf3a8b7cf5f38b1cb50faf0022ff727ad01c34c562cb00aa86cb6926f9332814ef00efa628927b88b26694331f5a10772feba67405c895a5f0bb8ab42fca9f2739c990c6d3e935602a4ffeb1b0a9982ad967138ddaf6c43906e90548c2a255f65c77f87c366b3acd3e7a786395adff51be29c7da3a99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1265cbd399ba57cc48d616ead5c73ed744ce7fd57775a4e92ccc9764d48c54dae3d94e79ecc8a4d33799d85171fdc264eba2718e38dfa2c8e20226a5c4976ee48abdf1286294751e98c46f0048257a7d135ec992823d86e12107de0fc505dec818eb073c2c12f5add6ffa162a3ea8824c968a8d8b5314a2fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h183da7bca7d0b19c322326f0dc03720f90dae8904f185a3aebea0760561f6bd65d74a7163169e60a10c0a69694975082e4f6d62054aeb461eb57080b88d954fc1bb071112fd0322ecc5f399b94095949bc4ecd6ace01870a317ee82f9864ef06fec778e54ed54b38d0545c1d3bef03cb79545ab1688b8e650;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h123d67c08dd69663cdecc3dde77429f1c92d7c80d4b68b5bbec5b5f5bcd0ec6bcacc07b8afd57d83b9113616bd5c66e3788171c863d489904c75ab908dbc09944de68696e89533f11bd5e7cbd6e74e86c37c216c0288e2007242f0e1d165c53ba244c4713cb692048770d838ffd9823020a0e8116d06e7bd7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc188f7ed5dd54bbe180c57df4d922e4f70f9f8b93f2f0e311eb4545e37508b70c8ba455e352be13fffc058ace89fb2f5814aeb89b0f30353b605c63ad6a8860b8e2ccce9bba54b8b9592c0f5168aed8bab9c126ee66468631bc02a7b3ecbac4c11ada73007851d4e09814d1199651d27903e31c8a127fea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a986bf2b62cc0d0df12ebf95750f25d32ff537c2e1d7d1e75c4d1e9e4715b22d97c02be36e6967ae6eba1f20bd429da64ef064c4e619025184166ae9df491e62763fefa030fadb330e15bf8d84558b794aaa28fb83c085e8fe987d217c2ce099e47a250f80e126abbb1f59b9a54dfc0edbff05666cc415a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h49b04fb72c1c21396ebc20ff598c6042f2c1a00e7ea502c60b9607b70b82420147cd1efa48957fdca3580b2b40c29dbeb31fb1417ec3576287b1f38c559f9c4fc6a67dfd8a820c787c28610a356a30924f196d4c2e4e0112b84fa3d6118536719b1983a5210debc4ac36c3e06e96faa4b128c2abfe516e7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9e84a9ccde04ca666664d2dcb7927d96664ad718a9c42e08b01a7b2e42d048147b741d5d2b20e646fef38d676edefc9a2383dd6038406a54988d1c1221620b584868a3e3808960e208379bfb6873d0ee97403449edff38ddffea7f53b735d22acf502af4dd39d5adfb91e44cd12607d5b036a6e790bd7d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4de103f1eb6be50e2350aff88ddcba3104de65942ac4e6dd93401d8dab77134e2b600d8e487fb2f9138d91487c205184ab2314f5f5e107abb350a6481065c7829ba8cc456f2e9c31fe3cfe3f8c2d6bf9e884d9ca4972d3d824053b17adafc05cb55f7f3c4cf25a4df9e5a6a6385f152bed45bd50b0014ab3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a674324296e17d87a036990bb640c1de983803bb545cc6d70e63cc1138080e6241308e7c9399bfaf3b890e3552ebaa0d583be001625bf91237a60b4ca4ae07e02a8f6f3ac917a347dd13665c60973724723e7c158bdf2fc0a34a121d9cf713c59dbeb8a4abfa80a1a8db47d9eef8c4bcb3d8cc3ff4a2bd77;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117dc02a0de00d1d11eb6ad5baa5006fd0df4f9fb0800e53561ee05d6277fbc9646323d99c073ea9d93c6a1a513748418f379d5e4ebf5cba6340d09b557d3a4d16563b343bde46449155d9b088fd21a8eac232045259e6b46302840a8852a4c150301a12c4ac0eefc44eff03883116c49c51b4267a38f95a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h176410e5795d3592b3c2355e7197f631a6803852abb25d9aac1a1b268ceaf9a2d5238f813214352cb3c9d33bc6dd8de516f142e409eca74ef6eaf44dafc874c558d1857ace099aaccbb4afab6daa0475075acea98c5a5afced173d559f081c8eb511168686ee4530fcb1977f73e9374eaa2ca0c756f291cf4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a6e2430fa8d47ce86054395607e5e35e376f9763f0451b7bfb2115b6b86745cbf16a8ae54ef7608ae16363457acec86eb0633d04e8b260b12d48f363c36c9680f25ea08781b5ab1a61e06cdb2920990c81e8a4f80d63fcf79fffcf51ffe4e10e3b6a5e831904080ae3c913d9d8dfbb797344ed53270fc15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h178123675a49f42efdcbe8e9d44300cf533a6d74d5f2894adafe844dde9586502fab2476f3f1f896c6b37ac1053c1e0b554c520f72b6880315e199440fba2c96a6eefd50a8d64ac04d1ea7428db8eed30d011862f7b9335349c79fe2f57c5188de0f0cc8ea63be226afa415fb0783c4edeaa07a30f2d3e08a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc50aad1e9b13c4bb614697017f7adaa64ecd70f4c03187b512ecd3cc23948aae35fed42008c576df43299ae974535493f1665db6b3d8f3a034499299fd22f24e268421f9707c1354e7482a15ddddd4f7c567dde1431c3aa2c4137382314e413e6d9794c36101efb0ae0e1fb08e3e724840ea7b57d2de64f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc19b03f72a8b32ebe31a7e1865b3e19a0db9dd116611a4d3ccd25d1fe9658bdd7dde0072fb089fa166fbc244f485d20f2e312152534a11c678beaf817428e482354d1f69aadb61a67357f9cbb19ceb8a02fd282b5b70b272151c8026630ce63806020678059ed821049ca6497cf2b6c070301ec3350fb56b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aeeff9f0637f9baa7b3f6c9177f2bbfa270e18b022de1eb439ee88525ebccb5d07b68ec5bb99822e1aa33bb635c179cb0d70c8fda54b81174fa505caa40bd8867b2c2be358082ac8f6f7ee85d4a381a2fb15a95710a00ba6bdba523274176bbd767b3a5c6bf0181d19c0e74226ba9fd9fc20082f44fef92a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5bef581640a31bef552d014fb0791a70928e40e49ad44dfdf53781460e161f60e495254c085c312419aab828920e5f03924f70812ac760c9b9e772281a7058b2d1654f2edcb8c42fe94f87ff297768f50cfcab24c19eafb551698aa038ca90a7bb5d91a3dd26466ad2a36bb38d966e189f41fc3b2a58527;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f6381dab0e0a7b120634109ef69c143099045b28d7ceb1869a531864e196aa86e6a587ec5003f1fb2d88739d82dafcb2897107e023018d1fe310d55616972ed2988dfb9c0143b88048dbf482abd024b652c6897779d154e7f4d3df923068fa2c045049670ebb6ae71dd2ad6e39829318807d768e98e20b75;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c69c0f8cce54efce3bd6d10f7b7c3e14e9d56bc21c56c9084e3f1d80b16fd44acb6731881ca21f4f99cdf6645d1ff4797319e54ae14eafaee69b60efd8ab956fbac281d1cb35a112f83cfc5b83b40b19524417a7532e4cb5f10fa17225361533a80e3eabf18d07450bfc274de15e455a81a1581a097b491;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a1eb327fdb1102a01686ddb4c4d3e78c924f9e6f4a864f1cf7bf1fe0d650a9b7c995d5fc43dac80ebc15699b8b25057d2fda87cc6c22c9acc54631c54894fc41573ffb22a6e1a181781b7a6029a324da69691425ab9d6ca7b472b9aa8483419860929542a865cd2f644bbaa93299585ebf9ca3cde64accca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h780aa4e9cc99434ff40a1b99e1631b07501e788e443f59e3f46bc3a77d1eeda319361e179db8788726ebc39dbf62457c903c975b91feb9dff161fc3d314eef52a44e2441b9559cbeb257fa5a957b98da27b3e97c1de3f92c664c06fc12f3e3457ce87e23b9ad23b4679e1d7e38af306edd451a847d666cb0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a4e67c859d318a14b71a915acc803c927f1ef01c4e8035cadab7176722e49073f33018703563c235cb652f528c0dcd7a5347dcd26cd4c02a1b550918def342d7bc1048a67f3b037ad13b5547b4eabf727fdc1323f0bf93aa11f902c7abef9c53a5320bfa9eb2c5ebf75edac1f50bfd53654fa3c6cb2535c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1164937ca0ea89b61d74f3ff9d41652fa53d0c4a4f985da4c98cfd9a9725d47510ff0a5b9cd62ab6e9f41985a04c2e7b8be697263a584b7992eb25141cb97adf62489818c3d0d9de9f0050cf617a4ae804e88990ff7bac8c1cd88dc218dce07b5936526cf3e475005a443f66d2f7325444eae38a7ca8dcee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h166566598e019122068c0b0d2227511938cdc0f0062cc9eb3538cb0780b35382607b37be2599cc1a3b977959bfcfd05eaf6ed8b1433af19e884db5e2d9f631ddd2413dabd329fe8c9e6da58dbc7ccf54501658430cf99c69d27c56dc26e2fb9a98db669d1e32028d2b1d5e23cbe8e05930f852a936e01bf28;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e416a9c12507bc30c294b4091053f20e9ff3cc2371980de56f628b94a4ce2b71709ad5d7b745af54db0737d405b396025763bd2239c15330d862d0946cf943d347180f978709943e21aebd03b3e6699193d31e3a657bdbd32961b41029c187b82433497be957282a0a9b767fa0ce781eb2bc201be3f2efeb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h129a0dbc0788b820bcc94b9387a399d63d689eafbea6f3eb01f7e1e9c93e4f67b82907df87c0f5c0b4adc41ae5b3fe961b40237793088729831be20b01b4bcc374025fed79e11b5014b37fa4a9afd645d31e4a214afbf371e480811c78027b24c935bf00131939c9f7264251a74f6a96736969014eb2d2749;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12270370a29df99926eba890c878e7b4d4b78f2ab1383ce46d4e13ba9823a953c8514c41523df5e2ebe3caa6c4de14d18970aeb7db8dfbbd705374097e64689301ef516bd645f13022d3e4562acf9df135aa325416290dc2798c41e300e8f0e9d66af815f47e212579ccb0d5eb6972e564bafbe9845fad0f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f77d55320c78482558846c09b2fbbde1618ca2e7732bc5d119bb2ddd39448dc529a2d6e88c9d2e36e0ed65a80e3a9d741dc7b4cf5671c81e93f38dbdb6c90302d712a23f8d436252189d0695339a3108249975db9834feb2701ddee60462eb5d468360855ac2492b0386fbc384176cf0411035563ebc91c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heae2fcf13394aebcab0034ed725824581ca7523da22fc7ea84e4ba5d61f9fe04239e961c76e5124c5bdcb922446df6dca18f2d50bd5a99e159ea6b18058bb8ae43b4dfed34ba32b5b86a918e3f1ebf0bd090fce5696feda4eb09ec8a180d367d47ed471cabc27c1791f40c8988629894b67e2a3270248a2f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16374d25cfa1942371f83e120d0c94cae225bbf9524592d4f5bcdffbe9680460dbf269de91c577004b8e5a69514c48f0bd9dddd097cce00823b50742656f6f31b26a096025fdd19f4d6bf9a4b1700afe003e29b6d29f417d94efb30ff13e55736246a6a5133bf3d7442570e172257e8bd4e16bdc4a9a5eb7d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175242b2c8f2867a4d99fc49e0dd4bb4614a46c99863a83ed97ff0b23fb775c7f3bf058e311d6ef3b6fd06d924c651c0d3e59a81e4426c363ac19f1ecb5e1403389582e2d65065ca05a975c4d61cb828963fb87b86f50682f3a7f8d18c6766fda6ff112be3f1e81cd49ff7629ba3d4584ffb9a88efef8eb28;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18294b031ac945b4d811605b227fb82f1fd94c6d8d15c7329284252400db43b45e4ccb1ab7c3a253e26014a750e00d53b1ea8ac40b1ff63a64b35885f8c263564b32d98321e9db026e92f4c6d241a09b7ee38c2fced434e6d5a8a765523a7379ade268812715193e7c47ba6936511f74b0a140c3711e33212;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bfc255707f7c7133b9de0d3a96ce1ae76bb475809fc480e8f47e553888d1abb8d3c1cfcb9642cde520f114828daf8e2a04ffc9cf977c38677f3118df4bfa37ee83e39d3c12d732112b0f194c2c514b6c026b256a44eda102edab378f271aac308901c8dda41bbbc4616ba3572ecc0f8fff7376476e7a8ec4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hab4e8ad557fe7ee92d479469f397fa50921f15d225264ea5b6ed926b09f8bea17f8f1eafdfb5193fb14e08d436ac49cee4576e29c2f57494da97fb4ca9de7e0f5d397a679516de39fcbabb1667b815b435b490874556ac206b2f988e6d9fa3fe77143886c8089bd3bc9175cb538f1973d6f56b00d2a7b4f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2dbd0e3c651e26857160a093caea5f605e7a948d625cb0d5ad0ee91425244b76323ed0ad89b657fe46e5064cd9bafbf55cb5160da3b9cd044595db9f20e2077eef17b4c9b4a18ff965cf90e211b796d7bc1574780f1d61b360503c7c29d04342e42acf9b9ef68d27fb50f3874adb96b7bd21f241cf6c96c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b36fb8bf3686cda2300a28007550e50308faca7a16f4d9ba2718ab22fb8d21771b10212893f4e5cbea82cf2f44b82c6b3bda6419507e27e87757b98f7ff5efd61f7b305b5b2c5f59b50f9c804ac426f0a059591fbab4230348a655c5f803ba84e4f094fed02a7389e03189d861d1aa07ea86c232a640e15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d4b4e63b72e5b5f5604f66aa378eb687c05417ba56ad2c65719b4746e1c9c854617f594b1ea117f19ca01a058fb3145b2c5f9700b3d06d4d628f8a603268dce89871a11149c9286d5af0e96d371cd921ea66184c1674e8ee556c9c45b664a0c1f3abeabdfc5751b932e88e38f9b38d010fd391f95f2e96e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb62805e191dbe6b579e1b01ea2c0a7b53fb91ae3ac756c59d4936f18c669ee8acecb7e1aea40df7a38f5ad2a29e16ca7917a970624b405c366cd35ec17cbe8dcfe0e202bd439cfbe368207c4da30e5394cb16bdcb13919cdbe2a7334421841f96484cb68222b5f811b34c05ee0a13c599ab9b2ad6b6ce1f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd8244cf8e49c93501f3a15c7d27d31daf4886974e20084e4ba02ecdc70ae1aad001501f1cc00fa14302e76d5c7e3d6cbfef20f3d3d14d029d0bea61f98cf648f664b997a2a10e7bac2fdc68ee10403c57cef4f531c7a9366d58977aecab800fa8e4eb4c5285902247366247cc69837370a0b0232861d9dd1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h131622c0851351d526a55817a2fabcccb99c10889186874ca2cfd0c73f748dc9f575826ded47d8693064b2e8857b6a9bcef1b3cda6b7abf8eeb3b6a8e0f1ca440a5c4a0c80f7ecffba3e514c57a4877c030e992ad3c1b6c5932000bda6c35f5add80f64f6006ba3fdcc2200a65dd22f37acb7e58885babeec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11828b83d1c96c4b3fcc63dd2dcabfc453cca71bde0ac156987af685b77b21f7c4493bdc52492fe3fa8e0e6203977032e9a4f20fccbcd098612a12b3c08afe7c3b53d75252ef946ee0b72c5831b72fb60c17d3246e78cdd2d1fcebf0290b0dbb8688d9e0dcf23cdf078ce62ca09cca7ae878bb3b095dafa09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e0ad8fea335e03c13705eedf56c2df29f3fd01731b8079d1ed2e57ed97da3547e5f53001efdc5e17659f869ca482a74970878b5b419831ac11e0766d2f099d5a2af38ac1056be4a2a0844d4f9460967e8fee05bdd2e8df744efa6c1555a4325f7689b50f186033a9c1c0054e0ff775205357582ef5cb9bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eecf62ccbec6ec9c735eda89f1b880ef8d73218c4e330103c608245a47b6fd14e5de159cf0de84c4d14000ad3f9f280d49ce5925592353732082e3ef93c5a0d9cb53bcfcbac856d8db211586e296aa8ec0995d599c0d2b47d69dbf0014e3e9ec12098eaa44188298dc82ac54178dc53fd6c5e1d723765ce9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5b25a45eb0810d9b973b514586cdc412a118d6dfe08a7c0d0e5a2e4360692281a13ffb20e2260d62e8c737e04228189eb4293c1cef8aa46ebda501ed6461b6176b2f13b6148dfa30d45e1ab9e0d347a54186830988fc1765f2b00fdd3253dfea45f3ffbb48512dff6247c0eeeffb960fdafcfde83d0bdf4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b8c51334caf8bd5d537f491f648d3027043a7e46d7768f250a56f3c6e095cad36d45263c5eaa3d0186a72b09d8d8e0c1e4b9b911304a5b35eeb21b8b63b58a01c872ed350515847f2102c70f89b83e72ca061f3210725313b0914bc82fb673ee5210f0bcca6282c1a1080db02df0cbd13fd93e2b7340f5c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1682e12682069fe52d91ae2dd623f305542bc733d70decb8d5540f62aca205ce9cff0b3f5db3ac2ff1d110e26f7fb2c5776106d200566d5b777a2f29efca2a063144c137995add8907563bef1fe172e7893c87512bbd0da8537c7962235e8e477cdf72119c83d8f46b551104f92e3a1f03faf2728a65abe2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb9adbb08995436e2d6520e3c7a6998dffa7050afe1c285d6beb99bb8cee2fa4e65fb2fdb280ccd7ce972cb7a7d962363012cfbcdaf1fb3f7b2293454e0e2643dbf4149437eb14a3b7f8e4cbabde6bed93f40332c28907a6cd4f40b0a5f69fba75738ed358d93e1d2e2d29e1e335ca8dd728dcf42c99c67;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a00ee36e755358c68491ed49c1fd0211a29dd89f9de7adb6aba4f960092797ab9bff197d5e5c1a36b3cdfab0d532ad173570475af0a2f6078feb5d28b3da3dc32e158bb222e81001aedbddb757ad259869a9f5377a68afd61ef1a4c4d16df045ff5964fe3f16ecbd3ade706f7994624c67a944e86a5d8d3f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7cb17a1f01b2821317a860cd2bdc68a92b3c0a498cb78c64d9ee5a7dda4ebb2478ec7c5388bc89adf4105f39fdbcc8237af7dcbb334ee898b57cfa2203ff24ca6cf4c88e83e5d6b3b49cc89789948edc673d51c4c45d1cb88d13ccd247f5ea265d9ba0a7d452bf6494631ecd19b0889ce22a2fbe5d3b9994;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h152d282731027bc2bedef1dd54d0ff41aed691a1d0300ff960b164dbb4899131d358521a0b02c0c25776aeab8e4c1b598bdcfdb3145bbc68d63f4fbe6c97443bf73299aa90977b6f7d72c33cdc36188f3a85cfd6d8f32494c91ea6cf2f9fdb3a6a9878f457a204b4eaa9728beddf87a01c3fcc268c33375bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c7cdcc1d4d837893fd76ad14b66d7d230ead1f046655563fa796f38f5128338e0506abb0a287b58cc0fcb8b4c04c2492156bb9312fc1e85d4fa0b33abe148aef71f199f5ef9cfc045587cb26b2eab873316a0117c4001c9195e34ac5a7b876283aaa3322f4c888307dd9aa4552fbd9a003df84fc88c35f70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h22379952ddadff8c304b5c6ff1f2ac19e44519e600570c93435c37a7d81dc8a27f89650b06da6046fa13957029a662ded3d9573e7d481cfd4a7b4b09bc08722a1eda40a153c8ff7f4f2487880249cb6762eb7b402653099b7639d0853581d41ff29509c34bb39bc5e211aca90aaf1a3406f4a9cedef837d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb57f017f883669eff32e7622045af0c9c9f58322cd5527961469a54ea5733be682644a75103eb6190e0073aef81fbb5a922c2bd9bee237fcf977f3c188417476a6f3e7702343c1ef4e2c32820197a1d4a4ffd4cf47cd8ac224d9a66460f46394b39425156292fdf8ae49f40126ff2d1d00de43022158f05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6781434316b7d6ddf048a91a4c5b1c9659f0bee94773ab93c827159516b064fd1e718191370d9941f16c9714299acbff1d13d54c623b583581d1369cc9fcdc4ce8c8db48a4c14bc46f572c23894787cbfba6b12c68e46dd96d927e48a1e1f3235f1e375b8698d8c0e129b6cf860976cdd3494c82536bb0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h87195640398cce16b6763a351fc6ef097fdac5b8a985cdec73d6ff3dcc26e9244df2eaec3d2046e3d9819931b3e12b67dc701c84946fa62b2bfe8a77ba721fa854f3c506affc3c9d63ff8eddcd6d67fca2055c17ef65d759e92b933abfb6f9c3d915a1a4c8d381216d7835a60cdb592966e9e4bc47c98c63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1590a0e8b6f9cdab8b97ee6e81ac6bbaede14c18f47ee4f8964ef1399e17d6bcbf469f5580e23ba21e00fe9ced68662a1e6759cb5745966a8a4663b5590f094d8ac8bbf2b4b0067fae33b26b39a4211875932cb281a3781d944fc7d232ce3881191d1bdc6d3aa2a4306955e31a9f8f9d3e050cbd35b7b0612;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19cc851ce22f33cf5aa1a16d46c2c370b084329f1071e3aa96163722416bae2dc168d835ebffa796620f5ab35daf88dad8f35d4e2eae75591de2b678889ecc36e9af9eaf7129c7003268f057f26d6d6c044fa6ac4db438e92f8ff5da7f818d038d0a080346f7f2a0086fa848bf127b03339991119571f8432;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h702cfcf661630f8afe5f70d3f0d291605ccc8b22ea73098bcc1b67ca507acb4363d227694b4a00e869f9aa917de7079805d7dd2327977fcb46ce525ca1a116c07d8717e543cbc6a8cf0bfd3d92e94d52a25232abd11a7d240f0c024590a4342db18bf007890f1bcc1e96ad046639d86383fb3523606b80fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bba2fa023d6e360a695bd60e7953ce9f7f3df94c6d220cf58164785fc4b9799b4f6cd316ceaf3f38abc02dec05771e385b18c2da3ecd185c2fb83ef58df02dad7e463d9906a340bfb661f2e9125c5b3200ece8d2078081f120467bf5a87c156b9710f008ead624d9eebe67a1673c2989fb538c215c3225e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16efc413fec70b902582d89c4252140e9f4ec891136af521a49df2111991389dd366e9194ac14e4afb16be4d4e9d5b06c2533ba1f229c615c94d2d2fc26f0e23e380a30d6738db2b0e15880a229bb8db327693b980418cb744bbd48c427659371015bac72cf8416ab3809ea6c199e62a625953de2c5cb7542;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1efb43de360a153b2e3782e7c5731a0342a33efbf2fd068707a201c0c45dc2c103b3977c097cafd5af2a6b41981e5c10e43a6d9979e3b9a70e55f18fefaddf71cfdf9110114784e251ef706ecff294dbfece9a33762f611ff411f1f7a30eeadca164c4e64ecc503baca763bb03bc94b16ba64eb446ac04438;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1140fb9c972e79558c5202709c076dd4ad923db6bb2e718a79538d1743e6acbec59b70b7bb823194b00662268abb280c188b3ecc5769152d3e74418cd9812f92dd2753945a5313623425d424407c082e806e976cbf56cc7739a83315947c3b4c8c199dfea041c7ead2d475a0fb67c177267f17051ff91a575;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b9c3f3343f4d1c3f90a138cfa2df379e444725e6c877670846466dcb5d4c772db829430c25ab058700a6a147d0b19d198db438ff0c698ce274d07e1b3a906820a51a3260a014b80103b45a691504e7e9cf8b5b00cbb5fd219890fbe0b43260400360c625d89f27b17a2f4453abd8e4e06616c41239e8b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1851b130a2a23feed24048fe55c04bb9cd24d611103ea392da8a7aa96ec0b5f89c607974d0add1967faf84010685e45a8f158feb8dd3da89b3d4ad613cf4e329f69a87daa27b1c9437a2f0ded688a24cc3b622e155d3476082ba7f4b44cc3ea92fb4492698d43c1b3ed2ca076d7ebd15b924bb88764deedd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h502065bb8c3497cded0036855e0770e4c03042a25c28ff87274467926c1fc2484b1a26259cded838e1e0cb842fded839ae65be7dbd79b600e5bc6746dc1f55b1f5740df2b60246cb5549f531a44094f5e04d5890a905f3504e34ff91e422bb01b07c8fef5129431ad0077c8af047df94c6fd7f9cd320aeca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61a504b468b5fbd178f7193aea786c97606d22381dd54ce0e73a4da189556cebbe8efe3f869619d02f38536567f00c6057a2deec0a755555d16f3f735503e2a133fa90c4d351d5e99bfa4138f07f0979d679786c0adb65f89853bd9862541d3aee155aa6622ce0e7038e99d65a779cdba8504e8de2c46559;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a799e215b7a663975ca2e3d138b2bd71b2a1eca2dead284875ebbdf6b9e81c0d12f66bbe859057d28af1e98a38eb5ae7b80582a324502df627238d033db085498903ffea68cb1615c0495fc1d259cab2b7ae190c95d99d648aaf1da8104345f6461920ca9c6ded2f55528581e7fb9cc60562b5097ca72ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f29e3982c3c37dc913a869123e7bc7c49802a4d6202c96755a3537e48045d211aac1076d6fa5cf8aecd5aa23f63f23652e86e2e1d3470d70a89d2629ab89eae3e6d4dbe0f0b72f669e4b89fcdd22920f82cf1bc58b7a1ef29f5954019d1d2d4310c4d9b77b0803b3d795b18ae3417f7460904152311940d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ce6b83c9180112c11ff7619e2833373588858fd345f9498eccaa3139d498c6c34a78ce31544ceee84af37d4bade643a14130af32e91e5615535abad601a07bf1ea23486fa7c01c73d1cac8e08e99d71be0fa95a078d8ed1b6327ddbcb7137fa918b7ee533cd307f795c83dcdfbc0f225383a5f6938316ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b55200af593a438b3ce325b80b8d8378064e5db191c27d234e70e19298d9d8137a8e39a2c19386dc0b27af106b433fddb91e9d213de1ab9fd95fbd6805c2ce1f58a8e0b0b86ee292c039dc81fe9a945d994ec740cc5abd28d91b9bc54d27d039c4fae21658ce968f3651737657792c6555a62482a8d23cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd410c43ca108b88d12f7d22ec70f85a4ac1d003e722821e138c600de606951e39ab8e18f258ccd3f19fbdc0859a05503fe44c865645d4fade887d27bd44556cc641ca898ed8774f6ce01b2ff6094f5a2391dee4c53f3bb240dc3ad24d294b5b1130b96a083b2b50a33d0c171bf33b8af2071e9f06e1e80c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5014ccb1c4d0fb3073c38294dc03936246db914464c3d184ac521741aa8baa0847773a67609d7f36b79b8a1c1980c09cad7b9ee045518685c4d1b76a80f456c54e41398b3913d5be3603f8e3220434002e4a540aae045565cc9336fd9ff181cb65753ab69ddc005280c9dbaa7d641cfd304643fa2c6274ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h92eeba7daf851f91ef138bfc1cd64b0a1f96ba292dad5f3bf224e5dfe0657ddc158c8b0679f15ae7374abb6e723998eab57f4c16f2f6dc173db66ba0bc13c820b27fadb129a5ce6a22a70550200348938694771bcf972606872d44dfe4267990b01b1d6e257473ebbd5a9a916e7d1bcbde260bec756a349f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h55185920c4b16c0165d2bc0be0fb9590ea827a3ee7b79ef88a9691b76816589f1ad334abae3cadb042fdd0a6d5b8f4e21a30c94990181cf23f074248d37b1256cb923252d93b123d90828dc54d2ce23f6a6f20ffd1036c7e377460017f706a7ebf55b5170569e94af2244ffa5176363339e1c0b569b76960;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a9b06048e42f4019c27bdfc2e54110f5a310be399f929cb8ff012b446d9732ea57271b59640cd520cfc820ff975da72e3f76bd4a7ef6f7ff2f92f701e55f1ab87593df19ee077dda4c4753f2e00305e4b7d30c008ea4cde40678b6e6190eb161f2f5c69963919e47597c31148dba1b34222477b4618ff3f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f8c295eec03a829d3e8b7b48d4ebd43ebfcf35995a105854f2df279714fd10ee90501c83f409b5fadf8b25b4b26bce346777c19a3f64e209af5eef4c2c37dee0a331e778c8c87241a57ce8612c29f45041d23f9846f45488279bc5f23a07a8b210a34ebcfbeabe75f2006e57bfe83f79d869102475484f9b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4dffc9171d5de9686b7f9d54dc01a13fdddf607057974c1a67261f486695567209ceea164e7bc03ea359f5ebcb00adb94e5e0ced1a29e2beeb2cd9b3ac6c45f9d927651b5ae4ddce9f6e49762adab4bf6498c013654211198ab7f5e7cd3d75e5dcb41e579faabc422913152fb70377d6bd72d76c37058420;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cbb17da0152b1fee318641647d8a2d7d0141350c5be8967bca90e93301ccbc23e774a27713574d300947d93186349cc074e01c696601abb00273ad7da76b4434b4df927ddb6735e63b30388f6198b168db7102928e9c583b31bfdff7c69e92361d326e7b53a55bb58bc62d42b758765c76bc5d2e10842bdf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc14479fb4a9e2a339954b2407f2d0a51abbdd6823d676c08c909c0eafa6b714489b89b6a2eb4291b0bc43480cde7dc30242fbc6090338c9710d29da600a1a835df0fe7e006c6ac12da71cb84f136ba29fd7d5291257e51d49d920dca3939c1b9c8b601ac2b33e65a4f662e85b397f3aea3fe20007c926c6f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a37ab6e7174d4ab5b15010408bfc1883c88f87bd3588569f1e99edc949c18c72c0015d0b4d66d68b6eaeaa158ab0baa79114976e4f3964505d311805055f22371b710b635ae4f351cb5023d2fcad6a80a2fd22eb69c3a7c7c837fb1637c9af511b5b528747340c78a9df11d6a391ffbfd8528c9a3ba696ef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e36b09e718a48f8c063f4f8c8e5279f4f50ad90356b336a04d1e5fef87aaed6b23fd17d6c31a87dd726e72f9c4714e68dfb0c4d6a0266abc92345404f0f263f4f77e2efb8737f9d4ead2eb8d9c956c861578f15b5fdb88f2ea442d96256c6e2b50081cf1719ccc4395b93c9b8067a8bd00119ce50e7b0e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b72ffeffc29e53d706a3d8d963e1ac8501ed37dbb78bd7f48bd3d940fe2078994f080c852cf2eeb5b4914d2518aa3afb413362de544e1500d34d24fd3edeba3e6031e7be07d53f84eb1b3b8564dfdcca780a54f3adb385e2f8aba66808a2adcf30fd3c79fcf2a7126a54843e1877df3661b5fb7dff26cbd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146f6f54544917f876ce0471be82cf1f656db4a3b5f702325594a6d93aba6e841a211d5653cb671a54c36a08b07e1595f507dd05a31d35e66d091eef31112e1a7d4ad1be3335fd1f07e393fd36101d272d793397f9805d64ed050da4bcecf67d7c6a0ffa515bf0a4e2828fe7ce99b617ac24af10a70a5495b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4daa38678140a29f5c96caf0835cbbf409cb270ef9ed1991380c8832a149491cc9ef08a28d8e27a37dee10a4eb69f7dc5b3e49d3f4aa9c743dfe84766e2ed5d9c4babfc52746883fcc72745cdda49124ad58ecfba8e6bd3faa501efd4c038f557ff2d58f767e7bb7b38ecd9f5b08ba9d2d2608fea85248b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h785b147045284679e8ab640b5706065ceee577913dfb81ad057f0faa0d8fc6ffeb793f93196c14ca5ad10c58e44b81cf4960fb882ab7b018139cf8548d2664fde7637e13c9521c5798b3924398161f2b53db179065c022297521dd1cf51ec50ca9e6e217c2bec53dac60f945a91fc9437ccd212abb1d29f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdbd4b6e5c8cfa0d72edeeb84d3e065eab73bd07bafc9562a81188f5e7c4b94a271870fc0fbe8a7f540b2e3ad1fa7da1ae8930ec31f80aead7d2a1c7503bb31d91f6059a36af8407896ee050e8f0ecd945466641aaaf95ef9c56eceb80831d4eee6f77b38c5118626a06ff24365ca2707b3bdfe7478c54f85;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f2257432c37445959aae8248b8aa9399d2e53532fc18801cfc39bae0418726e124eb678a24d62976b53267cab02c51c9a3741b335052bbc37a01f21f0ac0cb0436824bbe60e6fe4904f6c85eac16b89734017e205d12197d0553441f9e8dbc64406f66dbc17f7272834ab8db99d07b5e5dd53719b3bc237;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4800089cba1d5e50300c456fda7152ba70f7192493b3661c155b12969ca3daed5f674156edc2bfeaa66e932fafac2506e336de82411e4143adf7a59028802bdd6d9ce701f6d2e79a36530e6261b1b93e1874126e180d540cfa3b0aea48ac6f58eba5174e545deb97b9a3f85a7dd9d41d9ee936f6838eff6d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7f87fdff137139812ea21995123113d96b4edb782fb0723eaba8673be57a10af0974c936b2f80e363d553b8a5e7bca584f62e5bcdd87f30a227753a35582e12c056346cd30173147328ed72b38b7dc7409d80e7a4d85b0745685981e1d71d50d846b2e043a72bd78b95edec78b2f6692cfe183d743d4fa1a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14325ddde7b238504d6567cd5334a10673210d580af76b9601be69fe62ad9c13ae816d8c85e4aa1460581f612a4986518060addccfd58f861b9dc5e3cee9911b66f1ae6fa9f10d51dddcd93f48aba50947c653b0518f51845e7ed3dccd093018745db0a402b565eeeca66d78b6068ddfac1e5169381d18598;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb2c7a7fc7be14bc4fccf185653a578fd1ee08d50a6d7517e72fff612e922942b936978cc7c676896415a1cfdd61426f62417f078654d4f90d18be561e184d8f352caef963ab56912ed6062e82568f76b039a3e69f4af6b2be3ecdd50ac80eb584d478bca786d966d2661f8fde1ba8b6a86589e193b411a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1741212ef5f56f149778481fe26796c22dcbfb2b3f3d1329c2d3de7d0cdde856ccdfc284bbc4c56ed582600cbf9f6494550d0f7540987d893b363413463c27afc2fb4cb0e13a79216070cbdb60e941d9600036626071feeb391755025251387b1a181d8748bb4af2a0922be220c2fea4cb9bb4f3ebd983b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8daaf7bdfd5f0e87a2151a1364b9467e3692bd3142ed1ebc57756097f3e9b29daf1f22979f2a634c926ba9e029ef7075b8fba1f68e4191de2fe0ca6c392825c06975d8c946cd4006043cb337d64d06968f9fd53c2fdf463a348794c8effe998d7095a7d55222f442efa49d0ea3fefa6cf254facd02b00252;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h60be700d3b471b06af30cff08d1d501ba815551d9bc0d260e4edf638d72f4daaca71f788f2d640adf97f968ea68efaf144e1eb58aa1efd2ddeff665c4c97ee4872cb7d8db02836429ff8f86aa8ff2a7b2b4de23ade9b402b2430c1e0f3cca74c3ae053cf81ebe70ca52f0245ebf933b35685722c1ad1a707;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcabbee1add4502c2ebaace1c57f956577f5d466d4ebc7efde9109e74ab348de7a9f2e8243314abe41cbbe158db7c6ffad884f7255f63bb886573c5fc98880a096644e5ff5f084ab7e688a4007113797ffee91e934ade5c80ee512045a35e5da1d82c038591a71a8b8683b5583e6d2fdcd60ae7a73bd093d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hadd34082722f564dd3c4bf6df5cdb5ffd158e26d32352def1c7511795cac4d066a81c5c7c4aaec2fd89b87fc7e495669a35364ca7149baa2ec29ae3ff47b1512a9ab82cb1e12044f9f8ec263148f633619e0a3058e90e929a6f011bc55c29024b1c811961f6b4407e7554632b649a1d42e4a68d792b04d11;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102f920f2cbd051cb786e87bc188de54c481c1f0ba450188fbf708782b384aa78bd4f9c79ee5c32c7097a20b7b6f83d1295c8ce20d732eaa7a86d200edfd1e5e2bee062ba9b5b43fa295d24c71f028701b9fa57d45548500ad8ccd16ea004d17b25f5145ce2828bae56eb5c99e2c3f4726d336c9ea4984a85;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11c49ca9e9a98ce82e78181cbf6208e78269c283277871fb2d12f000506562b88b487e6d073ace211e4401f3618ace3e783cf9fe6cb0cdaa0f43cad441e13ce0207d5f7d7d7db7d31b35e97e1a079997b714a1e3295ff84e33bbfbc0e7994d5df3d54a736ed18665e89aae9b7fc5d247c04056344a803fa11;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b2704db8f7744f49df7ae88ea6d5764546fa80f69f0a2ab71794432188c384b9186bb2d04dd9a13b04683068e26749a8c6b244690fa73380a7df0ab37f0679c54e7451db28b45fc281585d87668c0de546bc2aeb4046f950b2126c738ad0f9ea1adbb5e54a8deb151c10edc97ecce94cb755e75a2b38339;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1861b7824f302e9dfdbb87c57b2de49bf0a9ecc0575987b4637d4cb3e3b10db9b59f902596ad28e0e277ea4ded974599ee5679b4a702c16fc20ac6d1916974d6d73cb0168fa8eb5f090211bafe0fbb7cec20128a04862db667c22a00d3093b402d8c5d8837f892d4d6c9ec12e1b1ea39d39320be81404a022;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1949ee33cba5babd280b4b2a3e5ef11b0fd1f97bb1b5a33cbfcb33665660554cfe9d28a425ab4706b10cea025445a250d68fc77da1048a000c9db8e611e4338b7cac044633cb9e593446fc32eeb581b6453829b134f6b1e4d09f7ec8497d97e9d7a14b785c016ba651076adb8fea4558f74b3130a4d541065;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f2c846e4c3db0a020821dc081dfcda4f877039637bb2476557638c829d6f290f520db96b4a5f70b34a9bf54800ec192543cb91a593511ec2b0e684f4f7fcc1a639836de12c37b12e3c006a6764464d1706f7bb651bc0239ea783bf23ddd643fca8aea71b3292dc029d537ae2fe2777b441086e16e6fb13d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10fab2172778763cc98b0f608291073024a8bc56f6a0ce5194e372d334787fa3184aa5c6e4d9a2b2b038f6bfabd084b241c7a32943e5ea7d8f518cd2513808b284406c6e63f5ccd45e181836828cc8cd09eece4698c47db4b214448e27b231ec24e62ce50c7175d02d32abb5c0dfd01f3f1c546d12f038e93;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9fd3808ecc0ac85d3fba0d0fb5f30aa4592dbd6f330b29c55c9cef35b03cecad53850d42b03d23bd6b17a9f1330a6de44cee32c6b4239bb6bde65747aa79b059c6acd63e1d862cd3d50572fbcd697f12c81b9410694efe415484322923024a01a7642430c1a2eb69ef76745ba99dac17e24e19c59e833a87;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7489beb1c449319675b9ada85b562b3fe7c394720d1babf3b229c4a2ae6f59d6de1d1877a23f74b5baf597ea6da75403731a5a96fa8e1cc8f701df04db859f420de339c672ba5b9ae6c9d41012f988d1b88cf47edbb6ca37d1fc5deedb55ea0696eb18e3d173c954acf3ec0c02c9496198e5d9f28a631cd5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4537276a0492f78d99a99aa47389f502bede98d84d58d8c28b2ea58444d60fdab9c4b42f075ea61d0997d6c2f2f9b1e7f04e45620501674b90c1d727e11832808023ffbe117d87cfcce2ea7d63489b6f8fb724836753b1e8d6958e0dd4aa39d293e3ca835095338e098f52ea47134ebff6feb12bb33e4162;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15c8454a41d6133f4866660c41c7d3a06dfcdaacaa23bdeb8be3c8be78f78c7b601c5916448a631e23dffe598e5b770d3fa4e9cd8d30750d8177abd9424e2c2224973fc28b32f66c28424b591d4d4e9223ffdb4e4fde4a4594982d3880a65375ad6fb6cc427178b235436f3962c9fcc3eeb6585668c0f0218;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157b8419ddfa08798f3c2fdf0585606bec4a7d6bb91f997722342cbfc63c8a47478c669a6c9ce3724c99664523446d7594f23d3172e6fa7f6be00bf5e91975e7709fdbf116715e824044e6cfb29c55ab96769bdc3989405028c101ded815807d972a5d38cddb389c572df138d96e70bda328c9e8ef96d8fa3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6dd4bd9142579591385697929327ad2399440ed699f741a35fe931d960836dd0e1cc73c7927dfde01303180fedf60c8f79cb3fd86ee703490bdc2e66d0b14c81b0d01e1b2029754163e8241b89111ae47286c32504429492fd4555e87ef838c257f32922733487ac5b3c7a692a9d13d4060fe11101a80e66;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102459dba0664719f485cbbbadb93aa055dbe0b1dd775f48f278ef441bb9846b4e2da17d9faecc7fb67f122c7c48dff32a2f7a9b9d23ed97443f6ea64e52ca18864bedf55979deb8fb14e9471231b17a8d73d8480e8f515d8ff13737e3880cce727c4dbb3ae4d19f1ea847b714401a3cef54d9455f032c03c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4538092636d441df47e30267ec5afec832a49c8d9dd5b83fd38a617c36decee39b8fc123de87cbf85a0fedd19089d6b02d43d2438f30e2b88a80c40f67319887c4dad9f3017d1cc8bbbfd1d0823720ce2b02a5c4d76fbe23dd3b4c14707f8dbc22f75d02a4d647d73fb9748220f679daa8624e8c3a41712;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h676b7a59d7382ecfd26276921a8ccdbff838de7e70069711e26f3ae34d11368f87fc1830c857086392753019bb1c54b4f2c153ba3c68733d69d74c40aaac957a839220a60775998d49554ce4d7a739cfcf1b132cd4b1e01b31cd7e22c9846d6ac36c141a37246532a2ca41e2a497dd82d62240eea05e3a83;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7f200dd768425f08d1bbdc27c9149b809fd7969b5fd063c653b419a7979159baff6dced829aa150ac65917a76c54f04455f6ccd54855342e937b636d597828bb4011fde2dcb0c0e5a6e678cffbc698df41edb3df46d909cf6f854e7b1a965a351ba0510a5f331391abe2f9a711e645e2bb021ce6b2380b8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h134be57738e61bd3ce8446d8a94cb24f8483073fd70eeee1fb49ad25d1850c163c6d11b1cb55a43cd504dc426e4b27a9d8669e7172c040ad6b5df8c4db79c3b97eeb2c94ef2b588350463b3f7bdd531d8e1166754449fa6b89b4d14690b34dd0bb1ca61955cf9af98dac4601a6be9dbc823a59d3726d5ce46;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbada62e9c53870540a7a090b86ffe5eed681949be95141d0a289a55c7e95b3fd03d67b2746aaca242ea9a2ff8ece09bc54b308a75eb4e294a6fb14dbb320ff1cbf89ddabecf17bcd9cf20e99b9dad31c0b227b2345582c92558e9366e36e000fae4d96a5bd025ffab63d823de57db4a1f59347ab537363f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a3d995aa1d9e6e88ea845c23edf5850429ea1e1c2feb8e4696919375a6cda14565b5daf419afc83a860df7f7c4a4c165cc98ac089ea744dbb685beb33f929f50856494b407a3ef8a67ad54bc1e41a905f381f62a60c08b8ee1fd0ec4b6ad182cc2f0a92562c56ade204aa2069a136fd358cc5462882d68d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8d5da0d91fb255f24d24ca949c5831da7351da3e0d6daedbfc5fdab30306e0fe0e9f593bccdee6c15f79ec68c80bb2dbc4d166b80da026a22d2141f8e71d21c650103fd163722a1f3515b516e2d22a0ebc15e88713f5697b3f1b4e0e06a100aaba1eb704541acefc73fd3d6e7f8bf8969a3b76d6cc46752;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe68c61f5777e9fd53c0521632e9c618e615660480c2d37e5ee12f01234738e838853d551e86dde459003e4c75b4db5bfad8709fca01d23ce0bb7befa1cda98ff9dce7649fe82eb48bd2e6ad3a6663ee45edf9242ac226161ddb3dd400fe36417754cd7bac43175f6a072c1c521b4c2924868ebdd81c969c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0905d3bac3aa582e46b1ec8d35fffd698c352d93b4815bc93b8b8c9bebc252b8b444de16c4be8996d65004edfbee5d12504077a18aadcaa0be14ba58410aa9496bfe1fa9db2cc298fc49f457fb11017724f472aaf6ffb25c25e2ab9e076285cf913eeb8201676355d801bae9250a14887b0dab93817f12e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1780d7ed5f4e4f8be218f7c59a913a0c82de5783321e08203ed35e6022d1dfb3c23be8d0872d53bf1bbda0bf645127bb1529ae5c1b841563b8e74cdd7a6fe4ffb039631e0c04f902e30f4e66bb3bf95a2df7cda0fa66bbb2e5339d3d934699062a683c154bc77a4a04b4f8416974fd824ff06ad25d50c5731;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b95026a40a03d23f90a0e8a0ad8acd38b86c7fa98fea27b045a4a9c203307407652ada2c917c26d56177994482b668a85e24cda91a99fdffde21d83a83d947c7276a30700104731a99d355d0f27993b16c0e8a2bbf01b1cbb59998d8bc39862c25ef8c58ee7d90178019b504b08c063913b1895f8869321;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1210492eb8e98e261a5abf373e1082366e9834b09fe2d761a9bafd9bb0e640494c47a00229d28747ff5a8cce13bdc47a4fe1a2640cfc42634b107ff76ab35d92a1658f0e4e776aff1c481b3883f993576eb4bad0a8f91c0f8ef216157006738969b8290ca7be41df3f16091bda3e767aa3febed7d1a4f92a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e0e81e41b7d82b6c38309f5b8db420302c53af326b990baa0a17acfda8a26e5a62112c1bb35af14d97d1573cefb7029f8ba89a3d71a22b5710475f3b96f0e075f4c1ea0f6d6bb82094d6fb9ad4de589f559b31f3fb7ecca72a9f0015c772ca0d3c74eb40d83671a4c545bfb9b4c56ccc32a94acf458340a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15e47c2f4013e0602dbc362cc92ea5fecea31cabdb133221501c502f969447f36a211af4ad905b8437613a57ff8f7e5dd05f3d153fd6736993952cda541108e07148e15f0974293ef2784050a50dec3987680d1b2925354c092627548f17620b1f7d603e4ed7e5cc465adf809333ba3367fda5da51dce7d3b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h98c49c48348810b6f4f659143eba0f643f113a5a27af2bb8f5e88ea7767bfb41cbb6cc59a90babfcf92110cf21810f3b745b63eebbb88851128da580ef359ce7461eb2e294f446e06c3b9d7eaf6731d26b220ea2d344c71cdb1e32d440c7df520a6de621ab402074e591604a2bdee204d64a288e1f0ab13e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b20ea9150894c007df6fa63baee84d4081210208019e60af5cb326a12873df35d36b2ec31d4a5ed4a20c4919c7159b01b2ae4e5c13c83ccf344302a13a0fd577b88ebd843198cfa6f6d995526ffe302bd95ff9875d7aa863fff8a4bb0e64852b7160201ff4e37273ecbb9418b69ee030cf06fa2b2192dc5f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h51d8b29c53d566f565fc707d40391cd40ec87c9e12ef6be4054d3166dc022757dca8636d965efe33699f9695164b7fb5ca007262085b2b31bde68790854518186fbac33e898dcd6e47a021c6b40631616ec7ee3b1e90d2e36eb731549368ee38e9e343da1631910030afa414cdd7911c418eb61c005f3dfc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee3f0abea865287c2fd0c6ea804847b89585842b1eeb96b2f5e262d71c66a436707952b7fe3358112fa45433555e910bdfae9cf03a86aab944ccb4da41976df1557a528bfae2496bbc23020eb09b561a6f446fdd9723ee7107f2b12ba9e1e8da8595bed05a550aa0b816d4053a8d21503695bd54a12ae6a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4cc862974f8bbd4717af2788e0531f2fb811fb7eb56470e6c79c1033021009a6301b402cbb40cfd1e8a9415734685d1a4975d60f4571ef3a6520bda9c9bd4f5071aefac3b008dbb5f77aa16a6aa6f7590aae0408f0926eb078198c995d8c4972656a5297f01b4c8a7f32e81ac4a28bf2f0baf3a437db1b92;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181b9cac80bb647502ccafaa1408790a6960be3a52c92f6cc35a87a51e78cf651fc452685ac58bb857cf29774256b0adc0cd23198c8439f71fce7e3ab3bdc4266fbc0706e5a931392cc4f4817feab5408fd9891985b542f38857731fd8d0f17659313acbfd7f1759db7c8c2141ead005bb2ad589162ff3bf1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd6552652d77d8e9c7f5b22d66135b13edca9c35a7ec5f67c85262ec346fa5dcf7e792aed0548667ef68129cebf314662c13ed80576cedc8196ae57694f21f41dd033d1f976080f93d2e1abed6ed015883cde06768cb9aa473a3cd29d7b85b7c48a63bef6b3dae9ba0c007a2a311bec572ec69c2f7d5812e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da3ae2fd8acb1bf97f063c4fa0fddd7e9f70101c3e1e57bc3c947ccac1ff6e4f4a56e2b01fee304bd5b460112970f57aa9f7b97f195d8c9394d7fbfe9a02bc4a209211944a10a4a6cf3f10b802f1a5334a923dbf01f0c5f42fef02828cb6e49c54699024f6f9c6a32b6d117227e7df82c11b7f34a1fd1e07;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc8f3ad062cd15676ecd25e03f8ce92d55388b814f348ff3b502783aa383a995f25cdeca78dafe191cd5a71cd1f084dbb9829ee1d3be4394bbd75dbfe83c16891eacfc78833627c2ecc52747002bd14dafffde96d0102a4fbcca6a46d5ca5750f1d1fe224e88a9d1e37e560d1a4094c9aaa47b07477a181b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c618fc562b697754fd5fdd86a84fea7f32cfcdbd440af6c96728dd85217af390bb96073d27970b0258695de5807bb4904a71d7675d1038e9f0bb66c1bac7b5d131fb5013029c81cc50d35e0b5ff191829efced9c4ef7bf54ff44a356d10f1f223043f616b79e33a9baf0a61a6ab64d7a92571e3eb755128;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3b5f2faf8e0a4ace2c38dbda57b29a767e6b4c1261964df60b8fee5eac6f8225e3322e3657215234925e4dfee37ee73532b361bcb4d93a977eb034100a6eeb2917a7e024cc259095ac425f55c9ec83689ca21b6f6b94779c16cccb888461e69799aa6b33cf0ad6a16ce3b7de2831ca1ded87f104c515384d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9b9447f7e13b9956293b21a9e04732b7a7f362efe9431f3bc1a744fc1468e39d832447e8b76cf53d02ea0a6363a6102b2c338aee97e6da1f3861d8a57583e90fd1d3db3551d1eedc98ba7b77864283a9b652a32ec30ff6e8f1d5d8f49a1bbfa31ed69a9be4a7a3fb9d7557ad7d4ba47a8e7d3a28776c210;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h694a572df71e3a8343d1c846a8ec36ec1fdfe69e087cbce01fb044dac9dc3b97fcdafe5fb4baa9a058e180b769e07496746f552c034a9fa271496f1d75d67fdc391c5afb808f38c701c6e31c02941fd661349d5d733726226cd5be92bbdb056fb7a4710e25846a1ebbfb0716c15b5e963336d0814a1a3b50;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b0928ab5dc3e6775c2329f98891f3306ba3b31254159b2871662fcb30c1736e1b47f758d71bf3600f546d250098051fe4888a165ffb9876b0b71fae83cee2e1e88fe2fa6aa05af372b9eeaaca1e655612b5071bbfde47b547d7159d3240a438d86f1ad7079bdc6bcb9249a1692b24ec92279a93158b0e233;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c15828c3973abb3915583ab5efd697b9012db946096c36cfbb2e164f5e333fa6f7d30991a0e3cd93d0643142cc39aff2219d701c42554e5f6be333389da7816d33cf153151e082473f07d38798a54dbd55b7b418fd4a81333edb68ab489d9b2c78a822bb6858d4f373620a79889d3aa51015b2b74e6c853;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h60ddbb99b5c8483ea57299c47e35f763f34cd3f8f0830a0d87ade8e4c04263df756ac7f8c5810ece3b52daf56d730089f336f3dee9e3a6cd3db005925a1c2509b13c5d7353f4c04e65ceb3209392caaf3978d54c23f5a6353fd47b3bce58aef800730c60f259dea17bf3573a6e619e32edcc7944d76622f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1439c4c2b2e7e62bbdf7e50cb4f79d24730b11c27e3001fe79926c36705ea54b1db18f804dc884846190e3c805579a422657554c363dcead20013ae9ee506937ebc24a22ace305534c524fcd3d04bbc0f11c5001e01b65da37b35b3ecf9273c20d3fe6297cff4d000185c57cf2087dc704398d66441a857e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbdb6fd3491f36f9d9798b53942057eaa9400da14aabf1a4cdc54caff6c2cd6e718936ecae7ebcce612209f09021ebfd20c285446cfd51cdf5bfe45488f5befd1d352f6c5b83f52e367d6ab4f9de90c7983cdfc1ab1e572153dcec779920a50ac07ea3a0aff3196fa3870b9a367cc6d267baaccc8c2cb9323;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a17af1bcae716cd3c9283b841b9a63d4d686f05f2eee892825fa0da7edf791b59954bf514623d00db2ded37762e76793decd7c55d2913ab89d99e0c9953df02c89a8c5d1aa3929d0acb8ef726e5e1fe00b24b9f8b0c998b6fe21c950576ea0b5235b97a4c0fd8d54f7e0e127cabfd2b82b3d2284a8d46e8c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h20cce18c66c5e1ef0ff9e5d3c928916b78bdfa0004a6a03cc0ab2eb8ba7cd72543be77d541c90e99d0c7318dc99ad09f29a89711ebaf7021c4c731bb9f0d59dc484f8ca2dcd71709f8584b7d84c31b8f7fbe3c81437575c6ac76cdb06dceb770e2db778a31b4d891e25ebc7381e61cd16ab910ef6bfaf225;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bd1c679287abcf0cff21613665e39dcf44163a0c5c706a6b18ac06e780b84e1dc52317436062e370df7ae95f7a6f1b33f4734193c2419c145cbef87505da21eac62cb8e0735ce396bf978495e4bcdbf56dabca80b5c524b6c91b0e9b34793603a88d9cc2b4a02c2eebd7338cf897e83d329ac09bec3a515;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa232618d6dc67dd7fefacf610d016d446264903e3fdf772c76d44b29f9cdd02a9afdae27289c3a1c2431c8ceca132d8f906df422f3e6b5a8c041b220772002f87990e5eeb6700b0f4a999c8e9f7dbbbe7a367d6a1c42255f0c716ab681ae272f6301e3552fd75efeebb7787f3e24c9c15ae072a79423b11;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a6706744567a16ef2d1fc1187948248b3b31fae876fa69477f6a69c438e7576ed5a6616edf4ac68cd7ddb358d942b877dea4e63323f3b0ffde27a79eb306e3bf78323343cd91017247115352e03d81a39ab493144c2eb1ffc8bda90f04457a1d4f829ba109a5a50c6f417c33fbd5bdd39c657616eb10de4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h839780d56c016a630bf5d872108522422b81f9e3ca98dc81e407de3eb8280f60f9e0391fc03a6671d57dc45a3d9e4eee03bd3dddf0eb907c78b67d10c0d399e59d8e77a03907dc1b4f662ff4e9e7371a29bad3b22c13c699135bb48ca05206fc56952a333123625ac371ad74ebad88de60da769021c2d1a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4c35e5ced229e318b4ae0b07e77720d1c457bd6815a8774018343a7fc331ec52a8ce04ea1083a547e87e8dbe21b47abfa3e6b604c0435d261cd5ae2a66935056ae519f56da742c7e400f61fa89949cf1e60408aab2d1e4cd1484ce49cc939b359c009aa0fefb1691a200a081ab7b2a1888571bc00ce3a68f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h48cd5103454325e82b6fedb65751f1f16a84f2ae44b6109c6cc3d40d4741a6a1f062df97a4b1b8668ca72a598a4f05e7d392687ae0144d5b2a88225023adc1b8fe700f057a19d7ac923ca59f1fde25fbb9ea70ebb3676b6a5f3b7dfbb17709983236869301ea5211dead622bfa5be94cc79cf2c99dbd7f71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac764554b481e101d70c44943c2c8ed540edfada257ec61e02c926cbbc146b31127bdf2f3470f727537182d19f0b51217e981a7b84df9b833c6e315fec028204aa12ded279f2b5ccddbc34ed7319e7d6f323bcde6b385f0e907c6243f330c3f9dd07eba9c9e75f43011cb8a7a0eb33bba75ca12ea16f483;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h122648785c087bb9eeb999714512d7b6831405f403e5aabc51e0ef6c22e75036e97c7eec944751544786a9081078e66695832e16e0fd212012acce10a3e4a16aeeb8b98b1040982ef70a789cde149fba55a2d8c6009b91060d5dd37986390b16bcdda180eef5df52c826d6f24719c8f424d449b461ff868ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f8e42895144f4ff27c5649a6aa931d3c20bafdc872c8c22bc5fc963bb8b0f3548cfa42a42710cb37d75804d7e1fe94b5c6f21f84cd8c89605989125631cef23cacaea25c6192867defc8708df79ae703f140d9dfd0860c5829f4ffe1161b118ecff03516318b475b10ae17f9973461b311ff0a474ac554de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104d1443cc54d873fdf51f29e62e04a996653f77dc2e2a240ce9a4d695e0a7fc684bace8070283c6ceeb9aff73b6a10f082eb57be00321865eef7e114ac1b13c00436358bb215e9f7fe7a22db02aaf5ece6a76a47c98f116f1a5db9247a7f05387bc31eec232ef3927ea5b33b99671083cdb2a3e543d042;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18704c83887509c24c09054fa8fe65f9b2d2121b821c360fda02f80fbeb49f7b72a8297a42f9392285107a1a544200d917dce79d95b9ad60d55a904f347fa015878974934e118ddc9f1830ea29c23465111d39630024554783079dca40add8eb13b30e237f8ecf5cbc9aca84454fa9cba2493e11b1095f132;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb96ee207e2c4e79e80712e1a4db41926e116cc3ceaab689ed5e73f79ed7ddc10bd92e4f08d63ed61c015244eaab40f1e90681f3ac9bb84f7e687d6a073c545f3c7bfa521351cb8f3edf17f569f36dd465d40e7a965217af45e1c89a22e53dd1cfe40802242e7e9af910189bb03de08d39487b10c237a6462;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb3f594b1d266d515320ad3ab1beb11b309ca507eb21c27dbdbb40d0c6d5fbc8a38ae583627485d357de66efabff80fb1e5b56e1a7183a22be9898fa7224f75c92b4b1b7577fda47334edc63caf929c5d245a2c4f89a0f144f539f7c9548d3d7699602f0ebf72f8bd3d7e2e15bef6e4b26e285bc4b5bcb92e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5e238b1730df646f7d2f4cd2f7c0544265beb61a46c124099fd2262057f070084a91e1cd14b5d575c1d302c787fab8f77de69b4957c868759b74f91f719951842a7cdd3b3ec3f695af9312587ec680bd59e26af503907bc7e80c4903bad19a8499a4f177a38ffe4327ba933aae6a143ed45db6f79ca3a16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h221051c9bef80cea2a13c5630f221e31c77ef25e99f8012bb32adebe61ad4f8883eb945eea06f8863be627e7eef3cc010bc32e5609b9552eeec9f51cfeeedcfdb9ef8352c77826c4db5eeb72b0391d9bb97fa2933df634c59b2a06a4d54ac6dbf1da10a16023db5ed7629e5b9290b9417ab50d5c9bd24ef4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47d0dea88d8d89eee7cecfe2f6799b40a32cc633ed937c44e22a7464fec7ca74cc9baabf2b6d4f0e453e2155ad13a7b45c766e6b639a598f783bb8b9b5cb7bdbaabb68f5468cb9efeb10ac4d7baf3bc31aade54c4200fe173487ccffc32c3b639591f7619899a13ea3e7e23b1401a55fe42d3fa17c163157;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5b2b142d6e81deadb60c276700cfdbea347d19f2c75141c5e26ce438c083e075a4cd5a958b4c2af5a8c61ea7c5a86412f7346ca2e7e9d2004067e12f511ccd82713eb3eaf4df99610ab0abe4ecb45229cc308a40e90611c50bbfea6232f6f0c9ce5057fdc0f7f9e76d3a016d26c7dc60b98842d4fbbb69e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dd90c2927735cfc24715428b13be3db196e3f662c06f141e6ba02773cc3b5141e76c7835b8e24c273c2efac6a97e37c164007d9465f2e9a823263e7085b411bb4d62807b04cdaaf3ebdf70a5df4310cca22f2f7a3dc525b2f3e8205a74e3d54e86d575ffe90c2c23817fc357c5ec638c5eee9e6fb8e8a6dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1414169d7a2f05725e4a9a69064fb52bbb7097954810680d4f1f78b945899e05847ffb5345047880894b30040e8abb9ab799267e6fbbd3be12dd59abac228f01b53ae9a619872177b5451077811a3536844dd25af9ae7ad553bc68200e4675ab510251bc6944e6999888d3727225ae19a3aed9072e9cad3ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15897e50a33a52327a639a9c20ef784f799de0b98dd6b298b320469736c9f4e8b2797410fade9f6f5dea9e01a4509696ff24d05a59d19ce561d52615a004ef0b3034f729be4424e08898b7d44fa52f2639c9986362c24022fbcdbbb4b510a926263c6399e46cdf01b1f59bf8f44c187c2de49859b0509ab4c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h195b3a7b5fefae59c49de146acc9052b2dfd660d2d7992e4b58672db1994d0e53ae1488bf8a22b7085d0f2e5d15c9fc9a6652e71c1bb27e3c74b9f56625d3ad41380a8b3d47474f18b83d947c3c4ca2d416ffa881cc9a396c257b0668bb4cc483e40408b021b1e793510d456fe898e0aa7e215061bda652f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ebe0e5035a312adfdb6e201d9ebf2136cec3febc8856442123358c21649c272c72ef95b0899729e61f4249689e95b2dab3f071042bd35a9089d32b193aedc2f1d396540d72224e2c5073e7c91236c485014aaad757acbef775913fa5932ad56df86ec7a15a9492f282dcddbcbd9e48dbbdcab37a9bc8530;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc84b3c3b1695e574ea9edbd4429570884b9377baf1f9d7af3e207a513b59085ea77a426b68433e3ed814de117908bf230111f6c93d38d3626aa7266ceb867d8b6d32efd8e2550c8eab078383bbb897c3c7e4d5e3164dcc9665f122dc898043a2740b2db18b0aea2b0504b169204853c5da312fcb1d50fb12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aafb840fb7133fd1ebb9fccd69a294ceb1f21be6eb74cca26771928a17b27980a46db35ccc9f46fee3b6d10d12a259e4762eb84609e99ea0e63a86d7e85d7ccf33cb0698123d8eb35fbe60235fa7953255fac12e195c8e1794185b5a442bc5d442b54bb1fa8ffbddd101d95bfb9ebbae176b418a782fb82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h197eaee80c4c8326c4fb0a2ba1976aae1e191bdb3fd66ddff2d5fda89bb1dbb316884f2a998f4496c126c61d121d0081113b07e666b3bcf2d5365ace0a5bb78e0f3d4ac23c5fbc241439bfa0978c8f63182ec662e90d61903da867a56171cb71351ca1a68fd4892486147a79abad823d6f24649777bfa2c27;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha6fafd3546c2a45c10f8e00a31623d60dd69667d0721543d7f9a1883012259487cf093a58fb0c7461c947bac93bf4a7af96665fbac1bd7fd6f8138e223f927ba21108bc9025aa5676fa9865bca4efcea11543896df7c45aa1dd93c76614fdf6d9792d92b74c3f7d2273f9ca1262035b03379edc6c56c825;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f58755be2bd78d696753798dbd4c38459069f9893e154369ca4bc6f26cfd985f4be010c8e7cfbf26d6124991f44bf688f50aa5225907c3656c600a2d0d7ca9b8051247b676bb3215a55999461efff439992db71bfe1769c4c1abc65261ebc1f1ddfb761bf635d9cc74e9f3c95659f260a2a1d76efe513491;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15052a46587b27b44473b000259608862f806eb1f14d9909ee520970d2970ee727ee40ebd3d1e1a51d7851d19474d3fccce8bde1a5244c178dad1e36a7920ad1b4c4fe356d3be5888f1b617ea69938820449d48e34fb3218dbdaadcada404b69407ae6d90c9cc1458e1556ca98cf684428f8f888434465658;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c47769c9d78098a24d0753426be2d37e307adbe5d4769cc7e65136ca222a6518b8d628f848ae19236b89cfa1aa1b4cf9f7943995fbc694910b45d4a960a21778d48605a2e1911287c6b58c5ed92dd1d6780902db3b03e5c16a5663f3369ff6dd283c9242b19b64baabcef32c4ba23b5468a427412d14d3ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc6b1170648cda686363318c7d640cae5982abeb4001f13d7224d5cfb363c1c6a081e33e7774b893fb1ccb9e10f9f911d149f47989e799fdfea74c12439270d01efb2309d74e89fd22c85eac8c1f93eb039d5502b644fbd853f4e1fbd5f28c25158625b5698e6474d6c51a401e491164217b800c692fecc1f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb37d63744f6f60ffdcc31d327241d4a3f7594f035e7c9893569de8e10f1ba7422cbd822320d97055b1e83c6329a73017e3cb056cc360466d36537327c1f3578c8dd70b5b39166273ab6f658b3230f0916eb1c04838186c6f736d11fa0405dd1188038b51daa4d5ce88acad09db146629ded8c7853ed604c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0a8c43dbe61a65116728c232619fc3f3ec48a84b61a9a7c4c04aa7acd6410a42720e86549cb6bf9d152ad6c6cee7c170fff0a9d248c2abe61e2e639ee553e2d0884ebf162c9645bb0b913045b2bd7d4067449c8116a9787dc57839327f3001cee9a567a0ecb034f4f824721332af59b33d9a91457dcc1de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b6d0df38b40f2574891e8947fb1181c3e9fd74511a31f597bbb89fbe6226725bac921c81f77cb9fd8e8aa9656e17416634f6b39835c922600df72f130ed8cf4382c9050779e6ce525b390ff89fe1f2a720527841410d84d87e080f7c64d63bcdd5c4f59aa697c6d60bb46c6e586d7564fda0692477677a78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he393db1397d40568cf3e3692aad2e983907798c69398c13b29d10abbffe81902f78f9ddd94ca164f8bc6d61a1f4e6bae10466574127bd32eb52aaadda12476e2869aaa33e151e5d64b72417409b2addf6beb9bf5bb48f98ac122008894433424cc0ae739ddb6ec8fff37dbaf67d6839b44c2aa21650903ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9cc8d970dfe6eade194cb9b6bd66d784087577996d9ae915756a9406a6161f3b0a1f0e40710f268c6cf38a78d90c455103be2f867455fd5c45cbb345660516ce2add9acf0a7ee27d12014e581fe25b3942f67802dd08ea56714b37573236e47c2503db14b1764e5ec57fd7d2a7004ac4fc1454fdc440e4d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1347b1e91eb7819a27e0b9c280fcc38b6d2f53f6dfdfa7157e69cf10a629a92237badaf2bb26aa2e5bd5e4fdd78192bb93beec6d1061563120d5bbf48a9bfe31f040834a00d55fed474f9cc4fcbde50c126a310a0133f056a30bc56d0943d07ede2f0e21a4a2070ac15816350b59cea3c6ff3fbcd21c46c51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13fb8bfedfd5b509db039a2e09355553c33fc9e16c6c2a759662c4b87bd5af1108e7e4343bd7874b15531003b7c2582093b138bfe65d54794f81ea3a089eb2ff9ea6513cc20cfa91e05c6d3c3669ef3bdf401df8b6a28be5458458263ced0de07dae5ac486efcdb1e72934b3048bef89032d5324cd2c8588;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h81ba3200d6606662c4d1c8e0dd06ba7d622f1e76d3432532ff67401f8182ff74b35b7237de8aa0c99af072346d8ac68dddeb2a5fb0b83235df42c4219d85b6573257d5843cd7ef9fcd45979042edafbc27c505f6fdc8edd9649d1e9915c2320797eb2fea4ffc5d69402564d67c3309785633569b5b758400;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h127cbcb16ef002fcfd69d015507fc0b6c2bbea28741b6150c141575ef79befa3445d064eb7ad3508affd12cf53c8698f0b197b48662aa63890aca3e69b6b5691377397319153e514bb8d78a11f2dd4e8abc09880635db5e81f7eb48c1a40ca0f6b63f8488396f0a93d8f22794be5723422814216165f5ea51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h185892d64394d45f6a607cdf925bbc141e5dc747280be72dc3b200cbe08295965159e04a0639857ebbe36c7d34c3651be277a541c95dc52dec5bcc90b157079f5e42e2deb786287f779108f7157fe26b804f044b90e011bf17bc6a82ae63b0a940fff2beb382ebd016718da2f9aee9d967efbfba3e1d2cec3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h499ed8d7803cce6be3681a4dbaec6f0355270f393732f911657c7d5b486d089c970d0d7cc53e94e776b0535171528a918fb5407e05521f53415145bb838d931210515dff12dbbb3913fb3410943dd2b770903b4ba40f7f3764de0df818f0b3a8d164adc89d53ed95dc4008e83763ef9410e0b938f3b72d3c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f74430e647f0e5d353a37c5d3a66e1ca78af56f6ca7578049a7af86137b53883ff2750a294ffca69a7cad401798d1460be2f79a1d97e5d1ea966bbd1fe508bb83ad9a64fe3f88bcde349e7f13c36b045ead82e73f12863ebd3b0e57f9291fdf139550035d58190d921d51f14c436d712ca1a1a1223b7f1a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h543153163a96452d588edc34380b78a5b11b2f9400a550a98ac58c024fb6beb57325b41349a9de1bc4e148ae00b36d5b7c5cf91f5514ec53302bde9969076786c7335ededbb64eff896759e8c671463a274843aec98a2830b7c43668ebe5095b02195491636ecbc5526139028b679257aef6450796db5b6b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aabb4f7e776ba92471027d5c82812fcdb66ddd71d33fe9cb8506e7d8484b5a4a3579ea44134dd1ce627797efbc942eb2d177ac61ffc7206e187ae638cf3e7fc1efae62c4f9e15d0dc8de2f91b8ba0cd9f783678a93b8854908b11acdfeeae7d10eec68df7ec8f5f584e49e45b5b138e51e5e6e31cfc60daa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfde170cc983b28d45c7f7c7ff24fe7bdcf3c16de2f416acbdcefb6fdbb48887bbdde0032564d8202c03d335a6eca3c22d9ca5d3afd3de3cb31088fc4c6b8da5eb75b5f752a9a01f15a7e41d564c61732dcfd04e5d16ceeae84b98c2c6c7b6a13864f66bf7eb517fc6d4a74719ed05994ad2cfb9d1c0d818b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dee04664dee407c0254b2f74f6eae72c3b963c29b908e1201cd7ae9e32598ee2ec2563f12279d4aacc606c9e5a2405bf8563a31357e210db992b2c1141fba08d48a1fd7996c3da95cb0757d886c30042f4bcc3b55879a3f893c399de6769c92e71c159a41a020540a0d93516b319eda1aa90be447fb25321;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115b4827ed5e28c4c986d7c4a25cb9361d03451f3a01b3a37decf90b746508dd4c50684f56f0c84ffedc2e91b9831090f901722e047a91af261b71c5259710869fff00bf40315e131da502bccab74720f4e39814290d151fd1cedb96f56da2c3a3c9f6aabddb07f8253f3d8ce5f66f74ec9eee4da482f85fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132c2eb0835fec22ffd91b1dc91471daaa0fc8b730f04dc1252a1284c21dd00a370eed808b588b2ca1c78b4078635bdf7f6148198c704fa3753ee022651ce36df40061cab80a60565ae734289fcd9fa8f78df246d3bf57a8509c70135774cedef89f931f28eee75e3d4d74b7fd0076a3f092f2a6318273432;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82abb18c3d8c199ecd43277d3e94937f20559beb068a7e6fa07d76aad1a686ab6127ce17b3afad71d178da19a0e7d9617b3cbe99d02143033c65a1497b17255b3256be674b8a9aabcf2683e00f581289968a2b26b2f9dc63e864ab296ebbd4e958f9bd14e066fb4fcd4f09f8d90dd25ac72fa1e17b370759;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5e35a7ab056f23572fbfe6c3d41e3b0473435dd151554743bdde135abbf11a665b9c7c9bedb13052101a584516325e84e514f858a00625fedcade409615296587bc173f65438d48f1e20e6b31de268f1c575964cac424a8611db87606f162592d9870eae6e48b09f4b08ccfba5a6251128debf93224d953;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb7351c6e5b2920ff828d75f56209ae608c8411d7d7de8c8db163267bf8ea25a22809a6275c844573b42ad1b66681ea90c06fb07386b75dcd618ce5b8fce55aed3717009ea0294d079bb3204ae9c92b54ea21e2d451a8634a8b10db208aa312c56e4e8983b3d3d60bb898e5fabf88f4f6a334fbd8e52d74de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd29eb363f295721b29e43e8e07f270cf6692e03d0345830dd5d045e41d60004acfe95cc89144602a16eee1437e72c274fa599bde26a9ffa6bf37ace61b324cced68338a13739e9af8eb8c82a6dfff18c0bd3e0c74144d2abbc25776060d4b47bf415e784c1fe68b72adf8ca553bfb725ad77f31edaa52b59;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h162c812fba1ee82bc2ae44e5e056eca0a218ffea76485744344b5be36efc274812a3bde06900508b1be969ccd3d1eacbd3ecf2f521001c81f9895a360ff826a1a5e052e617705152030fa94bf6879e4ca16f7a2d79aa49f1efb63345ffcaddf0b5dadaf1a20a221770883045d0bea0ac9eec098b96a39d0a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ea6d136827b8cafc1c76503852e2f72f3752cbd81afe351b9a0fa871495d4764625bba4e239b36e44f45cea579c2139ef0f8bc223464e4187827fc18ca7d6a067441b9dc8bb155db229eb87ebba06b374c116643db7bb6d8ac19ebcdb28a40e9937f4715a18e32d7ab708d7a86b59d768cc03ec11d980222;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2197ca5ca93800648b1b92613646bb1eb0741eef6d554d4157f7a52404db703bf6cba08c0e7db37dc277cf0cbe94caaace40f34957cb03982469b916179d8dd966f8d236c506de677ab05eebd62fbc9896dcab1598a24f9ddeb8a1f398926b7ceaf99426ad559e4805cec0604a70340debb11c2e63400123;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8112afaccffe0a3350c944c2be50a440a09ff342d8038169363be3b9880c7b1795b84aaeffd35b122fbab841903de72e7e5b620262c237dd87bdc12d31847f923fc0c42d8f7806c2af0fb72732680c9b3edf182a98efa770122e57c285ebff144903c3b1ef6a741ae451d8799718cf3547355b31368746ef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13010e342de7883ce59b55ee965319c0e9737f539c7894dfa1c21cbda7c14682580a8fe41edcf61d6576425076823e4c2ee7beaf1dfafa488967724c9cc86314f817ed8b9b41ade5c2c2fd53dda55fa2cfb1801e9c582142be79b1defd23078fdd60141904893a7b4cc71ea38967548b28459383f15c3e288;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d2ee3d6e460198727e413efbfda6fd8a4202b9796928781b13c381e7608ad22fb02f44ae6bb4fc0f7e88b26c02ffffc8769114ffc6b472afa1a37f36062db130023e0986f29bce8c4f46707c26b5940d69b28fa2a69ced1d3aa3844960522ae83e46a54e84e3d73d2ccb4c9f4ca537ca83a0d9a678929753;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d626e17ef1fe7b277573c7a0b4a119c1c3e57845344be60bf9d99cf7cb757c726663c4806e52845b26882288b9bf02d9f0d1f59ffa52e36f2e478953041614e235f0116a8ee29f09dd72efbd1a39661887546e50883c5f3f16df918fda62fcc1afbad54154503e3a88cd83310bf3e4a66c9da400eeb15831;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h83c4cba963907e54cdc6dc47d2a89bf8021a02bf0c4f55aebebbf9ec84dfad655643e9e8953eebb43840d3d8e08047ba620671c366f88b67798d30ac8065f431b0d466c462f62f07e06f9ff874721fa00ccc1fee209cad665889277ff481282ede97658bb7ea5a78d6e89fd88686542c7ccb227b2e93a51f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7177b94db323e68d15676fe9cc87dcd90a85edbce101ba8d520fe985be113f37183d9906d8b6deebcbf9ffc441c4c621e18462dd8a097e8220e67defdb4dede972f4a437eb48f79dea226f8aab75a7f19b8931b10ebc990157ae0837e4c52d56955de6166f853cec75d5bd6428e4f141b7d1802823675964;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9bb576cfc6df0af8113c5ddc27889ee7d548b616fdc09f9cd2e3914d95ac65b53f8d748f713a07e80e39323fbc506abf702ff0e83e43982a0fb0dbc660064e3c67dff0ee80d3be691c9e8fd0fadf347ee70e6875dd5787c09929065510d47849b88472b921d76c859353d9678630a1168e39acbdf33b37d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b90e1425c8561ac6e0b25471837caee959e08686cba2b50072fb9deaba7dce9f3ca3decbd55d60048576108b8c7a562397f4386a809232c1460632ed86d4ae4ad9469ea99113d10650fb4ee37f8e4063a4a48fbb402eba828fb82dd980d1b8525e6912312c1eca64f06c972bf424158c1e7ad586166ea5e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haee1c8326a3ef6307c3824f25db723ca16a21385bb064ec1525e0877b97ccf28a9444284b26f2d9b234658cad082448c49d34752459531caff50f4f3e6b9f3bcd5a1ae6c678376eb4a8839e043cd2f23cbd2da09183b6641c776f42ce0726b16c2ecb8a2ad58fb946c44d166e73f83970fcead61d44d69a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heec047866f74ddc162744e1190f6a75e16184c4ad8fede08ad0c869d6b32d231f9b2ce35f534cdf84e7dac1049d38d9794138e56159bdc25bbcee14cd196bdad1a90e3b0a24d2de961c1a3d18ddce11ac5ff043297ece6dfe291db83d1dc6057496deb5487c5da35ab4e48d54645e4c61316610a0c1d28c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h161e1695ac458eb6836c69f41c42002fa78ec35e2c3dc8591ab91f3c6d5516ae7e7db78109b46c8c647d2507ad93d3b3950f9f6d0f634a9250f2a1d18ec50c5cffae2bd004b1e61660cce9ed81473bd7878f8859a29e200c05b2e2a379f22e4cce97173e8154ea963a4fd675b7026a94f29ba4f5bd1863f16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dbeb557befc44b48a8d4514a9398c1b973b7dd7a9ba28d528924514e3a43730a5bac12dc06d4de147bb3fbf2f22b2661f26e854959dad25384ed489712137004a8113ce97c69f9a52b1aee2d389bf42528664c679da9b161789c09599d6e1d5bc7457938ef9e9db98e0ec0ee19cf0b51283d095a408c9471;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bdb6ed57aa0b5a1d8e9e19c4c0c3c276784aa6a5788f83c4b5f5126b084440f5385beab1df199961716a909f16126528eff4e6bb4c99d0966f15bef1912fc35b1478257530e0c037f648242c96871e17455d2a31ca12b6ea2e1c48d563b9d1219d92a34cd34995b1f0c73425676ba2d2e4518f8045356136;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104cadb643091c988d75c566b9c73b0a625c1b61e872b380bb8c2f5dffac38034ad72f57b5908dc8a8f08f8385ae4ff665aa1ab55ba1fdf1c582796a892547b64da614b15ad596acb27eff9c9dd01b6a784e65e356328eb23d051b2c607f1631fe80f50ea49523fbf5635362d2f10fb81b872f87ab2a8804d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1139bba70e4cf09e6cae3f968b2499bcb718957dcfeeda2e526caf97215aad042438d6492c26141c9055fc6de98f4959251c6db2a4dbd03324dd210b71d5414e5b6f704d37369ca0c7a94d832ab8c0ffb1cba8456bd0d1ece0888021e6f8db6cc751aa405b1d8ffc1d262b8851a31fadb30c91a34ce2eec7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h187c77b54ee1ca33ec3f19eedcf3c0bde31947bf87cb01a00efa6b57668551db72a6e486829c980ac07bab2ed5b28c14a1489712d67e5e90e0215f3f03c29f0118f4b07986e22bbaea9b06b5130f344e07d66616b2479ca084cd938ce52c2227ebe6ab14387d7dbcfeeb29ec20642e295dcc0a862afd24335;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc16afa291900e57d510b9776251a7fa48038c252528571b62b0baeaf1d2b2e35c14f8aa3651b319dd001c91a93cbebe8dcc44c53877269835be759d863f8fb1bc413bd41cedb67cc7e95696f7aa396f231a53bd8dc3864d48b4775c1ab40e4fbf787ee1b7f2ad1da2516a4758cc5f0e1ae9048ecbf20017e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa2938b9c4dab49c943bcfce2004c5e938a741bb627ec477e8c4c934f49dcee8211b62a234201b829b5cbd9e5168c455b7c0681286025314466fdb25761ef4f7eccb674e352f0b9209beef9ea34bc753d9ccbf49092047efc2957bce791ef8f5d4a7f172fdf444a96f6d49c41caeb4dc285107eeae894b88;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd6c10a6371bb118d73c7507f6a3becfec881824b32ebd5a15df1a6d9a836b730b8961aed3f4c0014d04c9c535b080622acb6befa17d5f9a35d40800d15d3bac5fbe4371156031bea4c4092e03bd6973b948f8d8123f4dc41ef1888b391fc42f8ebf3a33596d0a730caf2080add5620e466756699f9c12713;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1dc82488963d712b56eb9eb3cd0dd983b17d9005b807634e8d0efad61087b54a3a1de18924cf0cad0daa4be2faa5a8dc8e2e9c0129ac7b5b45787d666cdc266e2b25a7008a030d027b680d855f6cc10fbff00a94cd01841860581f992ff1a5a888d5790008e9d2c8af1bc4a5b762423791558d6a1b7d770;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1484b87b82eea4ac1d0a5e38471683a07824bafbd6bb08b87b7b42fdfe13d6107727f5170a2578e786e58eba5b95365729a3b2273ca907cd6097f0918331c3a553b46c43c4dbbc0ec0c9d2794179b69ac08a0efbb5c84ac8dbbcf4083d13ada57c3fdd9de462f32680c4c126c3a0590e40a8604e54f8049d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de11b9569c9388ef634cb85ca41da75bd9531b99bcebcc443d52dea95582fc8454cd46ca94fd6ded132ccbfa24d6ed6d703f80d5ec54fa2030011e59f6fcbae1a5699d4f1e2930b2917b04888451e3f96394a598ea6da20fbabc9ebe58660fbe428bcd7f224b41fe9d0f6a82ff56dcd12219f826226681de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f7eb1dd37b972815740dd63ab03b1ef7eb6523dd9ff8d4d0605380ace3700d34609c18d26ac029eae7d0193cd2b7b584422595f15aea156563991b256f9efbbf6d047155fb2649ca89922bc3016c915649f9a6f32e7bfb3521f381bde10f3134bdaec44a5b372ee89b951e4555ccbec94627f25b99490b57;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6879a7c572674e43a96583dd09de35b55cdb782665ffaf2d959814dad88918cc0960affe10b1c453c87f1d1e6be9920bdf2696854503c140a99b5a7a6017f538306730eb2018eec624b3688d48f5f3236256f3605fec605ff68893cc930985172e4fdf6d06b5cf0dafa42b5fd51593abe29b00093cb1781;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h87d0e98fc9a407c1c3627fb3141bdcb2da25d69fc748efb05d6af8119c01188aff9ec5ddfe091d46d298e9c7d03cde105fb5e2d0fbc087053e0dbf315965ad2df00569594a68bf6602507792b54d4bd7eee36c9184fa4f8952790a19fd88eb0152fb9ddc4c7301789e7f76e715ec70a8765543027b58e012;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba7b80d4c44d16ac032898a0f394dc0a8cc2daa46930038c7a432621f153e1dd5af7f26fc44c96020f5bb3ff49e31f8c12738c52e04fd321370420842c916fd280dbd4258829fa0a47fd78840ded96955f13730c315b7aab5f13bc852639c45d57c8adde596bf257a6d434ae21bef73f404e75475bf78c93;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd92e2f8379118b777cfe042f283667d6bd3dbb90126dad6576c3185cc80dd44f6f68d0f93b117bfebdb0a6781663fc0c9a0f03fde16f3bfb6db8b0dd9e577387d255a8b02fc4914e39d6d6a17eeddd7b0b602991bb1a893cf67ecaf146d84b09c937b5b47ff221426d1c9dcfb38bc340d33aa7bb94114b0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10a1d0763d837665afd12a1af932534ddc827e0a2bc917e56d17fc259ed20535d35c13bfb2115f106b1b5aae681b8cd4f5209d550448c7fccd818769c470b32a209bec0739406528d336437177436661dea2b0ae61ba0e9c8bce2de3eca2a0410d65b196fd0a7844609a9ac865ca2637da78658267f362e6f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14fb9d67ea5b89ec1db80880e54bd0550d05a21494524040deacb36a51b50d22a8f293e8f20273068bbc4577a7a7db938492579d7f749ef19ee90acd750a777b792e7d37b042e95a362d09139ee36d95289961d1ba88f03e2d4852d07aafb1f751dc0f9108b80f4aacc72f8a43f9b84e113e03782697438d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18c316fc595cf194c7acedc1d80e414672d4d72c4f3ef08e7119cc7097f87533d52c407aa2c68156ca01f52e6c319c5f11c3d8a8bc7da189332e6bd3bd8b8cac27b2a6ad0021347da3ff1edbf248132ee7a5a2a2b1985b4fec7f16ce01739c7bf72b042eec2a4baa3e6f9700037b5c253dde5572bb7275c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106e40c2693a7eb6cf461cc3008c4b964698f234511377a40755f718b58a7ce28d189c4e4fdee4c45fdb322daa1be29b28a3a7c2f886a504d87d70e223da625dd23f2845e88c279e725fed1a5e55b51d772a683c718758ec372c1eca6da6e41f401045831b2efc0364e58e09f220c941662979bc999637a03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf3a301301206531e43afb4f820164989734c14d52eaade4f72a8cde6a3b9e30d374d012867292d0fa19cbd1468bd6670e289ef64af1fb86fd73d46f14ef144219e3572cc854a01c062f967f25fe52df7c9c063cd456502a0581673386de6159846570e85a71d688a29c762de311bf787f193fdd3edfc38e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a431b46c59391e73a8dc9efe1de1b822c53dfc21df24269167232f0144a0322cf644a6025ab5c5cad0b6113ba270bd978f86ad0ba6d3896448df7dfc2d4fac11bcaf8f93d5dcb6060c80b09b38f0245ef29079a86decf8fb6a1dc3bf7300baacafddb924886db1e86a098228ff69bd9a81b6c91cfd910068;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4199a7cdd22b5c2bc30ef4e3ff101c59aa3a4f69a9b8d837f689c809484eb4742ac246c2c5556eb89e1e7c13fe9892a0a1b1f68c4e817b3b5b5f69ce6d099934e94e6c1e2123066046ba6b94b60d7eaee3dcbb07478072955e0e0915599e170d30a7e68e8bdc682d26223e960385993e682d1ca5e776bd8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1784f49f424fe4d376f16a692ba6d58d9b866c3fa93aaefb6cc22dd794c62e179d4ddccb9d303b2610541fc633cf52c6d18b27bd5961afced61635f749928dae3aad53f3dcc4da9695938282f7c1bff5437a0c04713175523ad2bbe152cf71b3081a99b69a60158a8fca503b5de7c3f8c3eca6fe7c569b3ed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc0c5a3993505803b59001058710303dd8c48282edcfab991f864f82bcd11734de516db795e03cea1e1b229e0ba07a38871697acbdc7ae955b5fc779a658e191ddcc83ed0e80604de572216cd447c4ce0d568e830aab8161114460b32a3129612e77007ae5c0ab0411393347854caa2ff41c213bca963a435;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha66b6df90986713a66cd73ec7620e92d45c735c53a760a6e9936a602b47c330df51aca2a24008ea5b4d2dcb14cbd28888f7d568cd1873edbaabe9eb2f9536db397e5a0cab2c9aefb3f08dd33b220de4e1af13125f0ae3d7a991e6b0175e088441afc02856e607c7d891ca8343ec75a204d6eb6f199c1317c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5a9afd993f117eaa2be3ab8b9754b350638cbd57304c92188260774f31783435cd76ffef05d2f88d4bd60974a0792fafde82c1f9cc4929aed415947346d54d6128075371fe93f11a9d0e1227a996bacea45a94ad1025ee93b62ae9ebc9a83f513abeec8c6e719cae53e07fe0c6d2c7ee59d7ab524d19a6e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15fd760ed7bc313ab19effe92106cae78ad2897f0ce7abdf285e33e2f9356b9b678ca0e753ad28b33d033e8949168f80ca975358d90227e016283a99137501b496db3ef91958c1c8caaf9c235bfeeeefc64b803c365cccd89aeaed26a09bd05cf03d9700fea7fc5141bded1d558f0b6ed12f3346c20a18871;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h457292e604328d9eb72c0f44ab8776725de05a99f9fdae7e84b8f0ed4997f01b383105350f4e61deebff23b8336532d38557c86e4333444ec6e95bc93d6b784a65145359a504c45678a0951091177180b80f55638816f7b6efea1331235bd8cb17055fdbebbba2957f30dedc09d1e11661aec5e41459c65b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hca62c45edb8143edce2b4c6c24897542120174af5e760e330796e394ab73320899c09b1efcf59497707daca91873944665a5dd12f5b88fcdd7d963fd5679da07b915defecb7256eb184aeb44ccc7401170f8627eca870e9b945678dcb4597d8d4614afb9224d8df61d4008c695d3bde2860fdaedf3ee421e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h188291704ddf7c869f47b75d906e1c2917fac2a03daea9095c609e465fd797bb08338a4c2b564881cf62682be36a98533874b809202292738b9bb7351d384191414f05f2211febc6cbde77d427447de9117b3cd4269b9393d57361d334ae5a4738e16736305ecb5bbbc7befa03a5fc959b2d41c1c7e53a05a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9fe0ceabd94a744f654a8441d4b91265a107bea84d8c0a3e971c6f069468e4f2b76a0ff7d93bd3aa26d46d0675e20125889c91eab6a6e37996620f49de05414a715d9b38f0d069a06187600c06b4e80f8ac5f991ac57d5330c6436642975916e7b8266e9e674414af02a2e6b66de64542614fbbdf036ef6c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf11e76e89f01038080d0e905dcd37b9d1d73d24b16ce25702437eec75084689402e40e2935c483154e31a204ae03872a8276fad0e76c11336491ccc653b356e4403c42cfcba6243e037d12324793b5fb89f763a3dba52c6350c7e3b900cafc2e04795ce221439bdee719bda91986e99134adebdde5c01e86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17beabf6c4ed3b0e16ae95a830dd9f247ccdc79977acf0d389c028f004bfbfab13a197766f513a108a839eba9df580b19d638aa469fa3d3b78eb40ce17da134c6c87b40239056e46762448b38df3b3cab38e0e93aee5da436d630cfe931c33a1ef2119599c9267c425486a83fe08c956d75c18a4255704be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50656f6dc1c964b12222f5d2b57f595f5f7d6803f43b37db2bfe09404927fb52dd36e9e458ab9dc95685442d6c92d130706634dbd0fc063420f9afd1d7ebf8a6eb6b5b84e218735051b0208256583c6fae17c9449ebe002fc1fc518e7282836e80a674c3dc9079b172246292fe176e78f1169c38d123a5bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5751592757250c0ba6e3bc073111db94395843f71fd89eae4efde5df0aa9914432a0cba6f5e3bced184351d9ad4d0c31d0c4771beb940ca30ba045d21ca8898e23c161f5b7c998bfc1376c782d1a64a6dcc242b11fae659c12335d7c147e0a7f5461620ab84efb24c75d59707e3cb66dcf71d598087c94ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h23b1f9d3b09dd273d308b4c9c0c037757a2d0d42b3d2d1631ea4abb1d308f637883dabb551b5feefba08efe355dc1727960423264f03518709fb73a3d9785c7aba30258c7d4fb00c9470e629161ae624e198bd67d4c2524e519e09c562e2d7c8dd3678a22cf470ca5dc8077cf9fc4573c8c30282619d1efe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13cfe7ccd41a2d2c708e763d7d01f632202a57dd7ad9556ca21f1b1ca7198f3e9e8df55032040a73e11c81cb8dd2e8d56848a7628b056226f8e9a09f6b6235a4d25ee23ca7737d6075c95cb9a9896669e73ab13b53b8c7ac8943d6503f6554d9d24d09b669cd78a96dc3369069f98b1049a5ba4f9f131e236;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d2b7baa8a39471ba84a6df0b9773521e30de5316f63a4bc1bce32070d6d45f1a5d596a38a2836f011c805e1bd0b78ee1cfa1160f0d814963b93f0163acc9c84b679bd03f67f60f86ba89cb97453d6d9b366851bcbab6ed568d48300cedab0d0d620276f42a64515e5cc537f60694d721a4501b4f3d2b2bb6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1401891972ddb2b49977db49e3c33525d43cfc114d6856218aa9baf01ae434d14a5e6ad5867a3a499b5686d761e57a786fea36d53c6a12afae18ed6ccacee080c09c2884060f5169c8f87b01afc59ca63f94b308d6abf34bade723ae7202789b14404c2a8b79038315995a07fecf8bf3969341e98d6bb62d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13627ff516007a8b5cf3e1b19611ccfa1a63b0d5ee26311741f670f5c84164af40b857663aaa9fb565c3c45ca920065934caa4d67b9774d6e01235ae38e725eb779c6e03afa041d07d5aef48d615e882af7e148c1d142d2aa3fdc006190e0f5379789e9e4a5caeb3cd4d496af5987618ddb1a3cd8f141e95d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84a9b783b75b164b210b2acb7fb8f5bf06c4a42026c14e1f855a9d801486c778e23c1cddfb427d3088780667aac5efc0f619e63e4f80dd2f24facc3771364e6473d06c8bd5c088ab607fafc056199db10f8683aab1bbd4b1c7da2aec6ed510beff6f516af738383304ff2a1bab4498c46044ec4bbe041be2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h92e60c310c7842a2992d2f1678f25418d124920dfbeb5c08b10cf793c5fb3cb8eb4d42e84db5b76fa6a84e8030dcef23d238ca336e1796fc41f323f9e1588a704e88f09b40a1705fcd5dbde823000c324bec52333792d69cea78e30015ded9ba235a8e241f3e715f4ea688e2919d9f0c36d73019d6931ef1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h64d4f1e79dd3d3c58a33bf223bb5494c223fc10034ffc9a1b4cad5b3d7758618df2a077eb70062e5acc16260d9313388e245b05978ae6d3c440282675c18c916fcc8de59014705ab4bd948e9d8a769e7a4fba300950aa98318ef7948395056d4c97332434d534763345e9d8969ff53f947ebb5cfce82715a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9591029388de0d61e1cef6f7cad38ec8f1c1c89fe2bd1a93bde5f3e3a1e22d24602f5dab8f44070df6afb86948a036f6da8a2c705a3c5aef20276da5e4d5cd35fa64ef22c6729a3873e0bba2e0d0f3cd93cf64dc101987a4aea6693a8ee84e316ee4da1905ff98226e3ff151baeb01bd89dea1a74066541;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b09e0ab8180fcefdfdb273bb337e86b29a930d3a9f3ebd5003b2ffb55dbce666a88d0137d82b28d51defe6bb0350b7590534fe1fe1b132ab968af13c5025ac1113f42ff05aea9e2dd3cea72a9f68633a4f1f438de3f1f6b8819bac0200debbae2b264ba8120fef836a807d270e2df0c70465d314d293c49;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1044ced10e8116245b6d9237e1b6cf95e4247e87c78aef3c23778885c89b2922e24f3030a64e26323290f0f424213354450617b8145de314b5805c739bfce4521ee08c5bc3bc784915ce0027606c15fac95e9e52eddb9399a03c133bd838790981d7a6109f374df80a9ca5f982ff1e6f253565cd560ffa5f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18feb8775d21a192bbc9a8f776f9d3235371e3a94dd810796a7f25dd5b59787250e07118b57ba871b9d83959893350e69fe2eb44526b73a98c2464c7d3a8702259f8e5e270f26b3588fddb1137189b84cae8f04b4a7f904c5ead2a62eedb6abcced25d53a1d75ebbfacd7aa8c977db599fde9f2415a5e9a39;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186896ac949f72ea7683968438485ebaa94a222109f9a2f576c8605da1dc740c7ae25bce926285fcb860154cd6ee581a7f358a76df2d2fc0432e3c941e3ddc5559e5aca44ecb0acf87566ee89357b5f1221f02697425edd000bfc05145677c4d83f61939e6df8f4b914e8ea6641ffea916dffe0e0d9de7336;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb71c64cda924c341a9c9e07ed1a03a051822d454675a96106a2f4829c2b29c13e837b511773d771a34508390c487ad00771df60ef611acaea89d01221579b087a492dd6c5f0df92366a6c017806e6d0ccbdaefa685380e755c6feb3f53893c66709c7951b4221b61bbae31f9838f2922aa241f67272c0ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f8c426555f6467be6f38a4e90b0c4bc0ba7be9197533d79c3de8663495e6250a284719efa7fcf294d36479d062579e434f7686009858c498210c5a2fc2ceedfb3cb2ba40ea853b5c6f94a79025da29ea88fbbb9ec7c1bd99a065fe9000b4803a4a1a7b77190dee204c59d45584bd616d60ca32779386b29;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90ab04fa4d2d0206b54692f5526fb831915470a52b15714d986003faa680efdec62030eb080b46a319898451cfe104231bdda60bff9c9e8c86a8e76b2084856de63966d312fbf8476404ba0bb6dd799d92c7d91af05b32c6b0851ddb02709bd9cb761b60daaab4ba655e69c6e9c4dfbeaf0b7ff1581edf1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h122f334ceba9700f7a2306a720e5d9d701d4dc17ca82539cdc5b4efd11557ad84d052e1cb49eed749fc68d108fda65cafbad3ea29ed86fa3efd8ff746d5e52f69e800a030c615dea0458d2a1a9236a0e5561c3307388c395cc47c752de326d8a0356fd17d2385cd656abe5f8d159ecb7c482d815834d30d02;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50a2f63b272464880be356c0292d3aad5bda1b0697ef404850b2bbf8beab0c37e8e95188a300955eff608459383812af730cd064fb97b6be224d3e1982fe49dbec0e61f1636c740a884c7249e0ee66233cf7a2b12b4f14036367bfb377cfe8af607bf11e61eacd9319993ed0302e5480156efc4937f04a4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13bf5166b8d2521fd52555d9852ec9151d155939840ed7268c113213b016dfdcd570a6610876bcb3c577fd9030e3cf1886c97a1c95ac334f728d300ebef350da8767e23fa3363e1912efb1ad84dd4c27e22d9c9e7e927c3175506f1c3b119f6f6cd7687ad3856d3662b0c13f7dfa146480547bd5f7dc9ae89;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h66ccf5f031c07a8ae1f537b47b341a547402251b91df724923f46f46d5ff11a48c693930d0cde16b4e4756b5fc0abf1ab3efbd0d4da662d6c940e0459ef43399aaf2402affbc1ba4dae1db72dbb43dc3ec27f30556786692a6e1e09b01bb2b679460d0d7a2a0640c049dc1755cb5be7c55c77e0b32c88d51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b13210b6f23c892d45b46f0fd1db89749712e78422523f1c0b692511fddcdd1be0d288e18f94a5f4a2d3edf0d73a46e91f87f3b15931e180f6dc4a73b5f46f55073a1e9cb3b105cf3bffc17d8b6fa7891e229080a4417f8c386793fcb75b09144b9a772d49b5365a40ec7f21ebb4fa04263fcffa6eff277e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88eaa759285ac6b8215e88e5090140c6cf7fe2d84052ff0764e0274b0cc71a76348b703a0898e0d3d719bbdc633aeb83987c9986a89f3d1af192ba2bf29962f512273d35def5a54d7534fabf5ede6d321a09bdbb9d7378c879f0337671ad523d24609a57b4a4d6a499c4c7c8c23e5d6c4ff67635c6faf44f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fe3cda2deb3931d487591cc0bc55832fc9f4f954d37a98f4afe9b2b417d3648d4f419b4483a6b9b2e373e26f0766c10917c8fb36da89a76a807e055f59631b3e7e3ec98d62e75adae8e0e2807843abc880765eccdf8180dd932907a660242ed60e59e4c3051e75b99101e8a074d974a27e022ffec22abd40;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdbfb1fc8310872081aa42dc47238fcb0df3f9bfe37c95a21f658d852c7be81687488c50345d6d6da5016b7c267e2205b5c8f33c3a922dbbdcbf2397f23816f0c86552b4ed78871eef61588e42f6c06883866703cbbc2cf8b53a062f3291cd8bce1f865817406e2eeebc36da4a133c3e8ad78081f40ddbc27;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e33f5b7358d40dabe053802ce76dd8377c395fecd283d128e2089e931b6d29e0543e8635c9eabc9b4cdeb2e6c37f5976cdd4711a88167f270f26017a3ff8760a4ac3ff4f2adcb86cb829ecc85323db034c9e38eb7be2e0a09804109a53bd4a2e59beaf56b5b90e41fe6f5e64f6b3485403cfa0227bd4b995;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fe56daf157c9c6d4bf1ff2bdaf908681871c96398699915e1e256835e0fd5b5d0d0dbf7f0e0dc1e0b50beb656e3835611d378e2ca046f6ec53e3c3c5f0b37cc0e4823d3b58a733b1970520dd32fde92e289442804c2d7dce1d773c5d7ae378a2b85561f3eac49cc4ced8cff77947c51873e80b4e22c24e6c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e1607854da1196f067cd2f0bb5cfd41085be77e3200eb8083aa0db891a515830d454ec3c828b59536cfb344b1ed5614e9dd9013ad9589eb97705c5b46ce84b152b28278be70a001fc86bc69d9d7406fd3a7af6310a666d9660e83a6e1d1d2d7162004c33a82b787b0699bdbad4d8630bb649a910b554647;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h169bfff8c65c5124ae83a90195e20bfba5b0a19dc58b778eff578efe4a37322bb19810c05eeda7147d272d6a9fa0d8487d21ffa127b2bbe1de651eff9fe075d32b4f6e82c3843f59d9489ef024f296f11f47c7e6a143d90d7091d1e96e8aa526fa954d8c41e14445c143214aa837dfae7d164d7992a5bd4e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1999e9937448bc500d21adf72a38da8acc80445a941e6c949c5a321bf02d90965b742c5a980be34fc363856470d6e8d08d4c08bfbc8c1daf83752a3934d0a741549d3043bd2ba2e9e6d2a0d002a00bf5ee3276252f593919179e5338b993b3208f2a23d7e9a9eed29dd2b6d2a139b7b7595d99c4078088a5e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f55cf6274f4b483b94dfc8ad568f0d90d16e6b526e95023cb21b3dccb9bb394edd1e56dfff80ecc5fdc7899cfcf4daaf25666f449053301f9a7ad258951215a668892e2ab74b7255a5c8e269da920a0070a80465cb06422c39a95514420d6f7b4565bf6a398b3a2129d457ecf8b6c1c22624f5aff9a1813;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17501fe5069678d6ff6f7a7064b9ed69ae70ad2f8b57363fd0e0eb5618f7f288930bd679cc22bef2bf24be05c66c28ebe0ed444bfe7e34b734f0f8bf629043599295c62ab8c5e35ed1f9f1a80667f37202dc2a7824a82bc38a18c97b8cc968f557cc3d3252278e0953ad278bb656f87b085b2b5fd675975e5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1935cfc974831ffe7f72d76b78ae0a259223f90e00df1f9ef9c1ffbacb4ecd09174695ab02cf9939309c4e1e70ebb06d945097aa87b998598eed89a8a493f55ec50b80dcd3a35405d6e978403f787641d38ce9f864f3179b485f3ec4b8d6264e4823bf681d1130eabd33782b9d840938d9987970b6edd10c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h59864ba4bbb99870e66df4861bd04468e7dec4541974e49f311e71ed68973ece968377e69e22272def0114445116f4fa1d09fcebe93aeb8a31b3fa16393396ee2925c9778aac6d77696b0ea3728dd1e78f8572f2ae41301db7be2986f300627e164c0d499437c32e570cb679b3cf8f5e406966ff30b97f58;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bbbf576f7c2e8dba79fae2da092775f22f1bdda5c4c7d6cb0775fbba0536658f681b1042ef9093c5c63d2952172a22c2f26f46829322e93a7f2190e0a35aa8648513ec5195923cbf3554af1856157a30dc02dd159848fd6522b17655389e7d4930ec733e7059b5c8d60d90d3b8e630a7c11819edcc64bfb2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h54c4600f49c6e2a5ee351659c4be1b04eb5c36d17ff34b493b994ef1ae2c393fc9a0a75e750f30c765dd6491da339eac922cf1611204873412a204511cde1551cb3559b1511314de98d1837970c5e9583c1735a0073c9c564ca24328414d4c12f1ac4679cdf6bec2620bec78f97ef9afcdba949c8df7fc30;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h40b95427ebdf869e489916241c426e0c4492456a9ca7f269840df5502f506c327ac5a6c6abeff625703a4349a66eec626de8030bb491166e08bccf46d8b784362b9b3057d529c2497405ec56e8a8ca23861d88999cef4a22b6a3b6289538d02579b24f455d2afb88ed2107731da66a937c6ba5eaebc25a40;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h376c52fb1d421a16e99bd83597fbbc3f7dd9a7cf6bbe8930e46de813c067f7f7a1bd925decc79cc580e2a9acd0cc4dfd953754b97aa724dd39ecfd39a4c557de00295b738899f0a11bcb742b7e2b0c7b15e3d5c0e768e576889c85c53f51ad99116408dade167e8b920945b18846ebb2e349652f39440764;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17874235250403edb9bc569ceeb0ea1d33753a6781cb35e999d335574dc53826667875804275ced2e802cbf2fc0547f6440c9d3236932be19106cf040cf8b32b37a19d5a855b7d5af344b78985b1391daab3ef7bc698284bc31e0b618879b622993c63308116f3de3710b2daecaa2d765c5c4061ed164cbfd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdbfdb310663a5684b978d7a34e5fbbeebb30b1c08d4104be01698d43ab97b411008ba668bf9cd75456923978c27b500a68c8d0387c093720ebf628886152d1679536f08946e04f6c49f259b73fe4fe4a528d30afbd94ef17a183666598af0fde16b0f68a9699829548910b23e80736c3344309ba9a5ecf3e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e4763ed2a77ff0cfcad0ceee593cd94438ce619a31eb3cb408f9a395e5c0b4be67746f930e479cec5ceb47feea98c56b8457360493d08cca5ddb8cc6faf55edb6e427f2d6717ff774300a50aef5b6edbdc452057f254132376e50506ec12a79b9ca5c0651bd8071b170fc8233832664bf18378583812127;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f3e5ec0d2e8b4fcc3e67ce8bd26134041dd3f7b792ba48355b5da6ca5b23d236328c91fdf79606d2a927782ab677b4c393c89c7434ff91fa85b0c17f18afab5572e96935e93f8d0f0f62a791546010e2712cfd4b2eea0c9903a0a2f272f131ddd1db25abd88e09699540319b90c23264049d25e9afa269c6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d2c0cc57a6aed87388ce4aff15c68a53bbabca94cc0fd986e8935a7d80a59f426e3d9649b0c4c8624e1299025953850f98c38e9408ed7e16a79f1bf78f8aecd4636ed7abb779a63c308b9352bb8c14ae6dd754bfaaeb0ebbb97e74979ec255c5a6239f8641fe2083375630d1cf102f763d2317ce1fe76c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2fdc7b3eaef4bbd958c7dfb750cf4fc94f51861804b914eab0c4bff7f75578e5f5ac78045f351ae0d2eb52104762dc874545651eebaf861d6b7519ca39e8daf3ea8b2c66c041f940d10c919deb90f1fcb63a1e3342c17e7afe163321604dbfec5a68ef71bd141a5c70726f9c977710bf97429ab2fc195a86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e46120b02ca93cca7372267006fd590904610909277c358759f4c88185f8c67ce8eb5d570ae36057939b914ab5cc277ec34a37866ac4406ba9faee99dc51bb6579059475ed48c4c3e16b9707e8a968ee9d4068f053f85a2fbd5c8962699dcdc5c4491c4b8fdca6dec0e354f33c388d48199b6fa4eb14e05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118fd9942d7ee0b48b54f8ea166a6de828a38c492dbd4f0124f2ec3660f1b09318c7240313e412d1929bf38cee599aa5c61224e6966b5a5f18077f87135a17fb4cb638005f331b1eeb715b91585c6448cd349ffaf3601e6e686f76ba0b5dc923da92101abe8410a2259141f53fa240667389928e77f55d265;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14cb019ffbe256d057019c5eca1808703dc60aad1901d304a2cd67156fabc5ef7cbd18b1ec6f8cd98e98871bfb73c21ac937bb1d7b4008bf23cac4c59a6bacffda07c5124ff11cd29b44b0c5bf2e4215151bbe6f94935a9a814a318fb0758a5894844e812d60aab5190342e33d3d20e7b185d698707f14a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa61b7dee8d71ab12168e68000f68b251a920d807bed9a71fbf65a5e3441fc76e62d1a109635fc1ec56ed77058f148bb25e891b5aaffdec157aa0228521464e4af0ded0c52181909d4735d7a786e063254b477935e5816e4c29ca528079a22aa4fab7169966aec6a54390e7fb9249044b48d5decf7aeb71e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e60c357411db3216d7b5367d345b4c0e4403a674abe7502eaa3ca9db7290e4d5d16edfdc681f2e580678f6b3765bdcd6d1a8c2a4ee1cefeab61c04fb2c5478ac97b737b6adb8899c9276db6d499b5a47107150b69b2304083a40afdd837a9884a18ddddd1e64417047dd901ae907a22e0f6e0e6617a08bc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1346adf8cc0eba32950825c5488e58c5e63602910abc3aaf03d48c5ac13f93ae98859b5006b546708f8a653273fc7638626d3e5e338beb650be72eb7e141fe6965958cbcea9a58c29d041cd7581489c2381099a623349118541a17782d5cc80e4eabc995515e437fe84396a1b997a20130f3551ffaeefc4f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha37ba15153ccbef9b7b78bdbc88eb290ab25b99cd167e1ba884554394b4e73d1fd5d96c09b4537158581344c4fcf682aacf8a2a956b94f8f2ad66e9e134353dceafbbe045f2cb66316e90858f188bd37acac12c173762f9d1058fdb0d6109bc925714c91d1ac7023dd129638cde4fe99777e3622f375d3dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha49d28d4ddddf659f20b521608dbe917f901f8c196dd61b40f13800c7c3d54993d90005f0106c515c3ef54f036b8f390906d6bb0cae7bab2c5bbd16ebb69ed53da4f0c4d3a9b118e12209520becb72808288885be522aed220fcace0ca185e9808d50e7d609088961bd4e885d019536851afb5a29e422f7c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1533f942fffc084adb401d44065926eaa5d620722ec79070fd99c3c1cf51b9310660bbf397ad6a7e69cde602588bc90bd8ea532f133cf4090a04faccb2b85b87def470eb45cafb89fde50a8733f39ca2ec3d2cf0a7dcee4aa19cceba5621ae71bfacaaf0cf108aa14e17b2dee2196cf00b758ceb43fee7b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hff0335323e6f66d974623da88d671faf73201ae2e15ba20ad7051bd059b8932db6845ca68f48ce7ed0912e6c5705e58c1ad70b3d09053f8a8349183d48e5bfa46d358ab0ac8bcf44912f95d0fc49918c37edb3e672a9d380eb2fdce13c227a785609613cae1c197fffeb4a86f9ee3d76d6f537a1b8ba477;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf4cfcce2bf314d20395b3f4c8ec46d8e277a9a62ec2175bd5ac18de003b1a1d35a24355e25abab5b55409f8a900bcf5da73204d11f9a02c29042b9299a2a9651d01622a11c145721b9b5735153df945680b527dc35991a9c905760ed64fe368fbbfadcc70c1f49a499e83178cc1c585595f54d324a174abf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5f46217d960d855d5ba290215ba7fa330df54a9b3b2684c0ca62cb3388c427f60c612afd6780a43ea768a62e78aa392e806b972f403efa63486dbab8d1a544aaa00977547e17953286696c47a96db98745126a70ce834ccddc69334f9853ceeff38605c64898202697328dd03cac9deaaecbd5b9ae5435c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h718830dc0f8f5bfb231d91265d67e1e6019c5c8312dc128642e214ba9f24d40be5f6c24b4cbcbcd759dc846ae3160ed7f49a9e0722f0cc4d81221587b8d599d70f896dd099add4d97530f53d893bdc537a7198c72b98679928c0285b9d378bd76f7ab7c512710c8b55c52d4bd7f103f48e4dcc7038796e97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfcc039de97b1a221148c8398c745f4fdb1c06b7b99d76afcae93e3dd1c1ee4688f3b65c41b69b1706c2e21f04d0789f487d0b4bd0fc9cd737bcae74949858a668ec8b79fa52fad14a5756143b10e23f6ed2339ec7de7dca931133835600e2600bdbbc268faef314d4f774d3b0978109653077833417e6899;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10253cf95c1fa81a086ac772cf0d8a36d8550e43e5ff8c44b1038399cc918f126abc68aec3f232795599c446f7e577ab5e6d22df85c0f92d71b3534fe0c8895efd7c7cd3413c6f988d6997f6766d2ab704754c8aa32a825898dec77dd5fccbdf8283732080032abd14cf504baaef7b6830f49ee2688a5acb7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50e3d755fe9271036f97cba8729b9097b88523ca0744e019c69a971219d64f54d23090fd1e569542fd44c135152060f008ce39a92afa0c98de9fe31d90093d3ab95466ea5d80e1d41a6f6479a7a4f7a625a2c50e3ff4325d608c62761b2549a312f02f22aea83e4fc20b22a3a07cb3e894fb7d63504371ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149c317ba728ec682b3b1581e7f667937d7cead5657e44784ed077f8eac9e9a3af2648912cb398c7774465c62bac1824a30c1fc832cf6ed6aef68d10b225f8b0dbbc8b97ce9f9cf862b9652dc524b5a4f126b5dfe1f70d1d4a2dc41104fbcb7d523d4db024b6aacf55284a7f864a7519b7fb29f2cbeed53db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14a84c8251f86d2f3bcb40ecde67699c15b53e3504643cd2fb0b775b572927cd3488c5d84347f1c17f46f8accd3fda9807cfb4998cd78e2626e2aa54c14eef8b1ef76e1feba2485f437971802d2d5c6da964bf8f70b45634d85d289eec05db40d28cbe6cf109e72ff8633ffbc8f31734b7935c5d3af1af1cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1723add826283c2c48dea74829b90e36244df8e35ebab379d538258db457b69f119c7c5b6ea640c3bb9a9fa879c4c1c1fd94edf7090e06a9c4a1d5ca14e43a7e9632c4cb781df0752dece6ce7e5abe3013455921f52dcf78dd6f0e8880d1c24d706defb7b24f6f8ef07f6e1986ca609a3f20e137895f6a215;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aac2889c1e39cd78995c24fc90d318a01c5e0f365dfc9809e20d2ff1d5cf58ed292a43383f4740333501a0b0380274a006d2a1015b70038015f4c21e41fe2d630831d51d154ed164f9a70c6019b66543b39f79d33d2486084f4e69a92f02ba4ab4facebb96cc7fdfb28d65edc1f314874bcc4763b9d1233a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h197ab581368cfe7324a2d7e5bcbc3e01f02a3ed831256ae31e39baf16737a60e4d376f564b3c83d3eb12ef6152ac5e13fac3b97ec38e7d920658d7a7c568df68a1261293601f3ed0f50c0f47d4bef779b0e92f08b79fdeb95910a867debe4cd662e147912241584955880514d9ebefb9a15d536b98d36b6fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17bac39048c81d122c2c9924ddbd50b54959ab308e8bbc2663e18b7b771fd1670b69cbf13911b016daf3f6210b3af6ed1008c36bd1fdc8a7d3796ed5eb7a0cda6b541c9088a96f62b0432984235a2b774b3f6eacaaba0aca50f476ee60f881754d8811d0e4aca67900bdf3cda56f5d6bec0f1aa474a8ce1f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14dbb61088e2a7df48b62fd3ecb3ebe3b83ce8f865f816ed72acff5b38f27535a8545933764b809ce9cdb3990fd24419d519722b228274c982be9c86d479e7d5c60754c0a7c8de46012e3731ce956a967a582323c26639dc81ee9a506cbc1fb4073576d3371f9d3d223e9705910e3f691a57f1ed779bf3e7b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e353ae0114958a405d0a306b68616c575f20faf5d151c5440b3e396e0d83cee834fec34c138e48800fac79039d5dacb5210b8a2f203fd7b5775dedcd91931afa225fea81031da115e3c09dd026337af9939fd7346bb19044083f4217184f4f6c89db9e867b3fe4b23fc4d78f766aa60204fdd074f4a1f5a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6af4a3d0a877188db93b4df02f740298b8785c41bed2c8d6c17fb87bc141481dca4a5dd4dba2c328fc243d65197330f1f2e070b6078397dc56b234a54978b709040419f7e7e56ab9daa865f6191f72b2e5719ee9d5527d2e54daaccf45623bd58ebadba48a2ade72f47e16e93e47a1f7f6e5ae66333151e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b0bc84bd565a731c5c2922caf224172e5572d020a4276805504f92b51553560ffd56e3622ef8124b770fa8118c58e150dbdc3571e16bbf0b0714bb99a9f26ba3db0b9526a44578da708005f09ff482533a763e5705a268ff18ad8c23b4b915106107bb9e5999c1140650889c7da071feabb96a2a554331b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h832bc85c97e82fb5a296cf502fce6df9733e8fa1d6cbaed45aa0d09a7e98b6ba5311bdcd8cbb616c8ff1031c4b1138181d8bb568fcb5cce5da4017af0e9b313f7aa1fe2d2ba1fe6602cd444fca69b74316bc2f18201d4da26196c555430ef1869251205138f712aa2270287e13593ca7a5f763c672f39176;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d57e3dc4f01f4fb897177db5b9f10be7d4d7fcbba09d423cc7092f61740a123b390962aae1b46d4830e7ed6733f825ac212914febddf2fbd4b426c268867debdc1e4a9a1dce96cee04fa2cac5a2c36bd6c0e146f5a15ee9a9098db4e7631475b4033a3b1ac2c9cf10479ac3f977643cca708b5ec45622665;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a46e284c0a4805b753b72faea3119e6c883ff03d1532603b05fa84917d89a1485025611237258e8b9263908f7b985fa50117029996c88d0ffb66be362461d4c5a85ae7736a9aa34a97366195291b3392d5686c57c98c6e6c2306a501979d5d31f05a1c195fd9b07a363d0dc14690aa140f6c56d901914564;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4b873cd6f3bc80b4d12bb75e0f71cccf3d71bcc5b4f893a6577f3e0c43f6f7993667575bb1a234c7c96bf75c18f6eb7feeeb9050dadb8af5d13545a34237d92547a4deb3f03d02bd3574a8e5482b957da5d49d6c1700b1e9110821a5d48946070a82d64f79d67786ee9b88d2a703819dbf9364dedb04bd4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15958454a4000ac8de105c3fc5c019a50ce67762f4ae782c39122e202cca0e06223a7fba14c8d7fefff85f77a7c13437559fcf677e5f855b1c12de79c2e800c14ed4194a6c4ba52a716740d203bf4320536b4e76b1ca6d3a6582f56a132d8fa03d99017dec37f83e6e46f95c0863d679979a26059d0509b35;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6708bdb47f853c032e9fa467395a7e30b10a4d9d88f558956b673632163cc5e9ff0b88b4195845579e6388d83060f2efc37bcdab981d7dd39b0a3b31b1fc01c53423e832da7dcd1295fdc918c5c1b69f3df21c60e8b4ec5a714e88cb47d8acc30b818c7c59245feeeb814f01f5aafea0cbcfb69044561abb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ecbe5eb78b77ea07224e3830489dc8728a0816a98ef83e76e26c03c4d52a649d5f3a266ed926a02e8e16367fff19110816aa8cb8f4085b8897881baab3c81e8cabd3f81d11c9ef47ea2e178c345c291313af5009adea2abfc535e5aa37fc369037e3a9225046f92bf2ae7a9b6765c7322d051f8a820c5ac9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10396dbcf4840b377ee616c7df478395a5774ea4a1977633dc2898d6e0c02af71a9e25e49eda419b589f2fa357a461411c3b679672c3707f43e84b38e8245a8dc573966a9eaa985c8aaf3216eedd9b79077cf9e01682cda2fb82072b2d931b99ec86fa0eef630147a2468f9679a85f03e90ff271240a74a03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h819d5ba06104b8b205e8624e74904497356b10e5f724e773c0495be1122c202ebee77895eeed2ff35366daf717be42b10c021a62b322b9a8a49d5d1ae7bb9823949f4173fdd18d67a429fff7ab71750c51e7b484b868d4cac19bce970352465b15c9469127cf0523e67c6e37fec88d40e6a91f168cfb96c4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd161387f5467843c25806b33f767e0af023fc31dc9c52d675f6b443ca354dd0e306fec0e64b6d1351a1b311e357c2341b270887c66497462e1d6ff21817249a17b8fe97efdb2c248db8e3b244cdee664c9c35b647a0faaab91ab7dbab404ffc06388bef9306b6f8a011c664846d974d2bfe49046a05b07f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5cdefdd97ca7663a0d0c024f5e88ea18a971e21a85b2d46e04eead51dfbde9f3fa24f900dc6b9e2b2bc4da95aa90c1f75bf855c63aa67617c4f6f4f6699a32ef9b8990b14198b9eec2692c2683cf948ab866e5c8580804070c718948135a3424d295eacea16ef987b5c23d9be77553f2cfc4d35cd74f2ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb2644c45e9309e89aa1d3c6e0126613450d264e62142e53d25516b9eb55abcb40ec7b3ba38bfdb4eab208a47f6d38084814f7be216bc812f25b0974fdb5a1b87ec6c71db4170deee528a91bcb937ccd275059aa776364cdb387ca61bb5314b550a5e6ac31372a4374c54c041fb08aa223c513f76ca7a29af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd37eba19f55be1557e48eee0992db9c6fe8ca18020feeec5d8d018a4336ed1a07e8ad8100433718701a631cdd034fabc1fb23cd455aa2172d0858a04935cf22cbe75ca6ecf59982ef7a36fdece75eb36c75ec9813101145f8080afe28a0e4ca1437682bcbbbc50ed2f31e54b8c24ff3d9a7ad1ee164b43de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e6ddaf1f6892af2410a98ed3953c9ecb80e31e27b1d317e2fd3f93b39c8cc074c9b85f2eadac63c85f8316674b1304ee7b4c507f42196227a0550c1b2db876684276b3a9fd31ef992ccdbc0881265032c6e92c5a546e4af684c7cb650f97e6750c52fa2570d66a6aed8a56fcb73e7b4ff71bd79afb32ea6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h60940b16c6fb2710d0667ce5eb7c0d05b661563557fe62c3a28708e9ecf0955d285aa1c4eee3c1d9195a242dbb15029f187764564a551a46dacbc047c2157f0d0fcb4c56659c6dd0f84f44ef7ea5210c6fcbaf295d155828f177b0ef20922d4794a6d7ed256559f253af8b93fd299b81f9751a75ee1d98b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha81c3b82a09fe3a0b2b3127e77e2be76afefee73efbb59178d7545e1e87638f2e295b04aec7faf6bcca8032037ea352cbf84cd9ff71525bfa456aaf8a56c7ce72226876c72f9e1558e6993e201420952f2ab07925876e61bd4fc99f25d06900ad86fe0a3c1f89b2c03719a2210d773934317cff2253bd848;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16cee48acd78dea4320f041a2943c032856d5e8fcefa0e6ea6d23c28bf854416241663ff1fd35ff74ccb5d2c6ca74f5617e891577828409c9677cd4c75bf7d5ef4a720783a0b024f5d15012ef98d2554690aabbfa087c471f9249c8716881c42852e9048713389e8c4aaecca82d520f438cbea39f815aaa91;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18b0f4960a1aba109707cbc46afafb4038ed8cb7969b6529c8f80e9ecf7e688c969b05842446ce83f26f2811d281ec1248f241b94439e35df7a0315b35c64ddb46d4ac2be419f2afd047b085abac9bac244f30b0664bbf7b5a380df7d9f33733457dc6932d7d3e060139ecc32b4c463c2b6719a1d41fb95d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19499c248a4055b6a044f5b5607ddf6d23890a922b831aaf9cd09fee4477beaa8770d0aa521664f8b1582a52139fde10221961bf258590f3dc3bb293e5d6fbeaeac0f0f62e019e805b0d377d1dc1a71ab586360faaee66c038ac9c4ffd7211f7563ab0dbaadc004ac85d6ccbc2c89217167989cb2ba95df1d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16513fda609c14a3d0073bceb4678340168622debe9b31787aa8b21516148a6ffd9ababa2369f1c138e4f62a7efba7160215bc1e73714d98104e0862da307411e19e6c7de5e905b0b2ed10aa395804e66644f2f4304a96da2c52555102bb8192cf6af660a429374769bb17908c005944ad5cc36d3b5e1d26e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a733d3dd0fdec83189aeeb8db2a3995ddaabbd7469aff07a5436fd1366fcce3c55b8c975ae89c04764386b59ac44be1147414c9492742583c9f28d2b7aa93942ec1f6234c181d3133bb6ae2ec5de61f7935de4d0c6401a17b3540198afc98c4553bb24e374ec987f51dec322d4b344e0c829bfc43ab6a441;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h176e8b5a5c2226f93037156cb59e1f672c885170dc956af90782a72b84fd0a81e05541d7ad76034ff5cafb9f4a3286d384e75ba7827316ee4d25ea9bef87251ba707d75f2618cf80096945966256a2292db9c2f34716e0bf6d4855ccff036bcf039219b3c33c0cad231591ef9bfc1e82272fa9395d7373316;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b19b42aa304aee8cc90a839c059ec93b8d7768a3af8187ab1e75b8914c2b7c7e26aa0fc22a71342a45c86a3e8bef56f9c347ea5bd4e88ae6ef388c15b503c3359f472e96a047fef14eba5ec5c502ea5e2a2c99eeb7d27f3a0c24a6dddc162cc570aa5b6e816a50cb755e1e19fd104a0b2b0d9aff7b2546c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1786bf49e203ecc0cd64b88d5984921c9068fa3e60e2ff08772960e8d0f56a2fa2c2decee04bf7eb2bd3607c2693788c761b175cf9dbad93027be4a189fb19f08c64c3d3d57e822a65d6f12563de0c3795c874a63448e23e80ede12f7e971775de9dfabc78ba83c1964aa943c8a4106685f02e4ad5270d91d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h717cdd337208d98253e483b64728c0a7529b50956b33e86ef365d0af89a7eb9f7847ac5d9afe1c4f69c0c5c6a781e184c35a7425fc9b261f2e4ed945d957317b145ddc2b9fc5a7b73b86513bd9c544755e1d35cde7347faba958b7d3e02b43737f9a0482d8df13db62f30f6f85c6672b741d930a55f52770;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2356fcaed18a9cf39a8730f4e48f78df24355d443c46ffe6d41de916adf1ea8902781e1987989c82c3fbdfc4cb0cd9bd4fa7d34049303c80682fd6ca05123ad6453d39ee7a89545d6e6f47570aa85c4b584610180ae3dbd73d39ba9d23257d14f35b6a8f9b9bf13b337df675b4fa81de00c7beb561c5477c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hedac14f55e4a7b833cdfe7b9bdc31b6af697a4c2ac0de1ecb0b2e793dff287f0165caaeb670f53035d971841c71d98b803af6100938cb4abb3089691bdf9355fd1cf81f1848477bf427b516e0acd3486b10b4f551b157d20011c93d5d3fafccfb2cf97cb3bf14b18c4e1f5d93f3a809fcd31221167b29a02;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fbe8d10b06fe4b1ff33bd501a204afe6ae0b34aa4dc11ca04558ca19f0d9a4f55913b53c96723b27504e73ad610193d9cfcbe9a9712cacc934b4b07cf450098dd39067362e8a492dad48099538887b09a7626c3644d03cec35a4c8436733813d29c3dff855eb35646c43411fda89cad7a6df388808a1471a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ae7fec255b37b356d8864bb0550d872d49387a591a6641057a58121378167086c5f653413313a313cba648abb5f2db1eb9f223a23147d572547ecf98a4332d700b395e30ba712dffa39245e524c87eb0c7f02170d1d67750c614ef0a259f018c75cc77179cfe351205dae16fabde96c68809a54f044ff17;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d1820868d2e556c6f63c3cfa257ac6d9b00287dfabaf39f54840a359706b01db317aa1e9300c13d15741810b89ccdc31e547d0e073b5bf1b50232837b1e62a5340025bcd1a0dc7d2d2d1f58357d5b9e00e9d09cf5df6c1140bf538cf9580cde9b53f1f7794c6c46ed8bcf5e4cf0c5d2fc884d214565a1516;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he2d230e6d9fa4081ec0e6db15c60bd014809031d543bcb0b500f5073cdc07be3396c745edb8e4bf4660f687418329f47e8b097f8ae6423a8f0f6efd428f8aa5a595ba0da4a6b92b8b256f073f8ccd83cd994f96d53dd15b2787703e7ff938987bcf22dee081a943a4b71c1ea6b6c0099c2a6f340fe87ac62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h183d2eb6878a5db06e17d96eabf4951b07f047b13074c1190ff6c0c8462c9c443bfe095b7e6ba4ff0b0d8707938e1c3bdef588452a4590015ce45b1eefccb743aff138fdf8eb7879ef34dd2422b34bf4600ce4bc043edd09dd9e7c3079853c36cf282d732069d9c1b2c76ad341ce43420b2610c66985f35bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e6f11ca51317c48b25933e42f8c3e9c18397eff29cb006fda927cc819e113865d93acf1088ef9b036e6f4ec3c0eb79ad2732adf62be2296dc0cdab4f3cde2ac2e8cd256d0eed2d428b1be90c07292e783ac74f150eefa04547144bc456218e145a0f5bb996b7be7644b089c0cc82bba2d79cf09d2a76c2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h20d2f3a7b8fa58355cfb479148f6c656a2a06a50f0a618854f507f51a3c5a02a64dda22bc2121083a8bfac807d1e1552a9687bd2d9c146f42ca2fdd43f00699bed63e5683972d97230b127b0a224df0dacd0638d86696beda12a255d95aafdb9ab0d6db9512b7ee5fb3184289a52fdc0f42137495a22c65a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a47a1ca778328c66f248e264baeecff8370cf66d77f1beb7ba5d6cba55dd53db3bd10b73a35cc473dbb694e92154c702aa7f84c090243a9a1170d13421d2ea5d1aba47da38a07b29a15bf6a5df47ad634cdc1686bc4d4ce12bc79e47fa4d4c70036f337397fdb0827df04368de77df6de09cb643626e70e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1096215d3ef594320ca9aa4dc6640cdc584822f1040ca5184c23e15f4bc6090f0f3b47b034a134f3ac520229fdd1f9ec86e9e9ec09d6478600a3a329a1d0c4607f0052c72823b129525471854111aefec22b7a2a00ab7f8c825818d4f72fde015eec96c54d302b1aa2dafb5cc09ca384e4be47ac66d77bdc2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196847f49ce67d32e1ead5bc3484af6e933f5b113a363c7b3ddae316c51d14cae8c757b7dd080dc99ce8bbd3c47a48403568190e2ee74b10bba5c10cadc5f6dee0c399a81c4e588c2ba348e84b9271289e74b172725736389ab77d2858d851f07db44289fc9016fb12b2ac8424e5a63fa2968a4e4a7dc54b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104fcf0a7228307bc79370b15f1f5c58e243b759553df3e710388d1f3ba41e4b7de8d6aff8b1102c84620af3f03d2b21a0b2c098d75a4fa539c5e646848201ab4846c5b7fedcc0b8c7e437ca97d1f9b2ffabe15aa3269ac3f54b48228f446d2c21843e92534fc7e821e6c8490b1a2349bd90d5d3b349016f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d53339d3636a4f7df076334cadcd42a21f4cdfaa06af0b6ee998fb0fbab075cd270fd93d3352e0017dc0aefd0b6e6d8914de456eec96061da1302b4363922d7c3af36c069a3c15fb14fd8c136c64d7d0cfab405b940bc814ef602325f41de348c8e9990628051a1d9e29a87e02a784d05f9ed938dcda1d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c4993900f6b6d37adc4ed34659ab5def7658baba7e3a7e7477147b91df4143c0e378096d67470cd9b402e280ee3308eb83926ff50e8c7cce97e4b21c51913e090a6622bc984728d3629fa2d1209b3c514583a2e896b01133ae0f98e110fcf079458379ee4ab321aad65a72e31f2aadd9b81aff038ca1e06;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84c896cb6417cd57f8048ece3778645ac09205ef052c361b69d49caa28ceae51db5890d9a179e2c3dc2c1d6139c6b0bc98184b39a25c12023f6d14d1dee9d9a9d09674f17ab68992bbf8b08165cb0dc1d372a03eca84e979423b7f782b6b9ee5bc26de7df20f0869c7b8733172a354e713a62530e75b5736;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h31a24d62842a3f7d51a4c197d4a173c7103a7adcf0e22ada17c6c5259b80e9959ba2c26ee1c8e332e6842546777a69b6e25c8c2e9d189bfc18a5edf400f41f29efc08d33bae472046508a62f6fcab15d2d39bc5f42097f834bc7b458a3f705c7a1b6d137383e8a55a3e85eb094d08eb8e150f1e6f91a3e44;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19282035e7000b50a997809acc1037237e1a45e5379b6f5fa165317a760e573a146fb8b4e8b08076ccf176f56cc851965af0e67245294fd76da0672e56ed14d351b6579468205d62f7e4bfdd622e562fcac4bc217776c30bc88f02e5852941d87ac02df778c4e7789a78050f96101f78207532544066133ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d1b5f3f7e427f91858047aa2617526ec3f1d4623217351f8800bc44288d17d31c2750bb722083e07d439b74948f1d88783aa651acfc2ccc69f7503a0980aacc1cd16a81ccfee77d551d3df6c332d3a9ef77b33d68783d62a4aa94b01dee3344498c7a49fe784c7cbe29cc0cb50ebb929d0d64ed892aa1bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h86f7b6557a034428ac2e242459827c5e15ac342cdbfe96ba67dc07ce92ba91ac77e785f2caed95daadcf3da55983ee576c40b7109ffd22a989f52af37f0d806a28ebaccd356960969ed7d129798b84beea87af6622e28654b2fc679361085086721c31aafb6d3bc3c2ac5a2bcc7f96f9eec244d04123f318;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hca177c975191a839be29752c6783925882011bf089b5a5f7f8876c687e7289b65b1089e34a5ef0fc9ff809ad294af664fd944b68d6f8fb9ca261269c9a595202a76490189286a73153b490ed0c50605d5e7d7569ab126200beee9237948f719ed7ee64d5f390bc4f9e6e996b842f1c77b021fa6c581dffc6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47c9002c972aa9d85251cde01b977541c76d80d0e11ef73d79627f67414ae58c21cb83007ab5d7b63949fc7122f3c03a2c4d71cf8b1b6dad699f79d6bcb14eea53593c7ed1fb91ce90342a11203fcbabe856cfe930029f112bdf38ce8228188b436ece6dd026ae1cd64308bf6984dd76a1e3c035b30ae787;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5825da6f0670937fa48a7308fee915f30a92ddbacd6886c6b9f8e1dea46b1cc23ed2160ab3362558bdfae046e28c0f3f7f0c48500cd367c5297967b1b6a2f340aeb504abd41b17feea1ffeea1304cf914a37908b98399df093ca88e693ae81c2fb407f66116ac0f0f8e16cd318f576cc51d5be815a560578;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173e54ee3c08f976171ce0725c264a6738943587b927f6bbe1fd8be58933306ae500c7ae8f5757f936ef8d15f54e0da56dbf82d9946050db24f721d9cc28b776ba064cf02fe408c450a49e68400fe34f1d901b775aa9939c7a494b6e19cc0ebf77613b9f145cee3b47037d1257dc69798419c3dd6fec910d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f18156be0fa2ecc3dedcdd5153c4893f422f85d0823c682da7f65c9a1c42c4b54c1f75ac15115159315e06953aeb34c6f84129beee807d312a098d48e49ea33c63145db33eb72e4d2bb0526cd99078d90e5402ef6d1bb96a80e6b4f4822f1ebd3453cc6a870823f830478cc4331ed5acd6a0e885246503a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he177abcfc48dafcbb1076328f2ca2913d68d06d341106767c3fbb30beb0805ecdb76f3ca3a2b4a6eac6c0498a3c03d9ba6358217b02ae95f621c1f61d04032605e73f32a065849c114a95bd11cb25b41589b72a9ba4566652560e0d091017800dfb40e5fe7090400a114b5d319411d8d0815ba1348640d0a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9819c979f85a98847acf106992ace667e86290650855ed7afbcaf76952a24db290497a8a21a4e72a6c53fec4e0b370a3d652dc0a7d041a80e9759c8e93eb8bb5d9f355a1aa9720bc6c427a9de2aaae99943e5e2335227931ed561f9dc7cabfb027c0206ae0ea319259cc7fc7f55f46a648f52e49cf7cc22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfad46c17e208d7462e754e7bdd9e1159d33935f7999f762b2a8e88f4d4b5951083127cefa1315ebe9dabef7962e378aebeca9a2428b82a519edd84cfba1bb5704f0f78020fc3d73cde0eeff07bba31f3d1f8c086cd425bdc6b9e595e9c83d81616724b9db6f293dbffd1cae58db628580138b25027a57742;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe3d6d00cd26ea7515bd897a3329dab32b0ea7a706eb1e50d575c71c9d674dc20708db0f00fac3820f53d8b5f34415c6cb928e332ac8be05174489b96b29ef7adba3e74fa5dada3995488c066d5c0d944320c29a12bf354c00f2c1939413f9ae5a917c5d4dec1a47a9df315dadffca00607dc3a9cbac3a17;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1af33ad93bf512e4eae2cf215a87ea367725a8dac5cb3370f3bbca3aca66d976ccdf31e1cc2eea2d9769516bb3e7ec169f6694b5864b149cc5bf4dfce8ff35c3ec634edff651a8e60d03799798417d4990143ac2cab54bcd9f050b3e3e9093803192476a48610cbe316c6b1fedb4620d4d7f01e5b1597820c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a29dedb1a46559a685ad1f7307a62ff478304cb1326309acae09262d91b6fcef45c9f55482346c0ddd0b66c0d58da3abe40d21e707b73cd0d0a66572581a0cd9408f9ef7679c24318d1cbe19a3527704aadff5ae7c5d393005fedda51c3ad2626d05ce67132cf23acca932af024c16e695de13d28483faa3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102433029899c4377de02200437718b785d77f3cfb321161bee97c750a7d2d5f9a2255ad7a52eb0e65666def68bfab0ef71d8bf5565e92c8f12fa2cbeb754fc0efe134a6a9aa7ae8036462f439eb43c556d5f79bdcb9720c21e368b28f2fdd7bb41ee231d91f4883e35b682caab9d6e400ae1e7cb4c9a22ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf24773e78b3c4f31cdd2f1a184eb69afea4b9b4befb787490f783712de3bd4a45614defb348c920c58339ee91d22bc3d761d2a911da61d4121939e43cf9fed5f84233db55c10436479e2ca0091ea16d4adc38a4f8c04c082c6650f1290bb6920e292fbc1545486867dd724685ef0825f5914a6944848abc6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfdfbcd8cf2dd0b3306b5a357e61c580c0958bb2bb50341cedd2388e0831ab6ac3f4409ba383456b8463378c082cc94b7ef5477afde85226dabfa17a916ed23ac0f46c14330c9710e849b9f22c0f6a5b4baadd9536d29f7b9e0ac50d4a3b285e070e76eab2da30e51394fe1e8f1f0b5f4a208fcd1d4765902;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e8867f5cf195f845c08b6bf36ff7f28240d4a32f9c6bfb602fab7f5e0a07f34e2c86b3e8368c428aba30e72885500507dd40af2549fc099c5a8d3a7a3852cab762d687893d659b8454726807cb852a5e9283d5c8882ffcc36b47f56fedb031eb91381ee174a2a383d5989a4b58206f1272e1d32e94bbc36;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a402bd1fa86c794f0ac93d917d3737294ddf0ec9da34d261b09292bf2655418ffbc9d03c7e5c856582b53e81f5c73dcab87cf897e228bb793922a3b0306a0c2e3de4807aa6ce74831c5311478ffa1ddb7589e676bd6b79560a5650b2c94355e21cb321ae7436cbb207f843367671e57aaf7ab0ee3d8e515;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h41fa2f1615290755967299d9abb307c1d66c5b55c70b166d86aa37a6bcaa97996dbb12538a4d5c662826189a7231f225fc483bc45905db0665854f2e86bf80294897cedde76048e964011229b28726544b08f7a711a7df494ff1f8bce4808dea7fe1ea7c67680ecb63e00cdcf2a933931d7d7bbd5b1e7bcc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16369e64f488e639f8d03e922ef6a67e5cea28da15cbb3672a46da5b28c950918ec23f77968b23ee8e0820d7b1fc14439ee17990b904656c68013963415166688ef9dc32a56442f9e5d9a8f06405bbd84116c019127eb36d589c2a1efe907d3df606c88209cb18a37814c22f77d7d23eb1f92b42ecb9b17e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had6ea20bcd0092fa9dd1a91f6b1c873c8fe8096aa47cb1c6765d4f43bc9a9dd20b07b42f8cf522b5d9cbced9f1d10ebf181fb80ec7b9648877519f3fb35c68441ad8cd41d1a95a9c3d8567728303ad3a8d24a153297aad216e6239ad937d5435d8a4aed8299986074c2f082672b413c7cb0eb8f5c7441362;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd579463755a6d4fb20212e2930a1a0f8283a063d6e893951b2935e9928f2d0c9fa0299c3e5b97d440e92c8bd13ffc64648404d8a27318bd203b834ccdb6562442adf50a985fe97d28d6b5d8b5027324ff48f365dd49d8711cbb7250449afbaeb453e781e2704f663ab50e38463dc8548713dc48ef075560;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe25fab1064ae0f347d99be8b04d496a1d4eef3dde73d44bc3fa02f426cce7de09740a749956473d336d2654f5fa61c494806abe46050cbacae3a340a1452a98cf01e6691afe350f9bae58b4090eb740493e64d55aa4a8f77b04c1394bcc2d8654b30f61effc24415df1f467c6a80119a2e7cae231c0dbec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e516ce1bac06073529d57eae091899b264658084717be7bbeca3faf17a689bb52e168e7daf03346f225e6e33a2e3ea5899c3dd069d4684651ceb7864a2d9b0f0beb7eab3e802164a9bf1c09c49a9bda77070b859df810217c2f52c2be4de32dc1d5ae97ddc9ff6cb99e3b443d3e3d38af0ae3c45407433a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f132e23e997a8f8b409e214abea7e4c576a6151006dad666f9d67d2b0de037ee2f52f6f6b073cb2d183749310e0e607c346a9662ef445d3f400af28ae92d84c955d6d74a973ddd622862424dafc0982bd3c12718d593d0805424fbccbe0e55a9189230dd2ff066219ef4f69a511e25bda1be18d279b5e42;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h184ca80bee98a5a58971fce54820339cd014a11ba75c1ccf56caaf9a5ad35f7a3bc9b3193b3a660c8a3d0b6a314493264a232dbe446cb4ec7224c8474a4025f7c66ab5063ac3fd784e7a4d02d38232223910d5b0eb173529bea164986d127faa5ca5c1536b0a297d82bc371169dda3a97d6ba2734164429ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h48a51cd62e1ae7b3b7a72ac3ff83159fea22fd0b1dbc4cfc479df206a8adf849609f89e75d3ffc59930c1baaf7415bd7d0ce8cabbc4a37f071eabd843506b4dd6c2d953f0a6b85c4e06c7f4408a9e32fe39b669bea9510e68582e7e24dac5c82b3278748f031d1c7bb78ce4f1c9a7a9117a132dc59ce47c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aaccea6e8485ab52a2e93bc4c94619192d3610bae00a9664508a115464b1e3a28ce7302e49929e36a1704c354c5bb948266d3f07abb303a71a5af08ff723079fed9da98024efb07dbc6ab8dbd6cf787411d7ed1054fe3b73134dc762e08ddd1b07bd94b1e797375fc90ccdead655110e32b4a209a97044fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h872cb1a2916086e9eceaf2db2311bcca002a8b10b02a95bd181b6295578667bdb9664f21feacc01dcab50984885aa1c281fc5623a32cd4d59292d9bc6683da6002a328d538ddd6cc3d5c978bea03477411e35b328b523a57b3b315cdfa32991509eaa07b60c8bc74e7df26833e5b999c96d68a8d34a67188;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h162f5a247bebdc36e5de59fbb1da7c9f64ae8eea97fc293e4b664869cd39f5bad106e702a5df7c591b33efaabbc75c0d2c545ea32e9021a12b150c5a3a77e7a296fd586e51586bb469da20a715ca26b73bd4351a3d462c4bb37bde9360bd43f4407866db95d6d8748fada1991340092b940e19a5115624962;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9dc5d0e48fdc0c1049872563b24658816109f22ba04f16a971531b649c85b82e329745039f3795aca518041d54b60bccf394dd438b450a041eabbaa40d3aa25f497adaf4cd0368aa3e780af2cb623b5ae2da5815c16fd0fa073493db49d1e8b31d97e61c39c5089f0fb586d8e57e95c5c04fed50bcb20f20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb99ad0ad4073a5080ed0dec6f3e5dc10995007e51cef1d67ce1b8e003d3cf14b7bd65d990bee36620964ffc0ec71986ada62c21b4d9315199df0e7e647e45087355a3f5f524bac79fef86e24d074431573aee9cb4964331a33c449d3c8cf73d34fba940c33ee037209ac3a618f8aecc06b3ec5ca76da70eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1f7f882ca9862dcdf909bafa1f8de66ef9e432f36c927acd3babea9bd2afa38b4c99fb3985a6c09410ad86b1d46507cb5a2704391ff519a9456d3cc70d255a6d8a4642e51615ce9d028ebebb264f59865fe78306b3d41d08525c4f2bd87ea44920ce4170b754a923247f4b21b0af3368581bb0e0b03000d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h163d3d2854bfe5bac8258d2c40d95559ea5d1e8ac76f0a8ee8c752e242db0cc2df1816999032bef37ac3ca0db4e50e4a0ad846c892576ed689d0ef1596fcf0f363ba8e32300f8b8b78bdaa28fba2f26bbc7710b0d30bffac32ef3f3a7b4c8d18639cbbfe1d454e54d8d2d593c9360ca73fd36db6c7d1227fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h56110488c2828c49c7da4508d019f78011f58830cbb6766099f7fb3e7b9735c5cbd66da1d1f845824c684f1da15cbdac1f027657de71af36c35fdae19e106a243858dbb34fed70ba7a98dfcfece4fd32f1364535343c3b384b23fb9521529f34188ea48f983939ca9d5fb272c6dba23fa5c28f201372141;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b3461fb4a72de70afd19baa78b31e87db12277edeadb82d565f69689449e3d4b6e749d93b8531b5377fa0a830789945dd1d935398e57c0e12b71f8e629fe0f199e4cf0915b66137f39944e86205676b44dc1f57cfd0f74b0a7cab1034c13b14b097662d4769e32238da2131c837e8595fcc13024c7be6405;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ce0f6eb58046cef9abf6cd8919075eeaebf44bc423721fe898a80a504f9e7baa43f6de8b7c5a51455e5863009ac0a45c962865f38163ba5c1c77e1ebd863fce4429d80fa6f007416b820da09e439182eb16c95e6e657e587e86d1aae0378f0b4cd57f151c5bbc3bda42bfcf6b10ecac862fed8ea49f6a148;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173a749e15cdfdcea7667db9f45a73f9cc311cb0faf2b9c6457553b0f6e7c1cbcb0d535c3e7b719ed3f69988d21f3d5625a4dd41674c213625db2596af82f1f94718d689b56ac2302725692753f3c56f80bee39e32b6613caf9867e83d642c62c09fd7925282e9f24d0f3b40f1d16ed859b0ce75f8c5e3c02;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h506d6c1715ce86bb3bc7bf0a8741c837776cb226bb654328dec734bd2719a9334eff16271e546da3b25da7c8706b6b95dbf5a48fdd3c25d4ad37cbd07f912a5e7c8ebde5cd5c3940889ef82409b309c10689530f9ee77660aafd521de74a1bdcd0242e63e4c2b76e94b8053be7576aac8e4558e5b7a46081;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he2d36a6dd16224959aa0bc1d4cdfaf7893620a255a50ffb94ff4431fccd63ce70b5e829bfd55ffba38c20c597b8e0a5c198c3679e59c4b9b2beae750bab4cfc0dc36f05a57a1e8190535087fc3931ddf3719d3c3ab1a43ddeb0a5f5f749a648a0dc74c78dfd1ecf6443fb5f5e2c1b331a7fbaffa8fafb108;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h796ed656518fe0e23f11d87f56786c7a11d58823cfa6859e35e5ff94ebe26f9b2759c26fcef419a336d1b886892f1f7762b84643e3bdf576510d2c296617ce94dcc07ad4d5e26761251508d6818a54abef0cc266d0b59677fbf47c4f6796ac5fb6beaa747e751c006ad5a91059c7922f372b0d7244876e5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c0f52ad1e7a95326c67f949e03a15e6d10eb4519d8f4dcde461af9bbc197db06bf2ab77cd3defd9f0f828326d18456849e8fc6b5a5d950a2c0c272d526557d3dc263f40b120c069d0d57fec694cef0bdc4a8bbde461826baffb1aedfdad5924f2ee1f17091de0794d25905a17cbf3acf11f825786b5bcb70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8f2a2adb5767fc3360b8c0de95cd58e39307226bd9418a243f7b473548a51b91d372f8acb632bd7fda300d9c691018c53d4006c918e5d57cbcd3f7a4c61f4fbae6ca14550415d69f37218189394dddcb2dc862ec672e0ea7c2e1108bb25dfeeaafc2b162a94d569fab95ed1aed156dfca07126b7c80abcb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a7289fe8ae78d5c08e0529ddc7e29c20510d5f95127c9cda494a7bd174f82da5b45cae6604c5a554174a3c48835b35c21fc5d72560770357fbc3e02f6cd2d927e80db4db253068a5dbaf2dfe3781ffd01d1638eaeacea4adcb5df8f84095b23b08c38d6576d82220cde1f2567d7a694b8b9e3cb2c4d2c863;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e8e1994301ab119949826c8733a5c4a486cd0aa6ffca0c54c91f2f20089e5ba618cf461df2dc5b992c5920fa6d01dc20d67b3b0ae81c946a7915e6a0c295ebe42cb1a0e2f71e65728e54b0b482143d4630b77518223b989ec29e3d8f9facc041c32be131728b73c04a1ca1556cb57f5081913a7d6cf45466;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f656336bb2963918389b0ae6a2ab0b15cbea312599a68ac584f407868f7f946c359862bf68996589782bbf6d6614d917dc06697e438f58ec397f0db36b5277990f79338fc6c1008f59ca602e5b45f209a5d1f7be5a2fe30c9913b71796c52890734bd0e964d98b077b049910ea3fba2f14071aa10e65879f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef42d402198bc2ae7c57bfd57727e6daa163426ce129d24c8e6ba13866b16c49dbdd9ce999afe65d704f07481a31dfd65a403be8f07f6f1ae1ce36259607119891a22803d5c95f07321e4a4bfd7b9aa0d0f3a444884b71be7b20dd6154a630d3544b3402cb47fceb3c8bd51c6ac277d83cbbae336f4e0170;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf920b008ebd8ee50611b73977eeaf253f778b8dc30a329b7e81e478d4279fd96f17b46e4278866be8d772e93f30252b3baab404491eac04b03c4dbcf12d340c78d98b30283850270f46b04a11e96fd28d95b382169f274b00fcdabf72a1ddc8299fa483afbcd1dcf1e7f698cdcddcb6f598d692cd7bf3c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4799b61ca60321cecde895e109340735374095de014eca25d1fd244855266d4e213a7088ad49b5e13ad48256e1e50ae22452ec12e456a727ef2ce433b9a774aed11548fd76341dbcd05f43b11ffa40f6a8f35d70649561c0caa9d1d70810c1ed10e99f972511325fe335a8d859b0daca9ca17a72a55875f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17cac5b032774a8eb88936842263c2c2ea3a04def9a85368aebf1a6973008d81c8618cc4579d38ec1f154bf84c9d692133fda195012d3727b653d2b4b82694499535a8fb350b320c8a34134cd26f2dea7a43017a595fec2acbaefcd188416c91c6caa7df51cf6d465d38927cd91565eaeede86e49272627f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h25679a438d509150a9dcfb1da3874aeecca60dd14db04cd0ae4f637f8914457e32c7cf42340ba77616451ffb78332d93ed3ab041fb465cfb8d9312a6c7eca62b34f1505fd10d2419cc95d2852b86a3a2a7c1b8ac46f7ce8abffb229cbaf9d29c453f998b082bee231377c6247fecb5a8a9fab51f8c2539b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2723593d5c37720dde0cc98523aab5aea5396b7e6ca390d26070bbe8fa5f29ef04632957fb5206d4094fc33c9b82cd3082cc49df1141871c8f690cf1bc4ab52fd8823c5dc57bc111f970c1d4d3280c29d766d31455fd0d263bf66b3ecf590d2ec96c905e4a7378195daff35b8c6b5440435e1a394e7aa4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8147ef7c3838414256885902ec64716f08b7e0404fb8276df1ced076fc573df8c5a16acdc3b82ec407f7e53807a8d2a7a90f17d8d5dbb70f84698c618c7a64aeb4d22fffc9bcb9f1114bfa121fe2727226b8daade6f82ec6a99bfe903b49dc2dd5eb7afcc83bc655d510c93edec517df003f901c14d7971;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h27507eac46539e130e52da4f83e3aff6d702ebd149308a924ede715f6ac2cd67773e2174b2709c9a474a40e24ea5d095931ca54a7701dfa8ab5c11dd918ee9b558d5401866a64fa500590d647f5a3a1bd239d5365d4bc5e7639130778f5af6eed641cc0bf1448b7d564d22754893c1c7f11a4334b0a97c4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h566ec8782304ccb1d70d05265db8fd3add86968751bbd5bfdc39aa218f642813ce197c734778959e2bedc93bb12b5701eaa054a641ff1fef6cb1a46b0062c46e1e2a0bb1d95cfaaf4aa26db01cfcd2c9ccfefc0f7d981da1389ad91f82c0434641f444cc33239ebab23a07a7396fc284ed31cffab4c4107b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175f141fa4178d4516246d0781c7c256af3779a4f652bbe05ac0056256e677c499dccad690cb8f3318ef4329bc0de481f378e46d945867c6cbc28d6f5a4ad21f333a0406be0f39146d7f22183bfc0901cecedc2849b2d0f520382b42ebd7e9e6d31e345fc85bd4d2ab276f970fd921e92006a5545cc46d21d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd7d5c360e9b2185a069e7c59fbaefab82a9e80a51320beae36c38d30906d4bcb68d7768ed4e55833787407baea1819d2b33b35a8c60ca1b831a37aeb25fe411a47f116d1db05a14bf8c16c25c11e89fd2f7b51d6c7df6e42a55129c6d814dca2f883fd6f3a53c9f951d0aab67c39c10fe3dfe9e68f8cea95;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h22624702c91d07e839de3df6fc25f7dfcc70d720b1d3294fe042b70af3dbcb3d51fb48c5bf8f76458820982e85b51b08ef3de6eb5ed234da3572bdc9127bba88a08c4b03f0ed2222088c270724a0b193ba0f06859a93024fc5559b829c4143961462cfc342152b685997f1955a886c345921010fd7a2ea8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12674de22c88ccf8d2684cc23504a9a94989447f878ec09d7dd71cac2ac6563de70d7f755e26f4298f10304f8dd1f307d67b06eb903900e0679fd1e176b532e14bf8e010a0e05b83ad2ec852fa151e04618fa371ee70fc456ea4cc8c933cf89620e9bf52752c20fb699b04d8142986939c0682dfefc91f5d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hea99712da0ed2a2b3cb07e3e2a32e120ef9c23b7d6c5789aefa95aeabc3dd125bdfae92c21fcfb544379152dc8caa3c209568c0d0305b4eac188d877762103e271138ddac45f3e34315824af78bce37619e4eeac14b18d6cc9d4fff110ef0f51831ca62c36e5ba267f36152ade84df3361d3deaca06fd089;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe15ed19bf526d5b7cc764bb617f58137f2f16bbbd60ee0e4cc236d0d650166f93db055d178a9a3e2978e71897140c1edb3041691b9cdf19e4978708d86a99564e98399e86bacfc58d490366db30c2ba5e90f9376a99ca7e3643e64637fa3218998221e5247a7f1651511ab958de36246561f6536f47c4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h326b8f6e72edc603b599dad174caa06d36a30edf2ec7d20f8cd53e6179f1a08e223f8ce80333fc13bd543eb4bc5dfa522ddcd5983884871de2de945a898f4fc599adba63a20b8985e17ccfd4f056814703fa4f86f50a52f0769827d7aadb0d479cdb18812f58dc7b442642de32bd6e7a6a0950bcb91cf714;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdbec892092e1b761823a190a20f4b564da7c7e404d399e5f9702a94ea5ad648f19fa600bf4f927a6793361c1f55ea317b0bbe783e0ce46adf7af837bed26b2c83eb00d7cb763ad84469ac0364d19e157a3bc8b8a7c89128b390fb4d0d3f0f89ef5223d72dd611b77be51df7c14a33ca761e5158bb186e97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3820bc4e51dba57fe366f0f2151ac8f9e1abe53346b762a8bf167e0066c431bc98f690a407d02c358e1fd971402effc480cb93a834c79b0a5d2f927ea336530164651f79050d6a44d0227580c9689ca9202e9be736bddee41ff6211ca25a0228b3001c6ee1da6e0ce2c53b59034009b69e617f2d9ee8ea67;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17cb029758ab0d39d51336df93ae75c4e6c2b69dd2d8c21bdb06949ff94c2235d1f28eb9a20a02165d2f478dcabc67ecb7a379a83c28b9e97770fc9780d01d431467d0c0a646aa147eeca3b2752669c5787d38c42fb985152f27d035cda4d21a575b0268cd62f3ddf022d020a1997eb7f8b93db260190f5b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h618783e2704392c9cb09f47810a5f225b93f4738912bf7219d59dfdbcbd12fbb7deedc7ee8a02a0a66ee479a879ae2f57e5f2661c3a60bbcd29ee18bc7eb36d8e4c6a00121d49dad7a8e543fcd1f5c6af9b8c1eb64ae97c8746477dd8743cbc3a43e3e6a5e443c0738f429e8ae8f557ef897e3e421683e86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he06ca92f18b9f84b4f8300d62da9dad0da2f1295af6542098c0d0902bf83a40bc0cc3429230b1af7d5f1e670c7112b1146e56315bde1dd3401357fecf9ac3beb62a1c31e7f08170667b5837517d21e80c94469342636fa72f05c890934c916e762cfaf8e6c82606d9fc1c757c708cfac4ff541257568163;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a145d1f3a839f640b0820247556d123464b7eb890025a7ac2faa2c1b322b57ae7c15636067e8cc7bc75585bec080eea6877ae8074739e46937ab9646647d6b9e685eaffd337c468002bdd0fc5b7fd689f378660eb5c83e00c4fd23c063a0c1beb0f3bc953ffb2b6c0927e321718bbe21d7010a45c335d07;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16d6e4bece899a37d8c88bc304f474d644cf4e55ae59f4cf678eb12fad525866422333ce14963c9ba70b69607467b2f607bb863d16d86745199d2278ccca533418d5d2b3ac372bcec767ee534abee0da1ae2e32d065eef088587bec51f8813ff1b41eb071cece398676d163311da301bb3d3cd41493fb8530;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h171b0157927b1a1694127a734ffc403f399696ba34a9f8622115c8d7867c543afafad277dcb39cd32bcc8927648fd7b850c202f946069a6d041a8a1596a6b8f447dcd7b1c61ac430396c64d3a5bca350a26c560d06fb7b8dad4de8468a389ca35839da69e4f848e228b651a9478490791fd6b097ba4c59520;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf527cd9ea2674eaaa09ab55d95aada3419d21022120d1a4a23ee86f0d76c8db6139a40c6f3fc1bec52bf4a1258db26c1213add13704c5c551ebe783aee5ee31e60558bd3e53efcdbb824d97533b859298b9533e455d1d29be6142e70f6ab14f2f2c00a708bd35c1c4da0e1e6866d05c26b8fdd99419f4eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h41ab6fa61384b7c3beedb2569feefc8dc6692a70a10f39ac0887744dbd44e3b64db412ca0b83c54c811f85c013c23b79fa5ca11151306f1a75300435e322d6064f13afdbe2e6e3fdc4dcc166c2010e84ec66758adecfa820d5de73b017ca731742a3ca7981bf64c6216efad950e3dffc484fd8bc82ac1230;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd36d04ce8f3dbec6af1f8348e474b1762dbf6152aaed158c38af3ab85f99224dd485dce58bafd14109f264be11feb5962fb5e50965d599f7a0103aa8c44786665f86ee0fafdd0af03ed27b7f100cd5e564a5a1a2999bcdc8afd6350a9acf176306be6f013333d419fc013a1b9fce93e0ed00622c1a0d93e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6bb75a20b601514258b204b53eba060dce300706ad43467328c3a284a671b5041717315e2536979a9dceffb110aa287f0571909cfea2966f57dc423bcb7cb543a1c7a2bb6c050df6c5f9b1529a18adec613d1bc7cf4845af07341a2d96a8b1dc0cc4c244aa25fe81b0fc8d63c48b1a46038f54966b9dde6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h487a4bf0acbfa993c7cfc54793e9a0549ed500201c5766388de0d183e2d38820d1f0064c87042bad6646880dfc98a3a51c1bb0157bed457a8c2a55786d11e9024f3d805211a1fb70d64ebe169c15b880dac8d415f78294df8e1f52743fac85b7ce5608ec809b30a79e809310788a63a82285077674dc3d4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8893a6496e16a8fbecbbd26d5f3d3790df312bf6fca8e066d28bfdb51d3a4d671e058f16d19ebdbf0511b443dcf361228e8d828f5f8dea816415179554a2581a8069309c45f7a8c412d1364db08ef4b75add184060449af22b7955954a521d939694e61e27706ba820bde95859790377f4128aadcead5ee3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bec5843c7b04e94b46b6a104e73e519943354f6a0793edee33e1dc8de6d1ddf3c0fc9535f631e3f8bdcb73f96d65e245360e723aa2ebc68edc2b426947011bbd1fd77f7a50d750025de3e941e11d6c487b4fb6b2085ee850303f6b632582e916b0c59681002008a532d472e27d2a3a5f3a0e5a832dfa3ff7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35e30a48211e1505e80cf408f34782a871e834a0647a1908afcdb7fb3632e7b2137283c32df6191c4a5f504626c80481aded77355bd6ecaf9cabf5a37e6c170de67e9c2a0b67d8d83beb0d4c47514b9420e2b5b84e4909ae0e83f4e128d316d91244b8a3e462ae9305d33e3358bb9bf567359d89dce18e5b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbbb711673b5a6168fdbd5e4f195de1cdd451e646e5e9ddc10e0477bcfda2901ee5e969784ce6a7bd075f8905230ab033ddd9549019a7bbb638324cf7f24a719cc00b20c1d71860bbb03a4bb1763f08ecbf336bc09074b3b374f725362ad731d90e1bf48ac5f130a8bd6c3e028746a4525e4ad81c956e0d0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4396869008db03f9e9870b1203753598861920c52a1d54b8bf3caaaa0da6b0dd1737d3afa29780a8f051fc4b3719ce1817722c21110765662495685e04741d0fcae94f4a985193dba812b1b19e368ab372fb5ae039f7f385a0225d68382a099e22cfcb131ad61c49ba781755c0f3f22b665bae1b755db9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dd095f524b30ca072d33221afc4298f89315333adfa224c6be01d813508f491673e7d8e1c4951bc7da6caa617e3532e3d57a401103e124624a784a8e2e3348015d4efe84c0eb5c33e0a64e2fb9a694ea824efbdd410147410401e79266424078d50bb79997f5494f067f485cefe70ce1c2b2b58996bc2633;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f43ef1b05db4eb6f49e9fe1968ebcd0e4978e33d0734ab5c19ad5eb4a49504fa2be5caf82ca29ad9428365beb1c5c0766d176c149f166aee65bcfbcc48fd23d5e7fbabc647aeca8e31c94ba4ea0b3658129aad29badbb4852de4cc13842221ff537a810802ec010b76ee837fb6d2940a7024bc1ad0e0045;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h166ff8fec9188662fad1f83a35aed537a4287eaf571e3f2bd05909359bc5f75c855bd7fc46e183dabf5c243d0224b7e2c6a179de15470a587ff48682393601189f7354168ccb9af143afba822cdfc3645678f2a31c0861d24c601e7aa043ab72aee0149f815cd9ef914b92a39778afa48efef21174d482c20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4bf0590738e625067279b980b5c3806762ddebe58bb70862d31d81e5f1deec4138e375e79274c57a94224fecb4b7922cb0f269ee074eca1b41eac49b36509326192e2779750dd848a2cff2cd50f4a8b31e0133d3ef8cc04d2a0f04a829b3712b3ae2f2c97a078ac5f90e9bfbc532d7da09e3a9814831542b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7209f11e0c7a7b33ef52a2014cd77c62eec2193e813702b7287883c2469de7d77910f01b3699afacdef4402200243c14a6be6aec51fafe6eb48b2a41df7ec20cc97ccf2181d0cbf3db9cb5dc954f08433b1e4e124dbfb5fd6964617b741bf61a55a61513d0622484b3c6cdfbe9514c81662cf9f4554b7f8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h39679b2e7c936a594ab54c1fbf432fbf42b4ba165f0be2c20523b4921b07b7352b62378c179a6adcea4be4c0d6473f2d22f0363515a93fc0e47025a19c69b812d22f4057bc28657a3cd92c856fbbc0a59a2d6fcd916170269536e28d5b551702c221f7bef52d8d3f0286a77d2ed18485508dedf84c3f1de9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eb634c8a8c9f407f18ed65f53cbb52993ae07c86ce9b1248ac1f345101906a5066bfb63089bb893439e9b3fc6e745b442cbf5517e3d8d24747852529a01c9c59fc4d541cbe5c1071606d1edbd2bfae64f52dbb3bfd7c1cc62d2d31ce54f05c7d032fc4530431f4b8c6e28d32536f5632377d42319979fefb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a16fa57fcef6b46f58155f77662359f9122fc5957459dca209e8e1b3036c22a65080f084bc2f79338951096985abd3932921081ccfe408239b08ca167827763dd96f157e759ec054e4fd1bb4a7d11cf56a6fb3337078201fba07e32a26e062a58ae7b70b9ad776040c5227dd3fa5b804010653d769c3534;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb38b5fd9dafc541390fe35959eeca9af16ac3c3c1efb45e5633a0fc71c12c5a45dd0381196f863f863e62e0bb116e8135eadc5decef591d05a704da12f5a0e97f5bc96f8551b072d7099607e50f87032a3548104940a5f8aa33816efa89e3b36622af5bb91931014d6150d0ca78e2bea4b42018e0cd597a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6fc16547a73f6ec17922a86a63188410b6537aa721424f9d04181fa9bf79423fe38e51d22fc9a5bb6d932fda0a73b0e852fd1ba7c1f2a3b5891e93aa59ba166c1522cf1ba55aa99ac188b95281aab6779a40c600618c13a4ad3325e8bd919e6d2bbc5be078b9c525f569e0f69bdc15190e4e4cee4a3efc1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0a75f897b35c5dccd66dcf7d0dbc0250c16c21a8a771354dcd3a4c5221f0748f366491e54559e97eeb485196eb66557307613b14864783bf9b1a17a25794f0a093a09babedea1ed5f2dd2fdf753067700be9bb3ebb624b12e5743c2ee4a3ea1c8900e8433f656edc85bb62925608c15b6ddd71cc676dee4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71f1fa72539ce8e94bc48205b7535ef4bd185954db4d7f76be146d0472812ee4d56921b85a33461137813fe15efe2801c93273305486e00d913fd9676adf51b91c7b1d8f8023d77e2486f3e72d253f96f9b3000a4a38fbfec6cb2e0c5c0aaeea6ebc3abc099f87d976063b6f93fd21df1c172268770c8998;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1944c1c49d33992829bf8dcf9f794ff4f3c683578fab938f199140f683e85186b0287545610d79dd7cf4d548dce081eb3c20c1eb1ab58663c44036b8fed4d94162ee8a2a2295e5d0988c820c940ecdb3d47af70cd456ab9dc6d9934d02abb68ce82147c02861e9ef6485de43fb2dc8b274e8278f9bbc18a3b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1578985b0599718aaa6a4b93944e74ea021e619c317462c4d0bbb98ebc920a4e1a76dcff193b0f7afd81faee6e3fe75ae421fccc8fd650c8ebf63a1b1ffa6a70be04c60fff7d06b168908a073a3c13a35289b418d974ab0b442cdf9b1757adccb9962e7aaf88ece4bd0cea753d510631dcb506e34c52c071;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ae035ac60ddfe7b86c280ab0ca62c319188c1ee7fb17de0c9d83cefd2d955568fee920f00a9d07ffc766cd5356a9890d6a068c40ded35d0b8627762180ed1f93284737318129e2fe739a8c33c23709d31ba5b9422b488774cd12066ab1eee30f4fa1f71af12970bfad259521f9dcebdb1a2e21a093ac75a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a9f03848af78e42fafaa6eb129c5667659f513d6630986e2942a5d8f0d4bd10faa973b1c999370bae468890907df972effd43ec4e48473e74d00d0c31279dbfeb1cc1d54a783d2897d0f9561214656191ae2130d08c388a469b45ea9232f426f31b0a882cbc8b8f8834cda968e91170e4783510dcdd59477;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4f3dcd66cc8b92c7553181fe228a3f6c04820b1c8973c6b361641f1593858816d8cb49de1bbed2ed1709d131357da6c7978785d3bf9617a27d81af960889b503436a7b973f06883bf7f0345322456af3be4c34dfa4946130e82f033f828543f26f9216550c9f085165a9ee3c460ef927a38a89682348dc2f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17107bbf0965394df1526944a5114682284cba064f467ee3d209a37aca8791f82d28e3c32abf495555537cbf6c8b53fb18e0fe28470b3009e093f3e9ce259cfb262f21cb1175bcfa66a2aa763a67b3fadabd93a45caddbd275134b6e13ac90768972f674142628a83d86c749ab7c401a799cb86c331dc4a37;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2ad49d6b5c054fd41a682255a4697b173a8eeb1151a25b1cec0fc40282ea8b8ccde6115ea10f89b39b6512fff35f3b79916909bff111a2e6af000a8c9e9d0e2351a4488cb27b86a59066968a7c1110e2c23e3de5ef64eb11908402ec3de26f388d9110bd50a51d21964ee86f9fd92d66a8f58705e91671c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116426b7acb134a15e5dbdec8980b62ef877e51b3e44d3df294f07d658c95576d3597d37fd216508c8b304172dde972cb4524571480ed7bcc62638763d36326c2df5ba902079ff0c1a2172447e5abcb6b3498f01ba806992995e2d006e0cf2e95c87b7ed4e7fc2d22f60a5384a4b54dcb817666a01df83f89;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc7e7cc674eca7bcc812c4afb05ec15b9e20dd91a8c1537d4c551f63122c2a5229d08686b9d5592ed999b6f49c40a18258ac416e755e2a55fe5ab1cff00a32ece98f2326efe09ed5c990ce7d64ae6668b09c832c8bd7a0cfa43f92fc38ab736e4c7be996a3e195b4556feac01c926bfed9fd0d23f62c4bf91;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181487b8d0c823e9ac3cc4977d2adb26b25f57c172925a9a51f28e08ddfe4388fca12a53f862095aeedfdfd1d6d8bbcd58dc9cadc14ea8f907c1429ad4b11636c5e03ab80f80d109a6fe8829abf7b1222c66754b4f5f5323d1bc5919ef51c81b7024caf8bdb03797ffe0f11eceac0cf906b6f97754ae494c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ebe2dec6b678e1ec73b9a7a3a329fe9d3c4c60d5415f7971b0aeeff36c86e1a2d01327fbc752780cdaa30318fa185cb5465bea4c01047b1a2111cb9529d2f64ac5f8dd69da2bb332c2b5c400c292e05a0e796903708d355b7e7c488b845e44ec3692057e6cf20efd4b472ff7e8ae67e7c0c483bd490f462;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17779cabd14f702350b631a83cfeccc2d1a45154f14dbfb533c9efecbf03726a9e1259474a50d166427119ee5146556605e38649a821bcdcd035461309fafe1b916d45e6fb30e92c73136daf67d690ae41e8ff693a4047663fab093afcf87cda0d005c8737b43793dcdfe4582cfcc38e54e1c3d70b7771908;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd454f70921a4d29380d88c9fed73a7da86b7922350ea62851e07e33514c0491fe526d3b3c8107fb198a4317b69bdb777dbd03be456c68554feee58df12a33381520e2fe2d3e2e7e5ff8fd7c03b35b1534b8c2aa34c14e4a9eb0cdcd415c6c273158587f5b2e79bfed59e577f79c7a9bff5fcf98379c145c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1843982f02f16f241055bd01e912c29cb6d10063232e4bdc031642c646587851be5c77a549d78460136a179543c7937d39a78dedb3c7ff0913a7efb46a1f152698e0bc194effe139e4d4a22fbdd9c7e360a56d3694b53eadeb0eb17bab57a3f99ac1d2da3bd294085e1950d5b1b9177ee9a07d67e1aec4193;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6bd1fc37e502433d948a1d2ffdcf077c860ac770af31c486a2f23d49684d75fbb1a8a8d592882c133d534416a4d4ed47b6348f792d6805363d48c3532b2943398d5b1f5fdd9962478a168e668cdd7c212734ad59868c94f29c56e4a9f28a8980eb8ddb90bff2e11b42346c7beb6b44b639025e748f2a9a04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1921e211d134ed383673ae1fe74bbff280c3b6f1fa9dc0f51e58d70aa31c2aaba52bc6eef994bd886cb9dc8edade7ca13751ac6d10a6b6a8a4f0556d2c41449905d0605027aea575f78b295eb3fc0b5d0df5e7ec441f24ecc354cb72532d79deec2b62eb2a395ddc17f18105fc5d04eabb5fd1a58269a6795;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c64b85ebc0f2acdb86deac8bdd2318922c9069c63ee8f5101c173f80ec8f02fea2d0ee5376bfdcbf8a218f635d1c50b79d92cd8f1764b79e729fa125b5b35993b315cb1f6f66ea5569891b9f36b9355ada05aff0d79cfe4cf303a23148e328bb525eca50c75b45591a840be163f581336fd1e425193da69;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h249dd640275ff48b8c2c7f611f073385fefacfec6ec3bcd573853b14442a0bcd779ce5139417b7740e5d4eae64934dd0d7f4dd3cfe3b5f65dff754c13ee49933d7e3d95a48fac164fe7453c546d24ae469c751eace0615e49fd19307e1f8cf15d2881a19e7f65f49a4acec0ae3f5258e0b015e248fda7c14;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a231defd85c76b4cd9445293a3b5ac148f0eea73208c2e19e37d48ecb61a44552be8d2bd0ba75984f263c567eea12f0dcb32fd8b6a91dd2ebbb27757ac8c6db819f9393a779feaa7e4663f72a8cc703476978ad6be9c30a9a5719a57f1a681e61d881f67bc471ce3f2b9f045df307d058444161a13d474fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d041ed876dddf0fd00b87998b6229c7516dd523a2a9ebc48a13be0c7dcaf7dc3f2f4a3ca3cadc72e13548c1723e724767f130e2f0a462cb98e3d326e927df1c1e707ffaad6d7c21fafa2c71341bc0f8d864da7304f18120e84285dfb6936dc4e2ad2b6ef4e3d2a1579a4ff7a88d570a9d44ffde153dc84ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc6800dfb11fdaa9c8087dbf66c6babebdaf464b6895b42c6e65bf03ac350f98089b8e04efca35888affdc218647c6e5ff44f72c62340c3d1e90af7deed444e98dc836a865ddffc072967fab8ff78dfd4b95ce37aff96b39eaeacfdcae9f5e0a1f300e4f70e386bf3cb81812b420202bc38881a56c509b75;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1415b67f393efae0981d46858639b57e926756554f1cd4b58d2cdcab18d7deb5885a9df810617dc22131215e14321ce6eeaef12bfce639fec76da45e4b87a30c2a39c8255ecafabb77f5e5e0488d06b691aeda426441803ce1369e0d5c8061215f5ffed969fbfce83c75c1df89ae7fb9badf1387d6841f3e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he93000a8d804248702e4a01cd9d60df19b6fb802ca3c62f323395cea7b21bd5c5bfa6284d3b29d2b03bc9aa3e83ba2ebd8e50a64c05445e0c0a1d779e427e472c89cc4f874e3d5a3e83b81df1e9715411647f81baa4692b1d5321d30ce8875fb09ee2e3b515e38248f51f5f62ddfec5e99418bd1c9c97692;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1480acdeb9ead17c6ef6ccbfb8307423e80f74c685365ae9a01050dd86e6137960344e3bbbecd877bb42de7effa5b47d598cfe0a9423084e28cc008fe819c4f620f02d68b571e7c0a993dad01dab2a508b21f908ce35003af9e8dbeb4886b63f078ca9841933a10e8c3476b956d5d7c810ba9a0164fb51fa9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee51ced7a925866f2341519d3589bd3ae201c51fb7bdc9b16cc4cd03ef7fa9bfd65d0a5f085446778b34b47e61e01ea640d68a612e2c56b11edcc2fef4e1592b088c82efccaca57b1f7b602c7e5cb6a16a20b180a7d72d3768a6bcc3cd24308c15603dd46f51187cd79057a100c8f66d120f314eae01c76d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18afd5575d4e13db492398798530acea485773a5ef09909f07b7fb73f540e26198677dfa6ad9eec9e7100c0bb8672fc4d4a6f6160357f86461b661f3363a5ac5bfdb79dea19e85bb59c11d3f241cd8ae960307853bc0fff1e28bf4ea5f365b579370f60efc40c7b3e92ab16b242ef7d3b68326f866079dbf1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5bea443278142a8965213c3abddda2151b334cc35d8cb2496ee8938a2b680df8f3ee6fc8a69457e52eb4bf271f83cc0fac6e60d3eeef4b1e942511b9197515c2f00d96777ff3d353b6b5c4d6bacda699d7d83adf59ce8f6a97719346d2537c6605bfd4964b917ece816aef77e7e148dee7e3a7aa7b4adf9c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha9b65d88a47971ca45a11d900ec4929bf16063fea910fc4a0865edc4ce45f13aa149e4a77a50cfe24786f872552cfc667409b40e57fec1602c0522d1e82556b8d19448a26541d18cc6aade2e2311c9bfdfb86012f5c841ac376fc85b968fbd0190567f1f32798001ff642f0ddc344f8144edff4ea801405d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128d2cb63952a4f3a445ab721ae29c2b9386b896009566706be906921ff38a160421e00766964374996265b2efcb73409bab2e0a0991b26510e7f2747aaa7cc67bcf29515b168d619d13b320232629e51f442e323e7acadd15ab33686759759b415f19a0aca3a1d8679498c731e1412fb6ffdf98598f12329;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1494186f83e8e524f82767bc0747da4b58ac9bac0d4d64ee6614b5b9f5abd0db57c91ae2ffbe55829bdc8f7d798e535147f53e19ff69bccbadcd798b039708e4560eed0fa64bfa8c764bad8145c6455a2df3ab4bedcd5061e045091ec50a336d45a0288c6bc38648c47ad4ad37c20713f9e98e1976a9f3fe9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a515676bc7cc5b3e95b2bbd22aa31ec85c63faa71662cf851bb9c54090d0e4316adeef6f7c6aa91516152982b5b5147b7b72a6e72dac2fb0d58308dc2d8fa3e1dbaa28d3896717b5a2c07c1177b406975ce20b1a6cb74b32ee989d553b0bee6b536b93b8c3494b82214e1570f71e3477664f2e36b12d7cb6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12bd4448a9da0939a5ac60a4c0ac6d5a9ed827c5b9bca98f31b2b93649fa843091c243f16a5327d8dfd28c894178d2f4599123327b607f09903e507394398f45bfd62e490f4e3d9b8d53c479a102db6581c1a5590ea64f474bf529493ef4b7703fd3edf8d5c3b41944efdacdcda1351ea83810012dfbbda29;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5e7f79afbe15cbe93ce8f69a9f5f7f892e13c45a8f33762d99f6ccbf2d97b67abdc7b9c7c972a29abf1605e63ba8261e2f7a23654d132987dac98e8641d8816207739d6c99fe557638660a436b2746c4576c586f75e4155fb14f2700098147737c836d8ede9c8d4247a5748523ddb523f7432df60d546c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a0283c83bb2553a2f0f825daf91a7d8a0a5fa96b89fb98ca510b337b3661fbe91f3ff01a60a002b903ed34dff99b1da9b0642a28346b8bc9f770fcb2016184a306ec43981b85a81b448365f0b683b65226b0cf47ba4b024fc472e3f1f22e202df7575885d7cb13d9ea99a81080bdd9268e43df3c17bf2cd1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6202785d156479dbf3c94c9cc1d103a00691508a91e8b212dfbeed03aaac86f9b37151a30a18c09667ecca2e0ea63bfdd33fe4e2c949dbeb2a0e024fbf4b1fa013bd28bf5e0bdc1ba98f1a561a6a1fe77f49e7a495c29b078f877653c0aff67a153fbf6c2baf1d95a72c3f6618a4c2a70ffd92849cf79cec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79a9b00cd43251eba97bbe4240184530d9c7ddf20e987de5fbcf4017fb21963f9d3fd3460a146fc8437b45ad966f547bff646f16035611360f8da83f48cbee67c1b6df446d7e2fb56e05e8227176d625506c6cb40ae421925abfbfeda73d8a1bcb9a3bc0c2a5c22594656f6a4d0ba905e485e040b672364b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he837d0fd2d66633926de27e0d90dd8b9123a386a656f5abdaf02b62fa2a5e082e4a47a2d7aa920aaebc92e2f601ac78d8222e1c3f024d45558e2bc20d281c0a3a29accc6d64cc58452caf31056d9507e2e4d586367c01526fd64af814a377c91b1b9b8d92a4d79946ce66ea67fd0695c388a0d9e4927c67b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1320972b2f0cf6d04e03f78c130a11f7aa1f6123fc32784e211cc35bfab777da739d491aac7a45a4967eb275842d96b74a2dfe1fe937a429bfa4124a15f0dd9215a4dfc5cfa183e4fc3eae28451b102b199777acd0304edd0f6b7ce1e3a2d90af398d65d10b3df5bc5338ad1157f4d11b0bdfbc62b8ef37a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha266b2a45dc4fcbfbfafcdfea56e4ee725f9aca65b4c6b9242766255dd81d723f23fb56fb3e488cd2bbd91bb4eb6962a780f08fbada64c78b3f2aefdf4ad103ebfd84f4be0d4057ff70aa21a2c41f07efd412284ce2b5cd7566a6a1582d979c780139bc056260f1d93e819fa63f475ca37a138de0ae73242;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b7a609a119abb01c24fdd67a7ff5231a074f599eb8216c88f8c740f9079c2d4ad4346edfd0a3acf4fe64dc0ac188846fc3e7fb3330f35e8e32c8b6bbe7dacf4ff96700a947914f6564a64919d58ee12363f98033e39928b38ac2b35a758813bbb8108a4197af1cc63bc97fc6ca1e69a4ac7a79f0930ca65;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c48e5e3c12e6083ed74f97fba90cc8436896c414e79ad4f3dae1bbf8b1405de4fb6e5ad86d1d8b8503bcf3e6e97e5a15d56cbf73c0d91a001bd168cc1f216b479c80e2078f1c89d1578dd0db5fc26b9be0f35f1f12e0efa75c3c4247c0bf9953387251813f9c2a824de42420fe2177059cdf87d8c7bdb393;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f03c58be99c320540eceb15f2d4ecbc25ec1cec7e2964d610c009e4a72ad83ae16c98b557cfd5d88b8fd05c82c1898bbbfca72896ce8064b5ffcead33de7fbc6d93b732e8d9af1a32b3f0241789ae89fbbfae652b8d72c02298c71049cfb36f8c0617f54c237afe8f97777257a9edfc53e8ccd03dc6447ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b3b901d9e0965d5d57df39ed35359890c8b2762fb15ab982aae204c6605c18a6b09b7a2dcf1ea67688d3733b08d84408d5257ba5417ea894a854020babfb92e68813184567a09972d4609cd1780ded952e3f09e487db870a3c955b6b9f58c0bd47de03b754caf5b5a5f3cd1352f3f5ab6d3426b5759e10b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c1f45af58a94b3878a558ac6a664ed57a8ea822136cbbb43e819fcb41e2ab765baaf57148cc44b4f0f92a0dcc42782f5af8067b6f85edfa15a579b694c7bd0a8baf9c8e64cd960998469d6f676db43ef2726967a42899cef3c6c69d0678fa236522aa177436fc07b0f881f4e577cd4366cdda57c70497f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12899d294e49e1fc1a16dcbd9d9e11a8d829c020bdf95137d9a7d9ccca1c4d33541ddf6817ca785c0194f6ce01761bee1f7bd998758382a173ddc1f0816965f8a04ac50ffce278203a6194741d9cfd068214b7c5df6268bcf988b7895320b72cc59bfaf9c67f61dc61d03225cab9252fd9d6651f0cd7caf3b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ffc7220d9c73a50b370fc4f973bed63af1fb87b995851e5d0676867d11905f776d15c2280cd44eb54018f31d552359fa95eaa76dad169969ca59be97f66a4ad5d2c4e2615a3db40fe0d3006dedb62d9fa15c4b4103a13ffa8c67d4f24c926b34af11a4e73fb07da063e5ab891f3d28b01ef02afd556df49;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a554b6e970648832b4ba2580bf25103add764c457a86a3930a81e56675735ae7cef87fd4c247d48158cd676168d070f4f69b4a0f786edd9e317ef0b19ce2a22eec25f5ace119291b333a79975406f82e279a35b16ad104a93295e125b243320c7926009c9cb340baf62b6e6616415f34c57f4ce5ba67056;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hff579c330d97862642aa49fc33191a854a44318a6afd248d8b171c20fc153b80989d31e97c9f6f03a618298bbc00e2c83c25b0c0deb389a75da617b52fb54dffb111e66fa800a35208b31ba4aa5d1c744200da211dfd6ddb52ac48e0d3d163c67f990b86d22f7ccec98fdcaf8d39c063ca2a441a125faea5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4882913f4df4c93de88a715ec9a9eaf707d17ed1917064b694003feb4f491bef8e212dad58f69b45cc483d762023fb600b88ece9ce6eb76463fdf0f930164f60e3a1567d00e28840bbc883e4a14d954013bee340b55077c4d6e70c16f4cdfdf840ffae9365817d92c9275a85d3c8892ba7a390f3a0d5b2f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h191ae7e0bf89ab121301c1a7cba6ca04e2d02800cc41840e67aa6032503d338f38e214038b04b32efc60a8caf7c6ba299048888ea5162798e863b661797aa715e88b3e93d44aaa023efd29fcd5f1685f633bb869cba43850b4078548e1e7acdfa3c6b83f41c29f28950a2b66972943666653f04dcd9e7519c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d585d4dd1b50f5b70c0f1d4b4910bed824f7a8015fb752dce265f3318c57a64056097a7538fd05d9a0d2bce27a7cf2ace0fc99dbbff63715cdc8b2ab00a68e86888cb434a43de2ee2584b6196598d667bf7acd6b255ac51ce251cedf5b55a9f1e88761b21e56c832210bd119667f1694f22530d12551e6ce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7df107bf64ee687364a89d86f1456154879505269e2f3f179f20067926358634e7f4781a320db267d23e4de65322e7587e30ada37fb623f401cf45d271975cd930c965220ad791b6ac79abbb1422706859b5080f48c7c70cd18e3d6dbd4ef2a6588d686163d2d9c068d31e61a19ff0674f3f2952f862768d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d504dccae68d9cb83663cc7f1d216a70c0a8593a29f27efab102d448cb1e573566e1bb77bc10ad7d236b8c847a65a0737275276b7dbf4539cb0c3e4d141100dc307706b3570248dd96c702b6be981578d688f9ef290d57f95c36a3f39594cff038d982b5103430f6ddd438e3d133c09107eb34cefb4671d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2e2c479aafd0e36d14fcdaab15309bc1ef1808af7c84edb8996aeaed6ad54f3405e1e261c42284e62b7e1614282af7ed7c2a15a9c68dfe22be89ab07a00dfa9e3ffb5533af70beb804bab6430a19d464ddc6cdca672736a70f9879952d5918af44642de78f9b88d46d864fe9edeffbe0d717504af80cf3c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47e3498a809759117608b76a7eeb919308dea55532a91a39aca8a18cc2fa8d0dea4a657c69b58bac0023966ffea590e0ec5cd4ff909cbc84c3a27319b01b8c3fddcb1a61eb6cbc9ed58fa51687eff92e44cf4f137ec030af279ef6a404d47fcfe59a546252cde04fa1fc2ac26cd386019234800576323300;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha568eddd64d69bf311725d2a9109d5003b5665c19c35fdebe6423f6a365188fd732184bb7ed1c357db5c276cf51ae25666a683a1eac5e5008831e0156091314c35a06e9406863847c493fce39ca9865d3ef7f665834387f5ac123b688d6429f4799afc9b1ca0c61e3d24034c3b3bc9150f61003bd5754619;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e95f04032760416b0f4839d7a1f7e7ec11f6065bf12b3695bcc534925d0d40b3242a8273b28df706fbf983989298e5ffe26eabcd7b035c151e099923dbfdbb21dc93d412ccd69479e34f670b2340dec7974db067d620ae9e25f547d8083084927cb350ff1e1149b90143b59e4342030dc9015626b547cda;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2111904292c34ae914feb378c4f1b3ba1895025abdef7e1750f37d00dba535abc4df3b48ff87a593fae610244ac243c6df9061a08bab08b3ad29c6cbf9078d9af9ccdf71e7810e76c6e0c3fa845ecfa0c75e2b8b78144951b97c8d101f687ced812d01d29fd5cd8bf0109c3b571f1d706cf020429ffd2aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f17ad364c1f8816e360190425c7ec070c6a07959a7942926525780122accddf9da998f82550591aabae38ee25b1cc732c414ee02b7bcca199897d31c16a9a8f34a56c4046872db7751653e3cdb0c2494dc0cc2d57d340f0958bf8ef8106e6bdea91b4f632dc269f22fea9cb0bb7a35cfb43017452659ede;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h45d4034924e66bd8ae83c45d4d785c9325d2282f37b84f19be83c7e08c1f55b53c7fccf0bbd8c76786d28a4978df7407568db0d77a14e133723f182f806a2b9974e2bceb14ff7b1418c0176b38db962a0fb721df8f0c7ecaa14505c5334bd4308584fee5b3634b9e6c34eb499852cd2fbcc274a0fff7cc51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1341772166e6cb1c60f960a74017a8c94e31279dfae312dca507ec6f1ac04e6e87699c6858f26d8539f5c21ca09b2456eec948cc08786e699bc630885ae430662d1f56e8067b6666f23234230e56154f9835b982e362fc7c97303f096d54c59dd3bc9cd4419f06b1f2568c6502830cc8959d787bc97d731fc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfe86ee5d0d946e9f009d40abd95059bf314de9336814c649894b8a5f257b5cfcc9cb7d8ece6a261f18b555549fcbd5cf13b8ba173374a57c12b1d5dc1bb4505242f4bf714c9806ebab7f99949f444796121c70a26e15647426f99f1a342c65ef738fd2369f83807a3c9b181416a0eaa86acd71dff2825e27;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h45310ceb94ed58fb093104b93415e73d834405e3cd7c5b10e106f76b82cc4821a1a9b0de792af153e4a339b002fea82f3290594eb85212255c8199c0628698f37ae73f7acece466b5a9863b45fb704dd8298aae940bfd78a4b8e347b1a973168406d42ee09941522e963e0f15b496d314d022e46e9f4b889;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hca7d6848127544f0cf2f41837d87fde6162718bbd229bea41d1c93f09d37893c0e59b9597740835b3b0ca750fdc5e89eeb40fb3456fc8a7ebe5d29f39883346546d6098973a108543b71b4e8d3122ab050f3ba193045474fb05b6123cc5d641f1a60710a7c3c239d74c4d1d58c39903435e215db5185c9b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h43610c2301c751a398fdf1f108dcac9567e181314d80b6251596c6ee2f1ace0b702d72dd6153fc6f76405b7f58337af5b0917972f722f04163a4abd214b7a0bf633b03d44d58a76dd511e7dcfe086233df86b879fe366f6627c5f1e0e52d856b69f884a22045d81d1277e04314f40cc24add357a276cfb40;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5cb25242b13cb9c2d348126e20c84af690f40e1d46caa2027edf1d281652889e2276f53560cb1ad4767c466fce935f47fe7f90c1bd62ae77cdf381d3e358085082387dad298484b6f4b18705a651c4caac286b95a8ea0c05826cb0d73eb266a8a1d37d50fc0d389d7ca43097078fe56b70e0ab7986c21f98;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h705d8afb666c90fcaee910c14fb54fbe5f1f9cefa2518789c8fb1c15b5e4f147eb815b7d9199295a6c933d043bd3d6b5ee14bae441383cd6ac7879b168dbd534421b807822b47e2e6ce5b1fd13166bd0fcfc7c047294195e45a743e7e56287a37b98ab65a1b52431c1b717218819b908a7fbedb1af8bc8bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6901f58c51b82e1c33d94e93a3050fcde4df0266deba9446af84bf015f9baa9921e62cccb8f3e2b008cfb0d482d35535ef0a3ab83fde7863d02ff3c531dec278b3aceef054e76203eaec15c261aabe8fcaa4042efd73085097ca59e2d02a4744f6b40cb3162f11d60d4094907bffa4d5e30337d9cf7a7434;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15fa416d8147fea8772c24bb767759365bb23a38e1c328948d356b6c5eb6e386192a00dcd9d4403372ee6246435705dd430338dfac76b5b8b39fb1c2350a9e91cfe9c6198e071f1d42c8bc340b149ad88a2e667ea625a350e244b6bc62f4dfb635edf45f30a8ec8aa15e0cb4c410b2eb95f34bb4e08cd3e4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha97d6b74258d3ff2ccd930562571ecc022aa4fa25adac6fad77cad81f74f0f87e876a6b20cdee730041927dab2f5b05b6045f5589d39e47768dc13c4b0ff13b1b812d41e5b4ef5b43fa4c8ed983e9caa9ff1c3e13c397fcbbfea5333867cd113b89d37a830a698983ab49603342b769c473564b9b466671c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1407769b363e849bd5372bfa69e5fc466dbe2d1e2af965d702beeb090ca123680f2c9c24b7bbaf373d60554b985b31f3e02d73b71ed231587c4da425760352bc3f5cdf3bfd7a8d66acc759f77aa84af876d7ce623baecb5769701d80c9852bae7ebd4a3689722554446bc897178ad8718b3fadbc81dc8d02f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd56a13a9435ce8b5d8121c7567282a9e8267c24d39ab27f6c32397c0701d91405d70922768556b42d478538be98e70038598cee19ed823f0849c67c5290e89c53dadb6577c4bc9e3c9c4f4922891729d8592c119bd673bb0db74c86043ae4d1883579203450a8338a8317c3b85c7413d7822b3cdf75058cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2392600252665da75f42fa6ff8e594703603a3ae65d984372fe5268597e783a88384193208227048e8ac80a7eb8cbde60cc9c120c5414b2fbde4f9f1c88ef471bf415ab6e20c26e52b588c436f9ac0e716813a2f20d445907bb8a539da8fcfb1af3afbf7304f725a93df58750ce7dd4ca3699c3081e06b3d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6ddb51b66fffdacfdaf209952336f6d7e70bbaa0a8c548ed7996b4952339af3a3aba6d4ce22ec70e78b21940083de996e5db9362e1a270f3169cf99d521af8f5a466bab68af03617f9e4392eb0b4ab30e28415a254b4fe425d80c09affa2c9c2c46cb6ef19b518be7e47263b0c784fba3970d94ac2ea2349;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8fa442c64292f305d6910e84a2438206c5e9c684b181241d4c6c5631ae0c1f9f50f7e10b17ad5aab14965185d10892156d9b512bdf70ac54cb20fb4b08c5cae1cdfd764ef460c809db495e0b9cf1ce61604654e2e43e40b5a334ea6642e4b0f30850a45d597cf01a7d26adbeb1aaf207dd79a84359bb88bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46f466f083adf8247ef77d8e4718170fb7baec4803b014cb8c947c5d9906363e793fd3260df7df517f7c6defaf1e9fba76149baa86bc473eed3ce2b303f7e228ab444a24cb90a1907ccaea84774a907ec9ea70abe31bc24e62b7a2a4177f258926f4da77ae48119ad25eda2c2c9e6b4eb5e9a112f0923f36;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h371b9afee1ba62aeb1228af8705147ffae9a7599966add971efbe2230c257c23cdd7e764288afe2aa37942212506471a9687836c17d3d2510393c15d00e4838e3c4a887c0eef9b250204eada313ac5180cce0a5a4beec1439f644f1f1dc2f7186858c04543569b907172fad43dbc2a79343420e7f9ee3174;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heecbf07161427642fc5b493774a40c5dde6f77507fb7d1bdcbaaec27f208f690a26b06fe2e5ff55f6c5f7981991ed330bfdb3f8c7931a5c7903e60b5e58120fb89ca0db5064256a0feff43b657a5108316a75d992d755560e2824298186791f98f3d8e8bfc4bbadcfe3ab5db3e72ccf54a869e4f6a50735e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e7353d4d82f26ef5e15bfb48c661cc55a19af3a53c7346a9c7af837080e8d08f53ccdba62fb80272d5021b38b7f9341d08f1a2f15edeeb50ac9208487368a9c3fe7a33ba2666c502f6cd4601a0033865fd5eab14734cdc3d882675da93a099a40be1cb7e730efcfb10023078ff485e988cca187ef3a0d992;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hea7b20f9a58c3e50e1ad161bc5ab3a5df5b67ad5c8fbc8996617d08595548ef9477733344ae22e794a42194ee99025a99e76608bc715a50af47e54d20d1b483d4c19924069fbfaa97afb8ef683dbc6da4233079727fe9749db1da008c92bed156871e1ae250db42ef3abda09a03a09353cdbb849443d5a16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc6416b838e58da5ca925e361704a96f6ee55c4cfd953692a4b7d3b2e8e384f5cc7d3a3e4f5e1cc1eb00fa8e7c1ef81d1469316e2236db02459b0f6e28955e8b09235a70081637c9526c4dc34be0f981dd0daaafdd5ee6b78533149ea5ac77cfc0c41cb78cb8a5c1225c4000f3d2b16565fd7924ff80e250;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha7c00bd5aa85d5610edc52818ebe3bbd6e6334c46f1ab9426c2a8ba5b960f3dca2f7ff1964f1d8ee41e7d6cfeb0b8aea6d07ff9653030ae78859d7451280e53cc96829a6712c35bdcd8165d47f5bfc9c60796e06d88901887eaef7fce4f30e9a67698ca8d512861f742aa89ceaffad64490aef8a43dbff88;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10dbedad7729b3856e5090f38d68fb9d044859e6fdcdb0bf34234659d7233749ab50d71d66cc4524bf107773b16a84f71c029b3817b03c976b44be8befbfd23dafb89c383cf4108282acc239ce10aa38ac0d85ed4b2cd17a8a5fe95c2906484cf6fc42eca261ec0fa5e45c99fc97bdebf4ade9c5e4ca92bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13475f943bd3219322a494e0b04702f14487ad3ce91a839b11bca6a0a575242e691965ed42c9e775d69027430450baee5c5d7d816cd7e306af7f9f547ada855579b87bff84135959d7fea85cf674efa341bb21a3e10ccef5f453ed8ffdeaead900b0686c9634891c63dc56adc0fa04b6ff98e9e2bf6530b04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a016d4685998810197a8035d72938c47ced1a3f0b109feba13f8be18816b8391b3d934026e4f5cfde1263fb51b5dbad8f20fd7690751e520aac6fa48838257ce3b359f4afcbb09257e999383894354966fc427a4529c1ae573022cae0027aec834e8c425072f94b025c9606b14cb071e59faa1a72b8d8b36;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h135ef02eee6aaf8256e21206186ca2ae57ebad4d7f321df9ed1278452f5624624029350e99d4e7b7f73d93a55e3cd20b8974187148de0aa56630ec10a90452e0570180b73514ffda7cdd7496d27dacb87cdaa8662518b15d44ad08d5f45c504c954992c331cf3ecb493a75464addd3187b92841bb4ed3f9ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3ace7813d9534656f77d93365fd6c05fd52c1ea6da0d132ca6b8db44423c495bfc9c49d080c56e493678e3d06c7c1afe9c23ec15facb13ccb290af64a188332c7f583f5f50c50b35cfaaa21816900aea75229853ce9b74798cef64c75069cc27b1daf6e832f320778746d44460cd49f7e03ad8555ceef01;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16a47179c3e32c2cd43f0aaa5c069a20e79a90ef0eb015d209382891b53369fb9c55901f636a6d5e11040e2b2ff4827f7766ecb148a0026aee9d6f7f7ae0ba418e07697c85fc5e06e1f8f841a758252bc5ec46e39bce25ff67f71537bb8760f41be272e6f54f3459750c72799dda8ed9447494bca1b88cc26;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h96788d310df5d2b9e73b206f057eb46d3643f1c6d1c42d398ef958a9cef27d70931a23cec467752814b55e2a0f460200a79ff3a41eb8dccec61f97eb754707380ae3b267312a584c9749621007c5cc5c1727344669a150ff2df478022f586f769104db3e4e14a47d5015982407154d0b9396c7975fb0db3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h55421ba95ba8945a09c0206c372e782cb2f008a17187cf8606ada05e2a8c581aeff333eaa7fbd560e3079aeeb16e3933873ab414741bad7924903820ceb96e68a60c3574e7fad904eafed735ea4f2af04019e1aaf4544a869934334ca90bad2b9e2af27e661668f562dff6afb1bbadaec1347695e1c2be06;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16685c14017cb3e1f8d3e2778c36b50c9dff3d39057eb28d239449a7050b871f7bf672449b39541447462aba6d15b71181f3faa2e4a63b86a35a130431959b7d204be8401ec1c43c48734b26ee6d0cefda8ad4625e2e9303ce1b72bd6100822af600231a652b9e032bf23126b6e1f90c6074feb1d8854a0a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd23ee549bce4dab37396103760a55beed81ad35ce7d2e4072cbf29923df0fabb5425e3493656a3ca7d397e72216d04342abed7ad1a3085ffd9e92ce098a26c4f94af847f83b543ad40b729aacb887a84e01b09357139f1c9f2dd72a5624b7153046b744bbc8709b2a39a4aef333387537216548d70083ad5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1809ebd4b46bdc7b4ee6c77887af9a7b7ca0cd15ad5ae05e8f3609e7e1b47fe9efbbdd4f3b2ed1f58d671b4024f7835d110cca415d807ab9eeb075fa1f68acede22ee55c04e518af233b42d4b78eb1ee7c7bcf297634802eac740da7d7d43b50acdb5581682612759eb5f1675e538da0bdcc36858d7986e30;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1519a1e01902c47e5724bed44a4f8994e1e930be41bef62c4d3ce6df55bebde1dcf87a090e4da379f76b076b3fa426874186b2bb30a6df9842135e11566c11263aa489ae555ece6412c1e59c0f90915afbb85d3ebebfb876597e1a73a73ed8353e13c8dd98cfca820cdbbf098fb1540c5e9bcecf9ef76330c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13935bb6629df0bf7cb1f287955cf7a3953729788f25385031b0aedc178720097cd2f9d9b94d16c6f1133993a1db698e293ef23a4c57e1efabb33989932c3c8d31a3615ef2594b24c6c69717421d386daf2b784844f49c2d94d12f11532f0797691f09a3168834a6cb333c84bcba63de721f353e94deb0809;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a6518ee27c7531088003866403327ebeca5f2734c84817ac2426e8773bb1461379bb182789a8f634947d8e906f442c13ec2879526cb42772b645dcbfe7e65d87a05fb1167ce9b8e8e8e74932b9aaac2ab01428cd137984149b433c145fc2c7f4c2dce3fc00c093a74d7e7d908eb1b9ca545aca36a70300;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8d5ec8a0bbf95c8e52aad911b36964a2b16e7aa3d97a1ba537aa89205bc217531f76c677dbed4a0116bbe438fff7f37c676d4874a88ecf7d94e00be6e95ca34f3a7d42f62077e09968c4fbebfc67d1d1915fb143181d3e2504b275b25a2d69edc2a5f7852bef987fbf4ed5363aff37a11712806f31d0d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h150992e54c277fd7b2099122285ca20877507279c22099317788fd7bb809673f69e1ea463260cf11392f375386a8f2feabf47da326a62b0fada61f8555460e9338b7f3b9e76b189e3c6800a55722204ed06cbb55397d54e4929d09d5a5d4572f2c06dbb9509a489b51eaa77fbbee07b508c4ddac105d09acc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hca23a38bc9ea91f83e2c3c55568f588d70afac96d7c0d35d44ddb4e31bef8496a53caa56defc590dfbd203be1ab9f58401e4e4d669a96b5913e87475f20e1673a9d06d28c1dda6f42fe6deb8366f3a3117d248732189791f8bfb91a26abd78fdab40f275c85e8511b01f84e511dbef27a4e3727ef7e83fe6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc6ff17c3959f6d058e34ebf7cadf4c2180874def4cfa6c2bcdc58a9b2cb613e9f9f58b1bd6dde888b1a6f1e52600dd5d60ca4d7891dbf603d764ef8862a84c2aec22234265561161db3634e83d0d83c3bd944f4c5d9dd26d52c9cce66c829344b32ea025a5cb784d6febe4a489558ad39e09729a4631210;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h139eb18c42de74de6e2ec80791c04b310947026b0e1cf991ed945da9f8bcd249dc0a84bb4a7afe3173b3924a9df7e858cef882eb02b1a34eb2b044b3aafb3042b8d1558811e67cb534a105efff99358bf661ed9d87c354000e6892e6608120b6da6091f4cadb0945af4d68b2740105020818d8357963f90fc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h417f0594a69f9a605b6a811af384e21e519fc212bf73f6357188e34263185534afc5b9f5bf7a078e2460e976cd912dbb272c8e708b7bb46e642be23194e32492796e8dad48be8e849b9ca36cb1279241e9eea63effeae4072551ecf91a5bdfadd00c072082275cf6ac0951022042aa4672d4d4305e97e45;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbbe7bd6d60f30a931a07d7aaa88c4f9828b6e3523e18a0c0cf11f337167de33fb7fdbd2d2f6dd5957a7e4008912bb0803c348636f14658c7f46b993ce91c24a887c2a5c902fdd06190261eb635498813ec1a386fb7f37974efe68932be2d03cd8dd6eed0ae49729be35749ae4e1daca7daceafa5a15dcd1f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1db9d92ba22db766f9da2a4874da009b4927b35d48e89e23f49f38f201e78818c22703995325178be5cf942b04e7ea074c63f254b355a3d793a23d601c1eb924da47dcfce5f6e35caa1bdaacaf5be3b5de6996f94c06bd5574551454016550233548b5b17f35acc7f5d92bca0e8e1c1fd4b5b51e0f0221f4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7e10c09309afd415b5db7e649c2d49a978d6633602bdbd9335316a68c3f2f6b116cbfccfbdbd236bd571e02c0e73a37d61949791383e0ec82a8bbae332a6044286de46ae615ede67389d1dd8eadb821cb71e1ba7a11f69f89859ceac7de44ce72eac906ea85db8737dc8066919c2f62c657499ce6451de22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a0581c41d0222075da140e4095b3b1cdee58f53e27b3759da637d4182f4313c87f1aa90d419747fced33fc31af132eee7eca65556dcd5249a4d8c26a21b777f0225c8da9f6dd703237a03d27ee85c4a6845f3686113cc65a3616adc2b5b59eab900cb71ad5f07c4dca78079d1a4339b2893cde8da367dc59;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h54ec18c675eabcceaae29b8938e216f7ca336c1d3c4c725702f88b76954a10a57b07c8ed6a7b0c0b5e88b2523b163200daae4ed3a9eced09ea5c2f863b799724211b68940e2bb2d6a86cb4938e1f942d62d0ee8f28cc46f946765023c44d007c8b97ca92c37876b16e93ec2272413c3dcde0a7a966555396;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193f34197b0e4543e1f2ed401dc2ddeb5e908a2d17d1db269088d6702f740ec3a17d2c40ce9b8c4dd3227eecb0411da182fbeb49b36cfda85e85172c9bcdec24cfb06f5b39b7ea5834477db0ccf29e63b8e5685bd97f6e555e1e868c4dc65e73afc955fd2581919470261fdaab27e9d166a24d119337398f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha20cc1f66629ee04b494ef7c439c633e4e22305c4190aa37880f41a5282587c205de78afaf18f5da8baaa7a3c37c5dfcf170a0e9f726bd2429e787dd7d010e746740ee641733412bdb8c4239a4de7cc3b0ea5a17eaac90ab89eb45e49a7d03bd5419e14343fcd710abf19ff36c2232570aad1bd52edc44c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d44ada11c388020d9597ce87914d269fcc53a1711b458714a714d51196c746d540b1e3b9ca7cd921e38718fab96ee52ad9660c155ea5266564196f47880d7908227252ae8ab1582d9e329e2c7928e11fff8f28c87b0010366497fcf81edb1789ac1f7c0680b93f77d926bbd4dacd933a0fe57dc0b534ae1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8eb12913d58de8897749d23b292f8ebd7a5a44d263b3bc35b730a37574b3dfbd6610c6565e7501480e487270c96154b889426343740c3d1576662771e46d4b990c06d1ca8635f091311cdc96452cadcb8b058984ab9ad330659659f5813806605b9b170ced61546a5b90513e984abf1cb6695028a4bd34e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1478fa9bbd5580aff6309240b300aa3e03ca1869a2289822b1d84dc54b0d7c70ba6c79f370462a9834717c34661e1251cef3ce47181d0f99f9970df4825207dac4d96d1040d77416a46a77498fd6e2fc45c9281b3e09e72649f41693369f151d9a561fe33dc1a18458a8cd76430b8ab5278999e5c28e39405;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h97ae7b145b12afd67f3c8a7b3f30d8bf638ca54e108af037e2c88c238486e39d128a493e83fa7c73e960e1bc05812a4b822bf8b60020d990cec19591b4b974e22f9a5b829c75218d86c0a701fe4972aacd7cd414e54d7cae731991fd19d08d96818427e1bccf0496b9a862b11bc8eae0eb4111ab7a406533;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2983869e0a8a54c9a72645a17c931613f3e2a070b13855b768206c79670337ce83fee7b6c87f213bf4e48c4a5dbabc2be7f826ab3f0ed528c3529426efde973249104c5318b9ec2b914648162b6e4e59266c798cc86503a6da8993f6b7ced65cadf46fc73ac880df97e191106b53758de8338fed3be3d23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h169437e9f4a900468b0018866dbc5bb3f7ac77a5b0a562710cc7cfff1d8838b5cf708a89195fadd9974ae8518c3186a95d7b2759e6252a9c2cf2c6437ba552ab2ed6cef7a200206223f37d490c77cd104983344ebdfd94a429a23a1a57ed44f810c956ddf941151cdfb8b2215c79639df9d2c05294e43dcd2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf264e6bb55d25b5d39077291f8187f4348f51e460861daecc0509dd7468af2d2dfbe95283b8b3f3e0b15f4abf00560e9fa12787f5c02647a1fadd5683bfca3daa8ed1760035202374f8acd20b5d6a569554f85eb190b619f6192aca4c13944aeec0ca8414ff3fe67a870172f3d685b6edaf5d583361cecb3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17100865113ad5ebda8f0c448ee12511bec822a17d964080237cd6ec408119ac5684bd220477dd67756cbebd3d85c76d86ddd80f27262fd94365ba535e2e1052bf870f2d107c6faca67c0a24b13cc2abea40cd5f283803ad7896906cb27db75944a4cc4e7837768e1cd34f13bbe9d0f0b3a416bf30654be34;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b739343a9c30963a42744ad9c13b8715c9e61c541ef415d46fe5a411a9de67503281400452df7d3cd8c43967171e609434eaafc6000c51b74cd1f336b4760f1f7481cfb8c0dcc6e4886598615a2dd982c49f651448c38108cb86683b5b2e26aa3d1ee7c71ea95792769f17f6719737397bb42a8e6c7641bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h103da014e5223a39da8f90a08401d250880fc6cd72946b7cd8aaf589ad3280f6160e0b0b12bb7e85f3e046e088bf03dfbe893f7115c2707a8be062729e381e79ff3491ff3aa0362cfba47dc96017fb11f8070070c428287a4f7ef9e1edc2bedb4b7aeb6c733ef3a37597db2c2c0beade8c2ffdde84f91bc4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha32e37d16f81b078faccf2ad057dc4a47cc33b1d96cb2d6b27fe55685e3d49e517ee7318e48e041ede1b199c2d20398adf9f3e4854b03893406a8458e248d552aa7526ec3882757f03d63dad6efbf2eaf1e8e5251b56ebe4e1c311038f7d87e403815565af9643a98681041eecde9490654dcfeaf9d29edd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb2e32d389d7d7c0827caae15fb9c3d797a45ce12e3aea502e83a133284e08e13a29f0b900f90ca9f2593396b3c2054d9f5ed7e8f51c4ec9b75bec8cc4e11591cf21e7c87bd9fe799e7b832fe13ee400007f5c7da3e3c23fc7cfed12e85e88ec950091a51ae784f707dd4d4e2f888d2396b308bf74889951e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf22f01e384c0f4e4bc12182c32cdecc817ac9242b1a3c658a5b2d63478897a4ee51a608351ff0d5b18fb8b4ed1ce1b8aaa181952ed01b1bbb494a2ac17f3897b7a45e87943c82f1964ec173fdb816ab37c22157eef243b92d2df68e7d016b284444022feb6b73c66445576b58ea1444e19d2ef5374d00d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b7cc2c98422e8a10a6463073ac55067075fe3122faf229bf2682555c1cd195ea4225ea63fc22d403895acf3cbad9fa0d4de5ec3188810a2244f7c8638fde402a004cfd6b1252e5b8cbc8f1aaa900355876b824bcb005b8c6676c7273f5b2e164d7cd741dd843fab9862435771e4fc0e356fdb25c3687af06;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb54912c22a28c7ce814b04a1d06919b1d70fdc59a03f03e01d18356dedaa7ee2ab54529e9824ac6a2142d91d805c46a02b57d422aca5eb11d4d244cb93ae6bcb0c4a64f7fd21033567b52d39d480181e5d6fab6cbba7e6109e648e4ed2bd1e34b8c339c2bf5faee4969c658618f221680c3633f976004af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6cffd6d9c45f16240c2c0cfee7eae30da32d2521ed3f03d492398c017a56dd4a43ef9ee83d9ed595ea3204435077b58871cf3fbb8de3d6da74865437a4b015a29a724be15d1abee79e678c1b7ee617ffbe14d1f9cdb86319ebe12d1604d22358c1b77d25ffcb58dd451789f452b3e1568eb2a83920898cc9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de75506abb258cba399b656e6f89fa1bf775c90d3fa0dfbe77b8a7641a4df5d213381cb1d07969a7f6ca991b0b863db8809d5c961edaf11325d08e1627809bbc17edb8a595fe812cb1b7205549d1cef660bb7c1ed0dcf91b3b53642054f63a6ee63cfb5e2aa62775ed516e5d768642e78f82992c25f11602;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hed5be05ffe742e1a36bcd0c3bd4006a9d113743b136bd0cd8dccc5da4b4aa94ad6af7ac7a80baec6d00b2eb19b5faa31b3ffe11864f14c7617258c95266d7fa9617d73c13e344d06cc2d98455286d30bcd36c66019d836fce286156b17f3f308e0e6c2fc2618396ef523fc661969ecef2792fc2db849bb8b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e83f9d8112c28c81696bf3f39ad7cb97f74a0160b45b3ca1b52cab954a3c542ae8bbdfd3eb9a241bf572888d3328856080d0f295a4507ba5620873084439740518c3273aa86d450a86bdbf84ebab3b676b542b6dc96810da26b208fe3bf51a00d8a28f10c7aa1ecd8b5ac27dfc7f6887ce61d82b34d21b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12720908ca0d2fbb22e8f3e0ceecf9089414d8a380b2d7edd1c40ffd1897f894dbb6cd5ed2f501037ceb91581c8cfece8dce543778893e9097fdd3fa5ca0e96336bbcf800d41e961a79449bf6f6dc5184e654e0db41eab22489a663fd9fbaf2d0f7ae98b1957e99dd14ee4936b97f3227f47cf6c7ce65bcd0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8e2d853e099f7a1a8691d0f785a2df7dc27fcb7eb54a87d0e7a772563fa8e6500898d78dc15c427f354e6dc67d74fbc08665003bf49d304283a892cdd8a90fcee7ca6ec7c59d133bcadb933b825346e61b9779d5a9d696d962de59d071711c7f941f88f348a6c76f7654e30acc31481d19c3544d72af34e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5ee150a9459589ea8893a5ef93b3241e8c498a690d0c2972a18773acd7272f4753b2f563018dbe93f3836f640a692c9c833320a4211cdb6b72272f0e23d3272077158cc3ca75fa7b855999857cda501bdb9f3abc8b27e4f9e83ca70dd9695d8c95d7e6e18848a210dc4258f21d129e05051d8bf44710296;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h40a241b6357199fbc3682e6170cfd7a2bf85effaedebf3ad61cda42a6d8c3a39ed256f5d73dd0431da2bbd4f92161cd1b7f144c4883c2b77cb56e270d6dddd35ebd530148bcdfc197e83d5103f5f785854c0d69f25c446aadf53021ce88bcc5a7f82520e76467a696ec03537c9973344be12393caf0db9f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9bb3970ec551c0d35b6f7960c8909602acc3c6b7742b72a3d428a8840ac30fb827e1a88db2ef72165bccb47e9d7cfab4af66110d592a706fae90fdaa645505e0209d6f975ec228e6c3e77ccf01933eef2eba50e93af1764a7abd5c6af63656e7e61de59761b6d5a2ec4dab8e3308563daaf5e2bc4ab8f11f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f9c774a3579221bfc357e81335eac59a66c23dc2cfb6a6228c353d98a5eab383e588d32e69b11bff0145937e86eb19e457689b2861a693bef4bab2e303ebfbd833281c5d96fed820825f1e48466c7936c7994fcda2c17f97c44105e70d41652da973de560ed421730c81d5ff20763682ec9d8d5772a7a38;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'habe8bf7e2e18470ecf964e48e19798925b2cc013e7f602ffdb7b8d5230d5d3e61800da612122dfeb56d26e2adea5b5b2c46680e7650f30d1d6561f45bb4efd8604f93c484f108c481904e57c76e8530321354e98f7faa204e7830ff47c11e1cac0ba2cc5c8ffc677b811e44d136f9616844527b5f64349ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1871e70befb6350cd16187caced9c96b035d349ee44dc41d4be8f19691f16dab47b1600f4e8bf15d8e91580d107f3665ea7cc718587ea76eac3687750acac79aa3634e95eab7c9c1690502b849958272fcabe6ba9b7c667ef6efc00f7d82a92830aac69f57020ce6672275c1b102f121ce9a240b253421e78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1051166c3d703a2981c2cce6ab6c83d8d815d1563f5a49f713042d0f1dbcb29f506d44deb46e2e87ba24e6a854b76c6e9b134927fd7897ec74bcf4d882c59f5df908aad68863a930d8268f98b814c1c98a137c2dc5b170b4c24f76f9496566bcc1208944e2c31e38cc815b293e5ead22ad02ac4be2c4a0e72;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hccc4944242983f46dd8c907d7a2f0d4ac2e5a28a74429c7b1ccf76a8d48d79b7cf62ffe9beb816c3da0c7c7e9516b02456406290d5b5122fd33a759ee98c7570534c82d23de1a4db375f637c7563544478105fbb3d7413d20bd2d88cb55dc5cce0f560a9163d256c2d4c31ca37d398fa35d089c490db68f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149a8aff8579645424a546c6cf16690efac943380d5556d8c61671518fd4f524eb63dd689a2c7695f28ea82c41b34096f9ad85ed2e529eaebc6801ea0ad2a5b07850039c90a460f6b4570e7e2c32a39aa0c0e3eda164499bdc5dd4825307338706e242a2e157af8ca77d12bbb652ebc58c27a3c80303ae0f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haecff0b88a35d6059462f5e88ebb04abb396e2971d90c9b62a40d6eb92a8f9b7b9d10cc853f056d9d7d553b24b225ea124f3c484a3d90e18ee2d4ac08d4d158907aa4eecfdb3e91b1fa566bbf5aba88980dcfd33b3238cc4c18e7114d026bb96c736cdd50eb9d0e7126eb4efeed0975bf8bbfebdd9906035;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f83a5a8ff4255279ff2bf2fd5c6041d920acdaf2a8050c64563a8c7dc42d8e5682430864d1b4b0fa7d5f54cf8d9710ecd5b55adf41c35d8bde462d1e2af55c486fa89b939f611796d247fd7fadad7f7df959bdc4f4f7927497c98e3059f5db4d11d673a782428361a4b7427877a5fb1eb5ae91f22f8802;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6442f42ad0a6208a7aefc7632c967fb9462b180e189dd4382019ac3074ec334d760bdf1055b3ddf3d4f103d36ee4b1e39b7cb1d013fb04ed46d815ac9e89488ec3f6ee9d9e8b98c74a4388d13c14c12f867c9c766eab001c5633d69a0945c429ff564f8e898023f8257bd77562265cc425057d8e5c8121b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f92780341413f27f65db1cdcdba86d56427e6d61e40d6b37d717451cc9fdddabe9fea44177a54c4c9d22178195796924959c4d2e7dd6f0c03f42d30a7619b2504e8c7a4f3273dbcdaf3780145e9bb172a9bd6fc4523dd991532a0b78a017aa51522dfd18c8a0e0c8397417d4268bcd6c6dbe9d10aee9dfd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a145f75603b910e13dcd2cb92aa20ea2287951c29bf9a5a79b593e7d9877e94a76298bd07fe05d2d4a3af1116643a88fe2872a43bb8736f058266c0296570d0f7cd479e3f215c10a93bdbf3a9992c15773eadf945199cf843d505fca371facc1e0953ddd8a937ca53e7e5b7d9216641a0810745341721b9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19a40f27b3b580cf6fdb537f1c0d4d5c090565188f4dd203dbe8fa45d39730cd3846fb6edb9529d8932c4a83b76e73417838e095f2ad8c23cebac29981ed62cc6178751f3761c826c903d71d608642e7e554edb0334d5c9aa3a48ad57ca17dc45b3be574da646525b805c8bc8be989e57f96a5db535602cfe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h825e5a811ee41f0cabedd0adaebdacf879eb82da256a088630b400ca6bb2487174bba394b9276d291a021293c700c67974a392492572e6282ab5adcc1d70c66b965023aa4b30ab78ae03a2bda287b27b4ec685e8c2d172ac33c0dbf678786b68e306f71cf0687f649ccd0f6000759b5b16a6494057f7d882;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h816551bd68ae7ecf44550d81d917a114358bd63d2c160cf29b44baa390b484345f51855bf37d0d3e144263f0791c2237a054673afd46d9caf64502ca59e64a06d198801e408bd7f73ed0c9cb8eb6d8fe54730704ff8fbce7d9c7aecf204532d7f8356449f685082576e1dd49c7990476e6c9dc748c0aa8b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146fef28dc15f0f9bd7a55239ccc815d8077a59c41a4aa7d7e3b314acddbc69be7751e07e69b297c333064e3a66056750ac2fcee6d7e80c5ed0b7c960e1c65e6e864be33b4857dd0b7ba28737e6bb5c3f993d24a2f4fd04e9fe2a33fc909a0a7197cabc4da132b4d9562ab9f9085401636d7357f2be43114b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b3dca7f1be7b64ac5716e15ff0c5b2e72922b7b8b949b791333fd7fa7bb773a3428e0ec25d0263150b757ab08e7fb848053371ec361dd540af3444600a96b713ec974d007446573161bd31ffdd637f3e67f74bb7bece9486971b806d5390e3e7317ddc2f0341c3bb183f3d2fa9ce3b244f5f70f0fea0b12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9279c0023cf51e1ce5dbcb0191feca39a8959e01e9e93fe33c52fe218d0167ebdd355124d523ac28f1438cf5586cc84ab4719692c2804aa4eddf084f58ed108c4dcf1a397c7e28b1af77fc928000dbe9b53afbb92a2c2a8f3aef5b7f3445c81208caf45fa101f83784f5fae537be0494faa669e03af9e4a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1303ba0e9e9bae3dc84e07791a32711c99e74127dd8b87ad14701917e9505b56a9ec4a0637771ccc80952b48533305c0cd40f8662c9047fb7d0cbc8843681100d410e6a6ee7a50acd246b0c8711ee2bc5f7d720d6251860bc40e5d32cbf9bedaff3781ad2d33979dc46ddef530e8afc3f69731f5a1e4e74e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ac3d37c4e8b95e135752b0595e0b1f502b3f787747fcb87b1fa8a7b4e491f0f1ebc39bfefd3caafa99642bd28c88871853cb19caee22791d2f9a344f0b00680aaa0df8636e59b1f04c8612a71926c5ff3175c11d9c9215ea28a4e3620ce25085fb8dc05a1d167a00136bc097297b2c26288cba85d456fac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d621c8f2fea13975b067f0e8ec875623a07f60dac7a17c788b7f1f514d3721f1ce9e31822b0aae79876c645726bba5ce78f7522f63ed23be69c19a7a81d9bef1361e8f24af1e5075a1c51b60bb739d54af078f15245cb8999a495afaeb33b3dcd0c02e20b51a86be129c16aec4c7d121cb7e5fd74179b7ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8426600a1c63f3023093aec248af7b3216b0047434d1b9c2a59bb367cb84624cd8cf5de56ff277c2bb2acba6883dc879d33bf310bc3612961fd1acbd797273897f310a6ed407056a0773729f8027252e2da22518b701036a4848e8e3bffb0b2b26b196879b6797eda58a4ea3ecdf6d2a1cbd681c41a4f2c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d3c723ce26aedc62ae7393534e291127d071d1b47240262cae61fac6f3c6943598139b837eefc22b304007c5cc1eb371e7327abeecb63730a8f5eb095bdd74ab63af1c2a2c5f623e58afe4732dcf91fe503e4aaa4b9e5728969ced5b2d8f1cdacbeff6ee91c9564cb84a2c3b26f21226bed1f25ca32a3e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb4f0485e0ab8efaefc694772471c6123149045c7ffb4671e24b971c4785ec158b7f40000bfdbfbf11386b0ca349eb265552938639798e05c7420266ec29a3a57c3030e6b4340eac2a21758202ee1fa9d0a3e5d63f077e215ec37bb856281655d3a9bb584e418dd92872a559312426fce8668ed98a63b8cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b8a36596ecc425067a0d0323ad026930c69a349c69834dbe29240ca01294e1c4d1c0f0b8d7a49058e5b487a38c289a29e6a987ebdaa308076ef930681f8eaa663988d8a95931114961a86ac2903f81d836d59fa8e1d4d6f843b158171b90a0fa8b32b9b725e13e49cf8696373bdb971ed4503d0d0691e37;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h67e93b462c130340a185c500e72b7ca3136ce795f529b036d1b378f63d7fc962adf42b1cfea3a1fcea6c2f1bbd499e923a0d24cbad9ad04a16b21cd07f3b084adc86d8c548ec86cd420d4c49cff8a292901d96c588c5f189c24182b4039ee14017853b50778f109a9455a464e1581cb4da4afc641295bb3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h185f90dd1c00af502142e1867587ae189d05d66824dd8820aa057eaba826d3a2a8e7f8d6ee59fe9495b5d3dc2993c2624eae463838471dcc82dee46f7e57c0a51527cf4fb3ae144269ea37893ae2dc20d12fcceb29c16ed4f90379fcfb6e00b9645c151a5df58a4e0b0d1a5ec65e89e24a4a682486987f828;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fdf235720f859341c3cc8734058918dbbb55ed745d8bfbe909937ae78059ddf4a59183fa839789f2d7ea16d2b9fdcba392f32de2aedc3dfeb1279accded2e99cbe44e4d9f739f4a18daf09148a7ab398e93eeaa48a637512b99c5e205b209e02299d53d463edf3824c4432e993be36c4885e38627de92410;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfb214640bb032f2c70012c9269294137223eea339a12e5c619ce41e3a2e15b4b5fe275881dfb5da9b31e253aae37aeede3455617e8f6765d0a14e97512904810bfa5dcc54fe3921128739d20835414b2c32cc1f0b30454643155d4ce6f2185fdd713c999c1cc4836fc004741865c1508f1cc418d0f865b88;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b34dd880487c4fa9ab3dc8024b185cc9f4ce2fd8f22f2aa91ef204c88de6a537466ff021ed974cd7af2791f47050ebc068e7a498825efef65bb9cad01f9b95358155122bc2357e94b45b2ce62a75e25e46bcaa9c267cae80e5944119687a230d7624b8020ec392f1dc8705f5cbaa4f08905ed59768e0dae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd7d6dbb805847c042ae179eae00eb79f28bb047acb983a7630b8bb2ff88a3af8552dd072cc5195509cae00ce650bc84f6bdcf9308e643db8a8196cf97e838a8e18512f5e57d08b61ab7a337abbd119354d58f1e6827dc32057c7abe6331c244f2301c8a054e4913f4593607f336e70dea48f3e7aa9fb7a5d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d68bbea83ff5f285a1ca62e84d3038c0d8f9e9ccf44bc5986a6ab3aa50dcca5aa6a3489a2adc48cca6dbcb0414c7daca03c578fa0cfcf9ff42dbca12e67d45124b7ce11f4bf6a81d3aa485a876275069bfa8b2c4e6f422f6bf37e145dd30ca39bc76eb7791444bfa5808ff50a240c8158f41617930baf1a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc015c236a8f4957f733d879f7a788966d1a3d59fbafb76f4c1567ab3277521405e8a765ce333b0ab269b000ea335af54e4c9338ad24bf84cbb955cc2aebdd4667b79c059988ac4999539ad5e37ee13d8fa26d0114e41e43127ff374294ab5529d7b8a40ffbb52b3ed6a3e65e15d32df4efa5dd12e6b8701a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18c39bd80a194d728ebacc2b8efdc8f8a5572f8a8d9cfa367aebcfe2d635b42ea0bb3cb504358cef7d38a994eba674359f9b083439be0055cdba9144c2c8f2b5e1a51ef128c4d6d175d4e02ee3b0e4abe538909915a6f49a2ebf147c5035467324dd247331e4a40623b1ff350469e03821cf749c4b97ab874;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe3b6bf1cec8f0d1e3045f18b58bcac4139616906a7ebde07f785cb23af8e1a1c3908c8a1e1cb1ebcb394df9bac6b7437004b1dc3b7dcc4b3f0baa25b6cc9490605c285ef5401fdd81028844cd2eda01747fe7dee7d614686e61f30911a347c4bd9c25da1eb1adac76abd2c6e341da44aa3b9af092437323;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4909579fb6f9912c31f6a9f0845a911bbfff4fa9907e46fc0b03c69ccda827c6803318693d86fd57d8c1e4cb52111fd9a1e14e62e0c1f45676335b93e9d1b809d6a99c6a0ed0c5387b60215e2bfe7f0a7a0b79e4ec0fe77e594aff0a320a0d24f8d3322c5683e53516d9d80b48264dd40dd4fab4a2e7cba5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2c52d35cb54d21e8db764cf1c5ef7e3a57002977235f0e04e275c68e8c138f1129a9f7be9d437355ae523d03b3401583ef7cbdff62e5270fdc1ebbb90dd6e3b9ed02665c293268fc0c4f0cdff2f352f04813bae1614a91afa2d49e22eab5d7906b59c373e156a4dbd4882602529a58813360a5e9dfc39fc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d240288629bfe3c1e49a95e55e50f8ffe2a246fa9c8a61ef3fe141c3a7ed71e004dcc0789b9dfadbaa8a824575216565d0eab60a590a5986afef19d9895b275ee9670d8d6370a4a53287804ba375fcdee0d1c1baaf4e764e757b7f03ad71968e32636fcea4b00e478727b0ebc1d8a21c06baae2695867ffc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88dabe58d932e8dbd273fdc9420d833db70f00261ecafefd3fa61ed6b467b06a51a191de48c154eb0d2181be61cf283d9350442478293c1e26909a3633cab7f19e9f1cd37d8fae7cc800fb7991cefeac0c4486a461eba598dd3808ce9b2aec31e444770f7553512d171647d5a963e6eb456cc46a9f77373;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heb47141e742f53f5c4d1d18c6159217fe3ac3684c2e3625c8734d6b997abe5e8209b0d78cb8103d9c1221f697215ebe0e16826f038f170e2a79eb532a69dc2dbcb8c8b01b71e0cfe593b6d580e640cad67f5df1ccbf735347efd6fda638837b245d5f84c9e177654a573633e07d4a536d6c48a203d6ece5a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h188661962212bf51b930176ede75b910da677ddce61b0efc487ab34fa35418947432fe1316d71fb3dc0b5fbd8df21b029a43475cfec9d948385ffe8279636327ea47511af6f7bc38ee4f40ea25a6a5b71f996d30c0cdc60fb6f628a3579a11068b726be3c0f2fad437e8ec28fdfd29d6b6671ae2e09b587bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1696f18413a4206ff8be7aaf9994bafb98753c545f884a526e607dc6bc47c1dab05d8950d9cb8a77c193b7e8877660821fdaa830c81cfee0ceddec7dba3862e307dfcb40cc863d1fd6eac76daf8348a2a6fb609f1c5bfe933cd6975be60ae7de6fab02c81b03e1fc98580d42cb70d152545e6c006a6e493d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h54c6a28063bae631ffc0e81141f55373fb1197b7718c13f81f56a09e656defd4b019d314d4685ebf2dfa2500c0d6ab4c8582c097ff6a87673750a81ac877ff5038332c86a148717e7d4557e45b1756742ce78535206ae2ae99904eb87ebacfb92489b244eb38f5d5e92011588979e03adc760686dddea590;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h909dd82ed32d1e11b19bcc016c427d0ed9626e0ea401a6c55e17d2c4088436a5c36280cbd4a704d732ebe775f2c81ae4e3b9d3eed146d4d274bff347fa0285494d3c3cfb6d47e28287d6f09e17e5123139ab362c3a9330db70918cf3bfd28e7e58954e059022c5dad6982e98b5c390f238f99bada94bf967;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h159795476e4b1582c3dc1275b346db6a455c80d171f0505a90e4ce8d3a348c170ed3ecc6380fafecd4015b7a3490c1ef41125430c4ed6b1a89ddb6d4ba1e07c91ffbd97dbb301ec7b730fd230ed4d3b6bbfce288a4bc67faf4e16f20ef0857ae5a8fd58f3f01ac13038878ef810e1acdbb0b8a8a9a137d696;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1dd1e4f72d6fb5b8e43080e67dc0c760cc18afcfbc86d977f0007ef3c20b079cb355cd17ff7ea2c74761a6e659c46ef4f0393d1abf86a20596362d9cc599cb3fbcb501244ae4a2b089814c7c22e53f64491e941fa1adcfe57ec85efb8fe196ac8272462b6b86a89e7f75b99388e16e64d0c270cc141599c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f8ff719e2c3be2e85e7ec8647fe792689c37668684bd0528b60ede35f90078e38d447213dc966128104ced92127a8682b142845967480f7035c0cb5cd68022844c4b2e664b714e88e200686a231020eb7f43ed378bf0b22832f04b200b85a3873b668ddc6e2a194b047d14d2e4b89b4f609c84e6f35d57f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fbfe5337fd65667bb1ca6f439e0869c5f0c1997e8b5a323375df343aa6b08d5262d50bb87590e169db09e6154e95788c16375d5af56ecf0b2f328ec4c7db3579fab1b4188da36129e6a25db54befd499dff3456a2917ee0569028d31051fe6ae984ba9efc88b1b42e958be1058aa8fe413dd36529df95e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d472be1112066341f7b99486eb6116e08e8c4655914e648a9045cb7e349b7503f7a7882a895fca478ddf6e584ebd370dd959475812a0a073a53b3be5983d6a971168a0650e2dd062f36a4834216e14f84704e870da4015d0a8417efc315528f87da3b8f9f5b7dd57da23baf0120cf6c0f1de0074fb04953;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h57379f26d9f19912a554660cfbd5080e614281b2e74927b6b24a3e9e550e57f495a2dccded80476e01aa5bceb64e008101a3da2c9eef12571abfb0740bcbfe0d9c3424c17fa8b4c8f8170069a509b618d3dc90abc2f399b48f9aea7aa4cb8fa564615a75295370e703166314ce8cbcfbe8a9c009701cf433;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2d773758b7a6c664375503748c848641c6af36f67e625dc0e75fef9b169f608465e218662f979dd1c6979182ddabcd40e09177ff6acb5e4daf1a7ae8eb9ec85bf29e70ce883a82f1cdd976901887c7315386ae1e7b7ad966f6edcbbf3b1d8c21eadb71a30c27b87abdcc5f828e5091170e92379d75412b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc06ee1cf3f203bb505fdb73c22fbcf86f47ff78ee8ad7228b47a8bb8428efd94919a2d8a4f53720c1f6d7f06c90769826805d1414682f3a4b7685a24fe0b8bfeab72b0402e4663c6a0327dbc7ded5457b3cb3da41089bd774e0914c71edfdf5b245ab085fb5bef84d9858c4e85bff55ba00a763bda4e652;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1522f61c347124cf951d8c2c5d4d8109f7e11d31044c83f4d941c34797914e7a0b10b04a5db9f1e83f6e9ff00e4346b2c46fd2648794492c6f159c5f4ec5ed38450e6348392bf197d7624f4d6793ed9fa2b340bbda705b86e490d136804bfb7c3b30b4fbfdd71c390c3894314be5262cff4129e877dd8bb2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16cb44186b4e491b27e188256c42416982b33e62c005663431dc5d77abae8bdc633f87c72d2a714cd4dc80fdd1f580fbbb9c23d7ce43b9a2a9aca70dfe2df39a1617ab9b453b9ce18b6d06285f1831c2e3c9082b39bc14c8f51c8f8eb255ff56a14a39f4e52da6497d7f7d02182a99ddb99dfef13d9b8f5a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102e9dd2658154c36eeaa0efe3a7107b4ea23a86c0466af90e211d25594d8e6b74a745966640ac5f3374a3357b7550c867d834881b86328de716d63b435cefe6a11958cba82f8299cbe30415fc55f6a86c48772a4eb829046a575fee34ba000ea9e6352083141f35a22f763c72a9ba9d99c5625ebc2c2cf42;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46c9a9d0932830739437bca2f2db4ef3bb537604368e8d953e0d3c79d00e3b06aba1c766d570cacfdc303698138197953e861ed0fc6ae357e21cd3c346587b5066dc81826d05ccf3b33f7413d4190099053b5f911f807a090162b304eaef317ba512488f0c4f9e0c29147e92530ded6218314b5fb6e7e503;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d6690fc6d9f74dffc4e62facb174f7dc7fda00a1d0542cee0a243038b6305553852857397b44450a3f66e36f2034169a3dc29ff2cb39cafbf05a63041b2a86114062da5a1648866ea22dcccfff5eef00a976ab2fe2d6a016aa756b4c550e9081c2b9e9a6cc25ccd1435d765b4506ccce699521b44057810;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h124b39f67e8abcded89b7e5c8caa4aab3ec92007a748e732e89b91494a440c01837613fb801890be95ab5124746b978f47e6468e00dc68d17baa1a8fb024df2f3b83fb21d7c57b36ed808accf27ea40a31af96470ec1088ac8b363b9ed7dba28cdb3e05ee090ce2fbd21384b5eefb22629aeed9c15932255b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1859a92bc485c1c18319f743443e1f786409decec609374b2ebe8be096d755a4f0ecdd206b3180d61f365b269aa026b6c281556544c3bcba79c9c0b363efae4bf8ca0bb52be077f500b3b241fe55502669164a452ae4ece4eb833587e8e546b18888161abebb5cb2804af0a14b9880a40daa625e133b26738;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h136f3fd47fa074680cc89a11e39327f73275d8cc9fc28817d2f6dabd98d45f39b721b0873fac07975d2f0428f4bedd58fd479464f180e094c93ace1908d95723b819e70651ef9e0f2561b4bfe63ebb0c00268d04bcab721fa6cb2fe57bec365e3081209fbb6a77fd31f1597e9e6bcccbb1e39811546096ba9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84a8c629de4fadecc0f20bbbad4cd7ad948474af0df414414ad22b267e8ee481c055d3c9e63c99735c431329b0588cb4a3aef3abeeb729909aea64a2ad9f0db39f0946b9da1d9bd6dfef399acea57184b2e230a388825db09d67106912765ad7422396eb9dece227c63581d4fa1149ecfdf9101d05c17cae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fabe6f27a52ff581671d7eaad4418a6334f812970e9bdd74a1ed5431b178b181c6efc213f83506239a4968fa16947e53f55840b766e3c37bf230742e0afd77ac9ed0bb5df26f75f4408470c928cfd01de2d021365dae2243e5da1ef7c5161bd813f674075a38df395660443193f7fe39b48c225b206e10d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c846368b9a640d8d0d23e2512720180ad41a1a13bb4cd6a7552fa2998f29122515c6958cea7da898252bd8ff108efe0102f8353cba7baf0ee5d9f577a620530bc847ac768210de0f5b2fbe754e525d7fa8ba78ae102fccea9466c5cce11b970d4693f61b44fdf355f3a719e72d3b3c8311eede65aedface;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151d7463e6f6c2a47b1298b9b3c94c071b545cb675f4e5b5e6c406584febd4d3660e02b0ea291ebe1d95c1c5a4933c095c753ad4ad0b5948a40ee22130fccd6af0147e42f5f477461f416af59d70c1cc7b2d3a9795058f2c71e5d9108ea94acb4c91737ec654dc5ff5cdc38206279203dd44aec4fe705503;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9a5a32ba105e7f760698137b87e1e66a6a8071ee9b9901c44a34850e62631a0296ae714dce4d2b91578c66aecc89310e5cd99ffe0c8247284428f2336f8bcc88d31e3dfa76759e84e3de72b7aabc408036e97fc756ba3f5c6f28ad05ef1765f2d3c76036b117df36948d083c82bdffbe6134f11207e508e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h67a5dfe3ac0c1dd469fa2a04730ef63478a43049b36ece8f093ea5af90d5ddd99dee2620a68f523cead1a919a404edc26f02edeb5cd889b87ca73dc3c80062d947019f66e50a8c6065e9a5ffefe5faddcac6b3a677d99ad0d100d039d505216dd04fa93423da8b11b9de24df0934eaaa736ab97ffe115d81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h30f39e559efa7ad69664c4c1a71a04fb906f7125c2fb42d0f97998e8a4adde3ee96f6ef7a2fba8a349cdce09b41cf768ea025d96b3e9bf0dc372c3b6bf4e3a5a3741ca75b23dc0c95343e38683d1ccd0dd2a2bf597f928a8ca41d8541f0f712d239a06c9e7bf34d2f96d947bea0a775e5092559054d8d326;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbd3de01789dbf4ffd24c1bb0f10b3047e8bf4af88d3a4764c07991516e1cfaf5aceb08cb3c39b5dbd212635c3add0ff51c81addc03e08daaa4022d061d109c70c55e2df0f23ad3aeadf7b2154df4bdca275120e305b0944abba243d41b5a2aa998771ba19157a7aff61b83e8d5f391a05053121ccfcfbcc9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb47a2377081d5ba2cac6d2dc37e7e1c306bd17c1b92f2aeb8b30bc2628b7d0b3087c8bfef2d3ba6c16ceda17da62931ead81fb60716317b40105a2d26d4211d83832810153297ccac2e57181935c3ebb9f728afe4fe17fcc175a095a7135b118816b2aa1b488b8ce8f00d52b0bc68b8ca40a1be7b9daacec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b6ca8266b84fe9a09cf8630de80377238835f11df874674f875fbe164ffb4a3d47ff5feff4285e88d65fb50ccb25274bb5aa10042e77f94c3b6c30e4a0c38fba60ea6d50f9c1be9bfda58b9d49aed5df0222922e4fe4488c7fd6c8dfada45de7c02310ea97e0e2afc63379c0f393f308f62ab4481b53ce6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b64cbb72861975492e91d91f5e81d285b28f294cf372c171ecaa322cd87721dbd8bcedbde0e71dd68084222f3ce5990c64f2f8c190d3308914fbb0798adcfe879dffd06e6cb62ea3dbc52af446f9cf00939535dccdfbc1ee4b199142b93580ec809c0ebe396e62b3ede2fc13f15f621a14a2918c073a6cf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h158c23aca067e3fa4f52564e643823e3bf684cc7c3739c685ce438908b8f7d16b802b91c98a3d411cffbf7ddb7378ea3e8bac3248f8cc3bbf744ccf708c3cabc19cadaa69b354d107a1b18b7505e4d39ae4e3d4d5e622f22d790f3498b2dbb648dce43217e760c7fa11e77cf2177d4c866cbf3c55a4a42f6e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h798df56442a6a31b5144ab45e3bd74bb7b769c7aa04f935573ab905d305707c1c1a6bc25ef3d6b207ec4979f481525ef8e769bf79d70b63c386d2868b97b311c391eefdbde999ceebc1d2711bffc40de8924b3d3657f2c89ac0ef2f94216b282d5f3918fa25e0ed237a3d48f693499ae8bd9f42f50b6ae48;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h38bf75d9bcc1786db67a11e72ad283dad2fcc5605540556681bd8f508fcc886b3c087093f421f8a90906af7b72abd9c51ddb289ec1ce6e6c903df2d44076045ce7133a8d5b0fdd097c345ec3dd409e6e3fda26817e8f7d7ee35444aa71cfdb367a21780cb3aa0214e8e920a9f56be2c650eee0c53bfdcd47;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hefc2e010c2225963914c8b2380bf1375850ec98b87ce37cbce67cc809f935e74d5a54518460bbadfe164fbb4c42e3128f97dd40cfd30fc50495772efa59acc012e49be046d8816194e65e0f98670a99e3c6bf6eac14f06547c34352e3283a255bab2b442ef0eda6f6a30105ae21a96866de6e764ca8cb07f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf69843e50bf1d489f8299285ae13cb95a8df38ae006a854a088b85c42135a2b3f579531f446c210d8a2aebe41525d2c357404e3057df5c67e6778ee6b1428bc377a0e6844a6cadaea301c50aa338f467e49d2b0f326a20f86afe7252765c1f514e82781e833a0ff627b79d42db59c952605f66ffd3bc729c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13179135cf85eab1fec7f510dd22431ab03d164fa4cc0a6f21a44822124b39deec656e53aaa437b71a4cbe5455f2661cd2b474397381cba9dc0d76e0baf03c59b2ab5857f30c6498ed7ae636852040a0c02cfb32bb518ef643514585ea04401154b91d892fccd5416b17ca8aec219ed954e0d496fd9ef3f5e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19ba8c723e120f570faa56e6109402c180e2d8e03ab88fcefa29381f0256b97d1620af3403703f4edb65822050b73ab7b35820c2ccee8a219e87cc24c4630f15d46d780f87ebc21935f9f7cf9689418e877c77d23fab05b006ec4f1c998b69d5d2074fd9add87c126f6aa0cf79fc64a34d84d6c5195594c2d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1526fc46cee7eda9c2da16a0b62e9e2dc9f5968852fdaf3d8d108fe2e678405a2161e57726b52b360a391e8441834e21ab3f2622980af52ee2e53b2e35e951766082434fbe3e56a76b29a74e475be376410124351d7b237ef529300a6ec687493f703e8583d828948804b27177887f6c0e8d8240c636ff43b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16a731188d2ad779e8f8c0edd53336445d504f003e556b1c0c02a242830b5a0de47dc9039aa2c3f0053dd16e79ab8ea2675d5911bf9fb3e409eb70233b82dd68ce2f58d580c167323579b2545c042d81f210568eb995aa160100136a03266e9929a7b6b3f027706554c609bc1b1eccb8cdf488fe189e6eb27;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9f3d04f5b29aefcb3fcd039ced73de88d0bbd964b00df6823d0c8a5c1b3175d8e522c26a671cc73c7a85aa7babb6a3336533b995dc16b629c660a50e7ab85ca400171a0c61f1e5716cd2cea9af1bdfe05f445d47d2cc3877b7ca4ad2962104105cfa7ae3c68df1321efe675461796d58f1b3e7f13051a4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17affa74d18c0660195c58bd317cdc176071ccfc10bf92a8d8ea059f52f9d7ac70ea9b1fd19fb2319eda221bd5d83d51e3f1515a5e01b0a8f1a8cf870dd152d719b96b69d82d871c2baa76a42f099ef9d83a3e52cb8b42ed0df20a417c898ba1c32c1a70a5fd71f113de2d395460cdf462247056dfd334f3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdaf6dbda811ecc774a43cbc67c6ca665c8ea65ed518c6ce8b6778d969eb5c5d91d06c53e67469e973ec923cf98df57a0777d7ad6ab0fd085cc4c058e26e177e0103dac096f63ead542d2506bf183c236fc1be451ad8793771488dd93fbd44bf9fd41a512710b35ab541a285031bd2ee26d63dbeff58f37f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6dd722ba514fe849ba46b94e3a69858d5ae0b5e56e2aa175cc03c3e9cf081f372fe695ceacfd8d53725f033b9064f99000adc1908f52ec662424b42768c75b878cbf2326ce08ec81e60e1862a333d59259e868cade0c08d362302d9d091d443296756062da793665f59a79a39843a20c03d1bc5bc5d8464;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e4e73a28f6eca976b7db6279fff850fa5b72dbbdfb04946fe51944610b679a8145d67fdaec5f53a180d3551f5c9d376c98f3d6dcc7122530b9ed844977b59d40e17103d885a2478b57bfa36d2922ee2008e68022ddc9bfdabffa40282eb3a95808d9b3db464b0cfce3df0a69ae90767e9370f826ab6ac153;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e7c4a33d0695847c53d7dfec2d07ef51b8c1c1a79ad75f458c414e49e65884c83c6dd64d80491cda55bd2bf5542b5aa65b9e35af4a3f55ecae05e5355df18505718a2d41965459d0176baaafe6c641fa56803caa8fbe093e709ce1a7ef781f7ede8f04f97bc70771496af6270c214751ab3a5bec80965b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d260a5fe95a9ccd53812ce7f89e0087c41b28ecd639edfdb3baa265ef8bafe9df2b7e1622bd606132807a528376613b854a4e7ec3949c656826865496196fd273fdaf187efbd56fdfc0b617a2bb79c1e118da8a9601457c74b68be840a7b63e37c2d5decd26fe37e30a47fd60dc8d86ac55124b43e495c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b0c83da6c4d2c5e14bca0255f9eb46fbde8c5eff30b10bc1aedeb1460e447800d7f07286190b0a80268364194f8b58013ac0d12914d8a260fdc50c213783a18d36abc1a7db1c95426378f37cb58168bf84a5526c1ed2460a16acf1bc896679824ef44878da8c46a784eb31468c3bb49ecf3d44b0616a63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h197e50c3319d3fe648e18c3df5d2f89d1998fa62ecc7a7711851747384ebea04d61a48692aa570e877277de6e3117f24f9aa201e564f0baa4dc08b01ad61c8fba486f50e0e8d00b0ea9f2b8d286566ecba308855d60f57e5389eefc21f289faaef5c41789fd8b9521b011ab30c919126a756c3caf0a3160b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82543b04deafa82e573f8a792daf4b98b0f9103682dbb8b4038dfc9f270ea4197a5be47bfd8f8fdbe9f955c7fb4c1a1cb872b3a0382a7c09ab11c6f17b087cba122eeed06ab842bcfd03b88fbf9bedec1a0de1dd26e330c36790badee7c64ebf29fd32ea35448a2a5c56501a0956b2f95a783a6f4d45f154;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2217b56c53aba659c249201273c7257196de589e78d8635ab974eface841bdbeb83d0093efba3d1be6a0d0b325fb1e4bc3c11da91709fb71b52afc1c2da4b2e5681e2b50e9faa134b51fcab5be8da00cc2fcc7a2dbc49fcb03bc181a53df38afcd038ed203912798d93e02ebdcdceb399ceeb8061cdbd39;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b1261c2d881ccd651974037728ad4551f2c5609a768c9b9b15425996d348a907e776ccb619863e92220ec4f715c855189c649b990ce62a875c4caf196ca7f292bdbbfe89dfc07e3649b23d7bf40a06ac77a06ecfaf10116942cfa0e71514139b91882d50d03ba3969282cf6ac61cc748880051688568a632;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1391b5abb448c1d986b2dc314d2686d0e689f88b72325c429d7dd94ba83e5fe2af3e9fa3d33d4bbf54d446ba16a06590f0d2355bcfc8947be4b5db1535360e1b70181c1c02a78adae25d4acb76d3a961b3d0fb70c5bd808ed7756f36164eb01e3d8e9d546299941660936223aef6ae16e7068376027a926a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h166a8772cdf53b87927597da67fe19d3ef1763c5297f9ce30e6fb148f5d543170300ea38eea252b4765eec7cff077ce2134fe0529db24414df5e59c2a714f7bce0ff77b100cbc2be8fecb1f81f8886976921089037ae12ec3eda4114d67ac2dc3be05d3efe93d3d1b530dbfb7fac95c2e266d0fe6bce8ba93;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf4f333617bbf8af0b75ab4105536fd90b17116fc11d3d6451f3721853fffe38de6cf7a59e57e27a2aa9975739812321c626492d714f40cea641bc0d69247f3b223007a8163010a0ecce6ac476f7fc6125cd862d77b1ab9a231805bcea4362ba99d406672893e2fae251d918eaf7a59c26f4a9f61ab4c7056;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6729659aa9eb54b06484fbdbd8d93e7e69d43801a52cd80e782adbfc028748953af3ffc32054ddaa327cd80b23f842abf5880d8d470918a0d485efb9346e114a53a191efa65c2ec1a87e311017ea744dcc1c50e2640775ed19623f814a686f6c3d9522bc37109e980f037b229155ab131a57d89631daaf3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he73c63d96a9c9db6ecf36f6830e6b7ace71641a161d63e45f9f7eba6966f06b1da7a4664d3b1cbe8ec672e0ce33c0c117db7e8585fb6c21f066dee670c92873647b802f329e4eaccc27d31b1087c5b8b41206bd25ca398bdac92f1e25cb5dcdd90b97c1de5cad715205a594b24a1e2b899ac41689655e430;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h161351159eb0d0784b6d02ed45a1682fcbd2483494d61c1e75b4bc7c9b32fac80925dbdebc178f8ebf49535db4c17c65688c62003db890869d7aa5e81a2ad5d95a683126599899050865df7e3c8f7788d6fa2352173f4eaeb020fa3d585dc2b41d83478448c0fa47ddcb1cc125fe404ee9e95d9b6e6b616df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da6089c8e697b8669fb0950c3aaa46f4ba606a16edcfd34a99fdd8c4b4104d47f2193a16b29ef6b5edb3fce21fa3565d34bc45270243e1420bb7a34188d58368b5b4eb2501a5c7072500469ffd2b32f6c7134838bdaa56aac86799fa2301f58f729436cdb7945679a95aba215c6aadc290af599eaa30135d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef5753f8a786fdb0e507c52f696f254e76dce542dfd8cf914f6db7c92896f6efa926e7a857db92d6b65682f8aca09c9eb3fa381b529128bf6508c95bb4582c6d033e99a868263360816fcb6ceb76848ca81cd2cb2e2a9cdd99618d3a79b0c5ed590c8fc89b631640ba502ce7241eaba2b2a442b67f61119e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h290f02ef401cd45af65b9fae3d41ab896a17a39d27869b8770171c5f7156dfd1312bbbc23f2a131abec0f9bf2c55ad8bf483f9ead862e71f26a03fa2c28fde521860ce8c2eac0b61e35d7ef34bd9f8a97e57c3a5f61c0cdbdcb18f1105bf67ed181349b3e4a471d164d4e13d2d72150de783385cdbb09c58;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h27263ff75e1ce8aa39037d48be4ec2d03c5be376a0d57f0449c3b6306b91488687a5f841fb5d219d3a05313c07eab997112d9378cf58fd1d06cc88eafd9ed5784d5758c11953fe39986f73b3df38fb8aa0ae5d66e118e32faa530a240af3a79b79dbf574029a8667523d619dab8749776abbf19f3e0acf04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd784a5bece46c7ea093ce1edb22bedcc66ebdbe5747f7bbd3010f460f481b6527416c000957b4e67ee5faf1796067cdc0c5908555d180569d05c3f97ea095d9c8744273560be09baa8da0d0fc48450f9fb2cfa018509b94fdcb6d7eeeee22c41b2c3e0b7abf1581933416ae686593d730157da031b5a76db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a32c45b865c438565362528e177a82aa8c2f51546524ebcb077b3f668ee1ca27273430c44ef6d30c3042222b09298129f4a6b796d08a5149ce3bf256dd1164e92d33fae1673dce8cdc05ffbbd183bb1ac5a6c53c97c43878a2fac46a9fcccd83eb68f757350e0d2ec55244318ef28836eb4adf0a35afa7c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h886112640c4b32f6f285d16274a165a9ea3e25bedfa41a639e2765d710de655d6fec5b43a97a3e11a6f1d7e44ae9a96a60dcce4749e9dddac4d7c12ab7627295ee8f649f54fcf855d95321cf4421344d1a59a9f4226082358c2fe8b8cda3aa6a72b07dea767c795028b3f1b16a761b290a9ce23e00c7b74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193cf93c1a574b95f189bfedf9ba871cccea5cf6c7db11997f88a5c18e20b99721a267504d8775e560103a7e485124c1cfd4bc574e4b3f3786faa0f703e271dfd59975e174be3dc048c1505fc562f10f99183f9c00845ecf07bfa3367dd4d4d6740ae8d1b2bee87977fbb3511b6f77e5a161cfa343c4cf820;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha1b188765edbdebf774349868a7c14ac5e6c7db2f9ad5f0666d3d6da422d17c35c3301d5a4bb101ed16bda10dc12033e42e695e6d8996134ffd5a3520fe2ad9e0da074b83f03068c3f27077eda9e11758a95afef24e62ca515f68d7c1078467ca02f8f6669de96b6af56e5314cbce03ef944302135ac7e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71e915a4d98d02ea2a97e83748cbfd199616373bd6faa7ca9f4aef06e6da413c4fd2dbad42df622d9415a2c80f22fd781e87e515757298d76fb43916b69ae67d4de9a3d5f69cf6158aaf82d10e5b07d983ff573af5fd5c8abb1346b4bb591081d5fba0cfc429f9e8a5554520a210f28aefb25841f9e9742;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1751194a46afdd30839e4f3030f3ad72729afae1845d47e900511ba9062ac95412bb7fd304bbc6d5f86ea3a63ff788ea534c6f4c1a811d2ace08bd0620fee551b9327c3cb96afdf9641b3f4a337353ed616215f369f6b27ee176e7ecee37bcfdbd8840c4594c0394bf8c88d1c46317557825430bac9d7a182;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf70eef32369aee660c16bf78a0194c9edd1c4ffdbd96529f0c0f01d0b9a8a9a76237237329595f1c2741e5baa2e80a9305cebe14cf495f577cc2546b868447ba0106dad07988cabea1317e00fa06ba38da35586777dbc73ae5eea91e2256b46811f110adb43df1eaa550356250528db3a8500867834092b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17955832c4abed6dd04c1ca2b5cb9e2dcd7ef273ae54ee8b0a94107dad2975a80ede458a8a655c24d8d7c2241aeabc589768809ae39a1e26e0f9574d86ad68dc2b4182230cf31279c52fae3d3e300d93fb5a5e4b6810843d7d7a40f08c31827173be7647a1e8da0ae88f0f6b24873a0b0504be2b566b0bfb8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd66782eaa101a7220941cc7354db54c3cfb329c9a959164d5bbf3feb5a00c00060e11d8d9a3e0b2177d0e483a6b9b5bb78817927989c6ca596764dc84c3b818f9de1cdf2aa41df094565fa910475aaaab95a10c0b6815b46ff1915fed3a0cf2a1ef0375d8bea2aa53c403e387183c9fc8ec4041b75a3059;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f23a33cecd799ca8eed8d1b0c009f7220dc1a25e08ca88f786128da5feec817141bb40177bd4d6984aba5e7239decd61db65d5482e161cbed9750d1a49626e0e3472d57c5491e0f9b02121eff889b9844c2c355a54d7cba134a1f88022fafff805aa17028d68f5a7cf85a5f90b2a87b8a1c1b8f1afc45f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b24b09b1683fd73cbceaadf8a34c02dadec765cae0fb93b23fab9f4b7acae58dcf49f61d27089fc9a1278e64a7514ddbb17f59d8b84efd4eac5eab2f91cb627b2406f6569349dd1f5c3bc44c44bafe17d68e79f50d7307e0f983b6975484dd65f81242183304c94f9a23f0fecd5e8ceca0e11032f4ed4756;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2eca7b28491d515d6ef1428a4e069a1c6980be522b8083b9f9dad3b6b4e84a59385e4f50472638cfeead194d17648b56993539ca6b74e77e808834cefaba26414b549f10a8cc9116124ff93cca2593a52b0d2a979b0e34cca6a0669de2e6a1f76571a63836556943b41e3785169fde5597ac2f6c3bf865d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84f0921b919b7bf21cce961097ed6b1cbdd4377da69e3f8d5d7769680613bde3facd1b3a2866863e55b814abcc4977e229df8283f8b71e941e05cc126b08d884b20025f9f3ba95092e3376708b7e649ab82755928c7bcc6b89776b2a5ae90ae2aa7460bee57a699d78acc2823487612465c95e85b0976a4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b8f821933e73a473ae2898ed81007b7331859c4ee9f2e9d2c2f146fd2a46e8bbdfa12562f6c7621385f106a641402c10854ef34bf7fa5b4c98597a50b8e0a423ba74a28077be438eb1a9f5ac7f214948f80b16c576d93e8b78dc6c48cc75350996bf3e3af98b11d274894f9466701fc420a2644e5ffa3601;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f02dd7fb9cc53f72c6627b6f7e842d34c7ad0f1e4b27d854766a917c03c4263b01472d0c3147e143c56029653046f16cb7177635162666f562ce2c5d4f424e0b9813312ba8aa7d3dad21fe377a2a92e2a8501875d9d85cf9b8f7e4f9a07e110917b49d8d0b6d8f19a712ed263bba68b339b498d2e1874343;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he48f432a5504695456b763fba7612548f9a070308b0b834e0cc9cbdd3e878b9721ccd7cb7f7ed467a41eac57c55a2a7d9236fe34925e30753214820c2b846cae90264623a1fe0ad1f7a7363e6cde65d4dd2867262a6a6125fcc25830678243968e51a150b1cc7be4cd9f6dedfe6b8e3ff172e7cf3f7fe783;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15ad5a9a4c591584a25adfa7ff0222022c2acf64ac37814289b82f7289fd18dfe9c7177cedd4dd3f8590f74b1a23648136e7573276360d55c4fc7f5fb02d8eb6375e7cfe0f34734c824dbf7f755ca2b9d571d1677b28ffecf4b09c189ef6eec28174f0321207f8e5774b86fad43585eeddcbb6661fed725b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18997732b33ecd97677c704e4db656f21e48336d58afa6800a0626e4b9751159b84d8287ef65d193f6a74fd382f7ebdc613e53e8b4320045c78e98387904a1ac66ada2b1abe84309ada68fe4bc10e81a6bc0fbd7f55732ac7b6b35f816bd254972aeb2e989f7b8e5f79b8fe36d412b6c2f0b264205fa51e64;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f9dffeda08bb837393f145b6ba578013aaa86afd4ffa1a49ca3560351612bda77bf64691d6e28749c9ed211e89ff7b5609c9729acddb38130627e0b3b1e44ac4fe5699418db6683158abf2d2bbc55f51e6e48dfba86baef5658bf8d015b80bbac00348db39afe3b88e1d28bac2028c75b14bac0edfdfd31;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1922674129250fd197d58742e47fdbae15a8a7062c8f6e94d798b612255a903f48a21849ea29d94daa976ae6b18a6aea1c4739c3b5ac408df5fafbcc4fd63fb95506dc6d3e4411f3a439a837fc45c67b5a7633be4b69393c567f4990d809395a7e1dc91abe1222f4250d9af0e33115dc311ead3548b59084c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147dadcba122a8371ad8dcfdf12a83effc33929715110c5f98029222535270bf314d1f77a76901490c49c7a36a58c0a68a0d312f86b0a8700fa180f546f8825d5afed92d6f65a2b6635859e0499460bce6452d9724b2ed78e0e05f8270003867710e8fe11f344e1a55696e30644abade2ca3899fb544bc2e5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h179d05129be37b60951013d6fe4742930130e9bfc55a1669ae6f280ff78945aaa944ed4f8267a4a84d009359f70f237f6e12dfd0c30df55620d42142ee7fcbcd3bc3f2f735d5c063c449d5deadc3063496c0167841c2438d1333f9a21fd458453861756549b8f6538dd9c2ed2fb171da5547e0b22e0edbe68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e97170b097f1c35946fb6639603dea05b34fa58420d789252f0017c5dd70bed122766aa820b4197dcd197ab816ef1e205822f9c3a0d7bbe805abf70769263bac1273272f45b4dabb30125899386c4497f4f31d7d0b56c1d546de42758f36a69699f3a59a4fbaec2b79a490f08792f95f0393abc5d4808c29;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1362dd95e1945a155609b2aa3cff4bb8925c8d3df7b1460532db56134ef5e0ae477b021344817469790368917173f02c3705603890f30aba854b43741fdda722b04cbdb2af4a3810cab8c3a357ffd5eada384e641328ce6d16c94f79d098f92682f66195428e5b00384796c9cc7e43dcd748877d36ad8f387;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a8c123aec1d0f9a354feab7706d5240197263cb43ab8b9dd45070babf8fb72da82dcd1c02a3d3ed3272835d7f24a4f3a8d3e805d3312d2d902181b198cb531ab80f95366b09487d941edc36cbd4ca87ed0b54b9063debd3f51ec49e0ef25ea6c174a17e743ced0a40a1f28688c82de5420af8a52925c52e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106d31647f01dd9cf02c79538ab7b3c4fa6100cb2f07845f559b069570264a532eabc7cc39055fc3b7773c26ea1e6562e8a948e4bf69509a77efd56e47d05d8c81ce447deb7511b2befe19efa3ba9d02283162e807c3b8793895e08a824edf8f90961e74190ffa0b077b8e0d8bf6a3988001e7539d3cc46db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc0a2b2a458b355bc8282adb2e22453411bbbaf7db9ae76ecb2988e26de0e5c8899e11e60784d41d23338e4b4457ad53463278416791d330fa0b2a0e2ba5391a8e9a3ba1adbddc315221d1b898aae5668394c7b053ce505a86ac49ff6491e08d0aeaed156d7485639798917b7679afb33b7f991c20f7641d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h78abedd80e16e635d2e012e6712eeecc212745df5436a8dbb51e565623c0eb34c92c231da0ce5038a9cd950d9fa9fc2a3c1be403242a00fca10bc8d43136100952a373c2c4568179644e447c707a952abd97f5ec6bace2248b5b18e60e12aa1b2c076f95cc190e74d46f2afb5d5f630c0286bd09c33e3feb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68e305f66a5677862616fa0c60f93b361717dbfa13bea74c6876425650c8dc5f05df8c02e881a84819227f048411770fe8a1e59e3acc8acd928bfb5d627de516f5efdc04b26b721ad8f1396bd7cb86ed67e753865d4337220a14ee8470d1bf2d5ea283d6745b30e548510806a48f70be6d7d09a09fdf232c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7139c2f23523e38648b11ba81aa35592aad4ac05aaf6c6092545c3d4e5532d9fb05c1506281d6567ac0d589918588c0821ea23f6718618d98c34b5fee6983144401bdf2d278c0fd9929bf91c0d2a19674167b33b91acb88ae33c2f9062e5ab1fd8d3b0ec1199526ad5f6cfa3900dba55b66899d99316ee54;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b72ae85bd3c496f6304de5ea3d1961a00292586d41901174061548823f714d5896662bbfba7b00ca91f31b22dc2e1450690c33bbb331a028900a2d0e01d1478e1a4d89f28082cbf9936e59f96832fa26e34927d786d5bc055d0493549335bf672cccd1fb867c2ff5ddc10df90cce4fdf620a127c82b3124;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e653268867854b94c6edf9f13318c9b418b4c3b69763fc140d5f3ceb3affab50bea3eca0846951382b47052c3274cb1455fbac76f4d4d2405da820c38d6242eeef622fd3d8d90c2cbf7103024ba6d734db58311c02243669d8bf168747348d347e90d19270c6caf3859d0b2e5323fd34249ba6bcda98a1f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h49fd714de4ed190ac86b17cc34e2f554c4cc7cb77e69fc5a8727cc9ec30e478e2b397972ce86f57fde1b90f47f303051bd775239bec52ceeafce3e40635b59d98142af5fe0fc59c48f3691dd4d0269100dbd7a8e658da2c3857b9a3adec16bfd966588ed37f0ac135ab389db42edd05c10db9b0c63e2a6e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5805eda1cbb8d9a1837559eef7d568a21bcfd03f691e05b253a12122b0940c8316a7d9845b9863b557e0cc1eb2cb24af7e50eeabbdebb07a6549135d06407afe8d767f34d0c0d7ffc264117e942b914bc3a73ebaf56acd2da9c09d3f8cf7b3973402676d64d406b066fc5e4e7863a88ab9f227033ce015ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111ef26aa0c57d33a756ea537a1f320fa0a876d3a50ab763effbd836caf46265cac3c120a8b7711eafa4523fa5afa566ffdeaf2353ae4d1a3547917fd3ddcf1630e4470b3f9f5e2df3d882b50d19fffad2a492742cafc3d2d5e960a109510e359b4de077d28ee2c6564025f0011da0b3aff141a906449f9ed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1149ac1c6529179463d1f4a0c9f56eda2963c9e1a49c1d300e9e7df233dce49c9e7837a8e738a8bdc5be088d7aa316ed318e2bb74cadc34258012b4f7b3824fa1b1ae6fd9f6140f87349749a519fe02906ac9ea0bd78604f510101fe76ccf866400a09aa2abeb5b5d03f41ba00c69536011a8bc10a692dbdf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf969379f07d0199ab0ba9d756a99cd3d4fa9e4c9173805b9758e5fa3a4e771dce2e9d8f147b9ca34b39124e36c716044b17e7cf2b0a890e90a8c1c1bd320b906546ceadfb2f2657337ee1bf232e5ef90fa79dcd932f21077ff85f9a1f8625a03f46a8e076cce64073fa51bc16ab1f71a37c1b3156e4f8c8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h95f4c4ab77e39027755dd048e78471e96dd2f320f0b73e208425e3ad5047624ae15d4e13d9c78179239870fed499101a58118abdaa71c60be694304e81519163bd2fd085ac01d593fc6d9546446452e7cd95f3466fa706499bd8dfda1de0c6623a3ad4f2fd653ed3478faa0c9a0c658e63ac319f80f65bc6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a669d3e49864567741e880d2f7dc782f0acf978ef0f7a9b4427a8f7a6209c57a8c7d474063ada38f7ada9399dc5d2223752191fa363548856502c0f95db7dbb732a845f317b8cae6bff0fc77fa00dc146f4d30fa661dc66d0c402ceb05fef934f04214d3c16359e67001e5d61770215fff195f4071aed74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde93bb5098fc915ca31c69acba7daa9e589845ef9368b31592a3c8f56d4fec80560856ee00df72733de54dab02a091eda513fbc7c3f8cdec715e721e218e768e04100db1adafcb51706357c9c855505ff12227e9d90c500caec827672d77526ba72f30f9705f12cbab95650b525d8236a7860b373236870d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18bb7f51f818ac608ca7bfaf50e6dc65b297bbcb9fce37e795771f35f1202e99f83115499e5a453a68e27b91d770189e40fe2eedf859c4d1f42b26e339f9615fa308726dad342997faf4b1566824aaf4322a32cf05f53d359c0f1b1b43a50e118ecf0aea323c19f5740f94726685762330e11c478ca447a56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef1b23d7e69ec48e0bd5f849c96938298a597948a27f63c595912daf09a9b639998c449696dcbe48fc1e713d59378203ee2f6df45b3fc2a8fdbc7d919ade0ac46efce955e72ef9dae5fc70e6874ec167d4d18760433a4187dac3b1b931f71201c1d270d63581be0fa7128e41a693a545a64862632c40be2e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90eddb9999d320db86d64d72b4e0c22ba923cb7819b035e4e39691b85eab353c946b9c697c62777b039cd0d017cf522e5695556a349511a7106d28f069fed0d00d79a827b22c655446c5639dfb5af2a38bf59ad1266ba27c7c39fe4a47ec540bc8a717e152fffd4b43ee5573aa5098f3695d77faac60fffb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h166a68c17e5cc99c3e543f90be1cd4b3a3196608a4a2df37536809120328bc2231033008fcd930b800ca13664c7bd1e1b3960b838707ae7f186583fa4f72117679e965b1f097e7697baffa2f29c5698d7f534c5278335fb49d5cb9d9a78a67cb37e8825abf7c22721d97b8a9d9c66f033a33fed80ee7bf39b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf45e499c989096cd964a90e4369fb948253409e1ea82322753cefb274ec1251c266ba36b763e7dadc0007a77f8d3cff9dff7fea93f8bb32da632323afe29474c192ce87a59a87ab4072e91b3c86d1c0df6df73d56744c3a1099932dcedbf1f9e637cd5b69fb5572e417f9d7108751daa9bbf75bc70f31514;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f8926d02fbe280960858a9cfbe50976f2b912bca40bcd987d5941142aa77e305a331152b70da3d50dec24f9da6c9dc69b33e1b6e3274032d15abb565dc3d5af069d92397237a18caccc2f311a46e50d367c2831ef60bb36aecbec251be218d4357c684f4b378f8063a4dcd78612588252e60762c3295e4a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c4f5f494a9781f8df523838d9cd0084d2178e42e2c3a29a04528e13a9893cafa6297b3ac1f4086768c04dab632b4caf29f8d017e9779fbef61139d639731033651d3340675c1b11f9b62d878c05193aa2bb1f68e4ce0bac00a23d76dfb81e557777d2dc4893037eefc931d5a0a362b506f17758d4229daa3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1005660a6a1e73f0987ac7b3647f6a4dea1351d7bee288971ba0a4bae68cdd0afb58aaef4b269863bda37c41d26191cd35a02b0b847ae84b04cdfd21fcf19eda936ff7dc5162226a53f86ddad8d5c5db74be18d83f946ffc8a474e028c153eb90c55eaac991e05aef8c379940f7d902a7af350c2fe2eff33b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f005ac6fd9054ffcb464b1d8b7e4b6f91f1a3218bb1141d366cb33a8fffd49909027a457208603779bd4c9da6784409d7e72999d9341ab760ef417c1d904e2804a8ef59e044199e37ea3a5ac4256e25df06b587fcc27bc8f63ac24504caa742c66e921ac1e4dae4384e8b46e6efc76030823a6ff752d235;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b77fc4f4ea1962b1442c43de662588beccc4b7968e5a7319118749cb06b79558dee28ca53077ed5c6a4e32d27ea9728e3498475fb87bbd1d0bfbe2f25ad893efc29030c055248859ad78e13c9b24af96382aff21fa6845403938280ca464337303597364f3719259c31314431fc80ebc9acc4781c118fc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14e0f2992b49954886cbf73d0462f4a5e5c0e0d7591e2c7081294bb8b573f47019a54d9b53e7480bec756464bf6a7c478bacb4a71a25ff7ca713a92c1af8c89b952045cc9488342b52f7866ad49f5996cd68c78aa76f4d0c5ec5e7bfa9e238bcfaa840ea1c962a790ffe8df02b46220e8ce94db74fab234e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ced108c043b6ff46e7cec7fd0bf4f9e66c97e844d3e868144185c5693773e557ee6f032dbf5bc74f410fab0fab24e8c93b108e2f41f6d964d149a5a86db347d45a5956f362a69604c8a49909f207ce3ce8b7e7fe6c389d164dee6fbcf086920e8c7e365c825740719ef5f5bad74400f506e9e7eaffedf663;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fafdc63d123f8128d9c1327afbac5a4f22b4734d0ef23f78d3ceb535aedf0c736b4c721ba56fbe82b9f9037eb8ef37c4266ce12980e873417173ce558ce55b3fe1308768ac5233aa90924b2ceb48d25a46831b006f4852a6bd905c6f957785f031895bad89e1c2d19df09515191f0c7193dc1c7d8870ddd2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0256915ef55bcdc17ac93a78c3ccea5b03ca01943bf8571a7ad56cfa7b7134fb32b4d44d0d1cde94d17bce593245b226eaabcbaa378b0eddf5888ac4a539885fa33067d650a0f7b654ef4d07a789a179c7e48222a4d952b1eefe681d28a917fbf70f3d9584bc0138b01cba69cf700f82b69dda589d26266;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15e49fe6ec4a5ae0d0095f02fc4f84e3b7526322e6e114858905b110791a1220acc23955fddfa55427a11c77c11c30273a4eab569e1c1bc55fb851b26bc0266225ba9e81b4a24a50010e921a26e650a18bd6c1d7567fdd50bf0688290b7fa3a12dbcd23fac1a04b9d0556c0243d555095ef61b6421c18bb6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f6b20aa5f10e4f38ffec1be4913b91af713a06b6cd4c4353b9c0153ad8fd761ac505a2d6918d0e01fec2890b46e6ea85c44e6609b8e7485a2b92a2f81859f4acd6cf52c6860a507a828e933f4838be45e9b074349f952a425a2f5e72d9f4b1dedd829cbf62c41f3c57d9a8a22caaabc534e7e4b019eb4e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd77e87db87a0db6f9d16de6cafe2c4d1106662576f991a057c446ee3ecf30c30f386c30c9123f8db20afeb9d3adb829ff5e9d1761773ba1c741459ff3bf59648ca6a31a4ede6516ed0b38723f1db281b2697d22faacc8942f75df098c90791f78d5f0437482f8e55c9902155b15b4bf7938ce1e3258ac408;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd0f51673766a42a5c332dbfa731ef01dac9c472260964305c04e98f545d47a8a320c962c1f2d507ece794cca304f42e776334f611ef3de17a620c087b2501bf56a5ebc30ee584af7eb3d7bb2155f89db16567dcf87ecb94e0d9e532a0661900949b9413f93975fe0fd5ef4f973841d901d63dbeff3684706;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a897c80270ecfe27a981eda7eeee3f66d12ec8979e9a089483a28442e598bcd1d1ba0f28778e1c09fdd9650e2d1ef733d58921f988a3c4220e1fc34ea8e25daf835e328097e864afcaf4db8d711f3b65f65b80aa7e3019cb258d25b3f18bff4fa90ca2227181e072a236ccf068fabe3be557c88873f5c90f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha708b199ec44282b10144062f3d302ba40ba234e9d80963f06f4e585f938af6f858c297e1a88b29abc45ed6f688de2ce16ebc03ed91f24f1f7ee362629e03644f84950469993920afafd46dc68dafdc01b5bc6d3d41bf26d4fa71b20ff75c9c641d088fefabab1d161f7871ed76831de1cb18b9d8542f8ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4bffe03a478ae9f861cfcda60fc78d4a7cb9815bed5a117560f258c8657d288e417e2229e22e2237ebba684925c799ee01daf0d49753ffbc6b6dcdc422d2006110c0fc41d1ee65a97aaedc609230a53c9799c768255e7f9a3c4d859a3884c0e20b430654716185b8e3aa16b9ae749b072b08f532a3bfd3df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h154ce1733a9058b52a935998a1ffb5e0b0a21eaa7e1d6682d6734ce6c56f54e900fde2be54486689cea43460f50c83bb3d2ae57f8c4c4db6b1a8725ab0f066a7fa8f1723bd132b9d7850d932fc91b1ccd8fa1055935e20146e6e1933ac17ef963386423a981540030aad66d88133d87211c710adbc17e7cfd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35d074e6381d4bd516875aff05bc9480d5019e7d93a994a12a2d304d4b4b22b573e33c7a83ec72b653c9fe72bbe52a9c84f507a034398dd70acdc301db3888256138586b035555b15c9a9c9fee8b8b5e0dd10935ade24717e991a04f60a51210497a9d4759884153608f9adbc556c1f1d4a11d4131abd120;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h124962a29dc353b299c71409fecc7586a159e71890884e584c0139648aa852bbd1483e4b74691ab7cabcef84917c56547ee05458eb73ad892339066ed9815d2e6628621d47128a7b86af920bc0f185916d3d3ef9ab6cbed745582d3b2687855c28daf494377caa5254a1706cbec0b2d6199c5a78032839bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44e65dcbc3293697e84fb0b7c409c8b1644c7bdd6e391755ccbf62f0cdf7dd7facd95b810dc9954aa9cc7d6d7e9c6a57f4458399eca4a09bc6cdc722791cb1a62301b1def1530359a5afa00e78ab8c4ee8017ceda430874f00472d742d860dd84949477f10ab06f2b7ff4e8e5b0ca098ea318dd0866214f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9f842d55b1e074ccc04046bf0b8d674974f111f09999367a99fc410c709b313a924e53923debb318b30984e6d6e8df97f847c4fd947f817ae27ee5671725ee6724e6f1968b160cdbe68e8a5a1cb2fc4a8a6d77442989a3b3c20f605a423ac048fdf9d2ec4c4f9d677d9acb39cf9dbf810b72d48342ec8109;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h163bdc22b35070bba085d60f35a0b6b2e91863a290dfb47ed3c6ba82b4b17ea3919a908371845370c4c086f20afbffee3f91d2ab6ea92c32335c3177b29a8475e54801c73b721ef50aa7dff2ce3e62dc7b80f249c5d98c431399a58002b84398c2be0d6c384bf0d057dd814a979cd1b7bd94825f0cb1f56ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfab6cda7383b2309288f03f075d6172fb0c56e0bdd0f84ff328268280a30e54b4c5e4ba95fd482b89161ffe285108489d127868c751af9b8c27f81dbcfe2206ce3e89ab721ae490ed2ae0ed855b4223641143420de45062620726aad79bb9373e34abe5f28aee17f642193a1807a7590c4e61aa0f4ddf9a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c818e59918c1afdea510a4ccc3a07208244d91b8a95142edaa1228ac7a1bfd99908195485033da9b5a89802e9af640c165483b2f7fc07ad2ab80a699de71d39e2b880ce1c8e22e6a3ef780d449a86200aa8ba195c47c70f427ede0969d9a843d02f06910b443fc347ff18012a91b4e2418ddf342e759473;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50af3c514232dac160233cae97ac37a96370e13cab87a70cf13c0f91a820c3b2d4315d340d2078b07d4580b31f82c5fa0a774a82ac95c0565876a8131bd62b1a7d59d565c6a21f75930f5a344676692ef030b866536a95cec79274447f610999d66a5a918dc3cfefa3dca344ab526b9c7ccafcaaa60df873;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9076a9657b381451d06b603a5267d813e86afe2ba3145fddb76aaefacacbe1ef0a7a55d1eb1bad1f01809ef661ddf8a9b045953b99ed582c079ebe0a0bb05f9c661f17cbfb0bb097bea02d9d7a70784badcf9ae28c6897ee483cf653414fa06b3d5ba0b724dc0ba0a8b8d64ee7d4adc38509f9cb0d23d1a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f658ab71ff618017f39ebb6e5974d7ec8fb94cdb267b74d347ea6acd4959e60d12378af6ad4df429fe4b3f788fa95dcf2eaca6d4d670e322403ce55190b7a8cd404fbca5a5f4e44ecfd93fae199fb4b6f010b35a056039a06cc75cfac0c0139ae16f766e061617499714402018cb3dcd7d4d0a725e23297;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h42abce231cb22e8ac4134bb7d3219f83b49fea4dac56f1a60f7348b48b456113b705932f9e1a406db49305177df3136a183900839b973323c0587f3367e9ff82fb0aa1fe08bef458a8d11b775e17361ecb616934f7bc744329e3cac30269adbe2f0d8355a846b383e89a951cc067a86c78f42cdc4b7f80b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b04dd7d5859ac15f25a0f7a6914fa72b299f420b7f36226f4f400fc9332f39d81e5d961371d750afe9c3aab80e8d9d167a27202cc23fccf145f695135eb0a8c9da4c1ac19ce509395263abf0450cf917d35256c265d04017a08c81647ceb3fe45eed3176f31ee323de4d09100670d801378c8b44b7f1f7ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hceb9a73c98ded11647fa837ba833225668a315bc02371708c1de3b2e888ed3c43beb2d0f96cabdc11b8c2f3ec7e1c56e6bdd2240377dddb2ca83bc6f2fdba87177e7e02a12e3e73c02bc730ff3b67d4c38fe7c81ad5be12ec7b0e1498fdcfd71475dd7a7e436a3d327365a8cb2ea2b574ac90e5f5c6c2373;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha809c731505b99b6ce3da7dfb507d2051657ecd9a51d10892c947323b5a62c9c2278acd8e80f7c337c10ca8d1ed79d5b01ed43b7109374f3afdda8bc3ff0102c92dbb56a7210b91d5a0036012851a729c503f621b81fdc59d3533fecf4ef8ea49f4c78e33d826b41d05c195f3cff81bfa36f649d964e5088;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h431068e21b9f82838c05208362019dc14aeaf79896232ede15f1d90ea764137d791068c1f58572cc7ebc24175d8d11cee36ed6b2efca8c80afa34c0e1a5292b8b4213d11a8a12fe02f93d23e6e0c9a74b37073d87f660afb6367a376cd7c0356599b3999e1a834f350b3e4dd3f52b751dd889b71c2514707;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12f81f51e95abcfcbaca5b5f53a135eb5c391535f5ec6e58993fe1a982144241d4e76f6d916de68a5e5119a7a925b36c557fbd755203f9cd922a7fb67f56e2db4d9694f9eddacfb06abe5bb7cebec746efaaf5a884afd84012c17505d6fa8338ee2409ddf2ee896c3f0a218e27e17486e68635f9220be2cf0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6aa457f82bd3bf6ce69eacaa72b5c5a42df42d6422b4a11ec2eba87be6e5f914e2da6ed90f673e5266b981f8f6c5397a2604b69de274fa9cf5e3f57242386e027e6a6ca7450387abf6ab9669ee8ee49430dd95daf20dfccda43ac9c9fd10be2e35e2fa9f3b48723e7b38c696730158e7c1dbda74c5f10f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h919cf6586d52496a5f084f630c3bcf6a787dc4683039dd10971c36962e5975edd63a75e8f882866e1484a7267087080c943028aeb8f5c095af93a31007fcdcd5ddcb6fdd30b3617a37777e0f8ed9af424a5899ea4638fa59bfcc3217975fc7f73bd0cf64087d574972c01f22a43f9e761b5bc7f0b4300669;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h185780bb4728fb1fd001fb409df0213fe50c2107ca5b178c50c260f5acf3d76a5eac2993f19063a24c7b534dc3ca20f90ebbac258972e88a3511af25b71e66b08057c13c9fb35ab7f7b16276e6e238aba235bac1cfdc2ccb8a73bab3e77e59546236c2bf0bd09039d1fc4359066f1748059c59b006c199d49;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heaa27a485da16c0d4ae98a8522dc6e0b7d28f65facefa27d505aebe416476a7bbba393dfb3a2dfc8690220f5c56d048d7bfb275bef5e3cc8a1be273da40fb0b90719f0c21e57224545d4c2cb262f7bc0e08437c2e9b89cdc55290582167e9794b1a043643e6b8cfad3a1e38b4e24e7f362f39d5440e0b7a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h712ee8a372113499ea7894cf52a0abc6af7f81cca653c40701cab79fe0b9b1478df1922968bd2615e82919deb61d61f0af3136026fb3b50f055bb37e0da36ca25f24cc82062d7ff2a686d39e48a754eaedc27ac9b358d8feb8e1fe2f82ec28bee72c75640647938dc589e9cf54fabf73c533d56e651222bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eb3d5c2a420d3fecdd75a3ceb821375678fec133bfca8f9142468d8327b86b97e98a1c14cce5c44ae1e115200abeb0143e7b4746c5b133b5b1e9fae673513816b88c651d7c11e311f45b689c1d6406a495dcd3b41286be33a946e53aa3fc60fb96b970ca5d3f86187ee2090a8ed33e5d1828c8e0804870f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181f16937d72daf4f635c10a1c4f6bd3cae0d9f8b57d25c43f0e8d8f4ffd96239701f8e906f0cc27b80443ee13163b4d43be81efdf63a15c5164e20b0a52098114f4d877ac89dc4d314fa66290f0b1ad5620bf0b8b8ef8ab72a72b38c4a3eebc245659a92514e2fe02ba3d0a4e04ddf71234fbf3d03bd4a65;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d3365897aa9afc03471b0878a087fdb04f2b432b1beb54ebc958667ddc0d516f57f7a898c15591adc975c3ebe55869372200861e5ec29d5d0d127ed8e23ed5f2440f3b70af2e76964181bfb70100b1e58f0a821c67acb154bca44cca0fb3f571988f335893c3544fe8473ce5c9a20c06fefbcf30f3e8a91;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9779907f3428c33934fbe26b1249012049c575680d5725df905530be3f54e73a876af3e077695105716ea70a6fb016efd70b33f5a41ea85c5020358b5bb9e1def942d8b596bcef9852c8da231e9b13125795ac2603c5197db1056ac0c2855942baac1f28593c6b2639afab77e862ef124124c025efc82b00;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h125cb0f15ea55196e45884e9141d0a418602d9b13eaad1cc2a3836b1e3693b371c93b894eb45d7b6d06ee69a4cc09cf35c45a34e13afd1080121977d5d294a45fccbe9bd43584c3508eb0b6d7b2c6ab60e565708f227a9a7d2df28c1866c1458b640ff15b88a5616e8ac19c01d42f1056e026f40efdf937;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b42c5b49c793c2b8c32579c60ee0fa926efc26bbf43ea86006767173b7392ac9275f8ef292d5bb040790c382fca9473f713b3f3c4819c3acbc7a1e7cd9361c6045afb46c672e123c7ece80b37c8c0bd4ec3c9df5a10ddc85431b69a2211db4d800cb037318f0e5c86e5d8b54e9201a977a9d0904fa65cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186ee47da1c630a84847748347db70db191042970db51670b462747c8d37f6686c223aa58dfbc8f400f67d369f5ebe4edd205d7e2da4be1493c39cc09ad4325dd0fa5b74bf9517ee5c405cf45e6045189a3ec32eb42cce094fc0c47279058d8565618c9f228576789a26896f8c5fe605add66d00dc6311979;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha6c051e3c92aa6fd739a87efe9027e73e30c4a57fa5efd47e15690cc4ff9fa8b29c7f0061a97d65727bc9261ec558d5189b1b0e87df0f0c88a8450f5b7afe6747ccad74b4732d568fbb6e3a7344d49017f20196bace90c8ecf0a4d163d0d546bf6beb4954f37cb2e997b6aef87d9de73e094952327c12b02;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e2421f54553097a1cfc03215e888a9bc8aef08dc6c5ff3ce39ae2da3e8de4ba8d9c705d86bffb3ab5915d8e35069d8eb7ef102857fed69211fff147c75b318e528b8bce41fa9fe01523073d877891e037cb451b69c85ecaad94da6023728796fc25cbb07e2000ca7720bdacb3e65552e3f8c2a010ba8166;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3baeb9dcb27c0f1a9c1649c331d387266e6fe22da9b1d3e7785c7f8b504a1c894b5b89daa79778746a6136774c3cc4cd8cddc757930bf0779983cca916f9b29221a72582894b49b050b9bd8b6e16c14bd44838c3b174aeae3453561622501cfd47a33473cfed9cef9be6b8a880e0c80a979489e3885c9ec5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1acca1ac215439d0cfbd51991ba2341a6b7466afb62b88340892004310455039b4ff92b8d321a82a5d6f9e3910fc6e4089dbfc595773b61c57ce244b90873b2ccbd1bef0eb15de5bcf47706ef85165218c48eaf841244bb828d8ef3c9c936106badc78470a510538e39489bc289cd76b8ef60466dcdb6fa70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8bf888f95017ecb8bc7a0ffcd376a3575513cc5c5fa5122914c2da5a43653bbce359278627a285200285408eaf43fa04fbb309302eb31c8fc058ee4910afdbe4c7198fdb83419bafd674455a5e5c8f2b3b2f83fbb1a3336fb6beb52ffa107ff23b498bbaee46bd4d039c4e9897f4cc24fd236c566c6f804;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15cdf27c278ed92bc4854ea3b68143f157cdbac6c56521d4d0f2b46d1d808503decb7479c593256918a4c9e417e2b0524cfb8ef646af841699a946da0a7fb2bf41d1a5ae738d11d1a4730bc8129d10feeb555a7e66845283ad50c4be260929be03a2bf004e752637e78f88bb85f11fd6af5cc002ccaf80cbf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e9b09a0360953030d8a1a61d749a7d747f1593e0401d7338dce24d0d0776ace766a8aece7409bdac34c59ed961369d91bcdd014ac09d0db35560b0f970126bcea64d5f03d3ed9e3dc17b0dece1d45194e23d2c122f6aacc977b0f659793a11a8b29d1c394cc116aaeb92c1853710cc8ac1aea052f56069e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h41c599b25b2249c76f8099a2e03dbd3427723461b5d2d875cc6479eaa9cd84cae841f9db4add91fc9304a14cdd9a46b9f89043f62c348267bc150997631ccd20a5c66219ab2b4838927dcac4f5fa9c1b68d0b94bb423599ae78d7e6310afa8fe1b272f77a11ffd6a60eac604d4ce00de0b541bdfff10e36b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he84168a1945e4b9308398ff6ac07322f03369aa38374bfafa46be18f14bb325837a488ef7b326ae65f2001eef02dd2284e21606e7e495346c568bafc03374933402ecdec60b4af8b6d14d2525c91fb820dd55ee3b6dd738741995bd38c0293249a3e191b36fa513f49327dea0d28ad5668fffe6a819bd84a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1272755eeb7343f9c19c889084848672e582ceb790ff80a63e5571b14ccae1006c695f41b0fcd9dff03997b950cc75e0db42c90b9da29a509af35b22737f8f7c946e5eca6e9b1afdd044f98d005a848e725f9e1ddf27d8c38696dc586fc244c459ca6c874351d4382dd2cda398591c7d6615926d8e7fa16f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a02a0cb95cc903d2e80435bfc999d0d8482f466519529295da7db06dd88c0e4d1fa90ef849ad2f2668b96a8ebbe4b430a3cdb54070f4558ecacc2bc5ae4cfeae912bd050c8cb6b52a379a27257224e2f2eb246babb45fac8d0cf5accb848320c6ba6cc82d774d4c997ac2b7ec93815d7ce5a4d7cfa720c22;
        #1
        $finish();
    end
endmodule
