module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    compressor_CLA16_12 compressor_CLA16_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15));
    initial begin
        src0 <= 16'h0;
        src1 <= 16'h0;
        src2 <= 16'h0;
        src3 <= 16'h0;
        src4 <= 16'h0;
        src5 <= 16'h0;
        src6 <= 16'h0;
        src7 <= 16'h0;
        src8 <= 16'h0;
        src9 <= 16'h0;
        src10 <= 16'h0;
        src11 <= 16'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA16_12(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [0:0] comp_out13;
    wire [0:0] comp_out14;
    wire [0:0] comp_out15;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15)
    );
    LookAheadCarryUnit16 LCU16(
        .src0({comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [15:0] src0,
      input wire [15:0] src1,
      input wire [15:0] src2,
      input wire [15:0] src3,
      input wire [15:0] src4,
      input wire [15:0] src5,
      input wire [15:0] src6,
      input wire [15:0] src7,
      input wire [15:0] src8,
      input wire [15:0] src9,
      input wire [15:0] src10,
      input wire [15:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [0:0] dst13,
      output wire [0:0] dst14,
      output wire [0:0] dst15);

   wire [15:0] stage0_0;
   wire [15:0] stage0_1;
   wire [15:0] stage0_2;
   wire [15:0] stage0_3;
   wire [15:0] stage0_4;
   wire [15:0] stage0_5;
   wire [15:0] stage0_6;
   wire [15:0] stage0_7;
   wire [15:0] stage0_8;
   wire [15:0] stage0_9;
   wire [15:0] stage0_10;
   wire [15:0] stage0_11;
   wire [6:0] stage1_0;
   wire [5:0] stage1_1;
   wire [5:0] stage1_2;
   wire [7:0] stage1_3;
   wire [12:0] stage1_4;
   wire [5:0] stage1_5;
   wire [12:0] stage1_6;
   wire [6:0] stage1_7;
   wire [5:0] stage1_8;
   wire [8:0] stage1_9;
   wire [8:0] stage1_10;
   wire [7:0] stage1_11;
   wire [3:0] stage1_12;
   wire [1:0] stage1_13;
   wire [1:0] stage2_0;
   wire [6:0] stage2_1;
   wire [0:0] stage2_2;
   wire [8:0] stage2_3;
   wire [3:0] stage2_4;
   wire [2:0] stage2_5;
   wire [3:0] stage2_6;
   wire [3:0] stage2_7;
   wire [4:0] stage2_8;
   wire [4:0] stage2_9;
   wire [2:0] stage2_10;
   wire [2:0] stage2_11;
   wire [3:0] stage2_12;
   wire [2:0] stage2_13;
   wire [0:0] stage2_14;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [1:0] stage3_2;
   wire [1:0] stage3_3;
   wire [1:0] stage3_4;
   wire [1:0] stage3_5;
   wire [1:0] stage3_6;
   wire [1:0] stage3_7;
   wire [1:0] stage3_8;
   wire [1:0] stage3_9;
   wire [1:0] stage3_10;
   wire [1:0] stage3_11;
   wire [1:0] stage3_12;
   wire [0:0] stage3_13;
   wire [0:0] stage3_14;
   wire [0:0] stage3_15;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage3_0;
   assign dst1 = stage3_1;
   assign dst2 = stage3_2;
   assign dst3 = stage3_3;
   assign dst4 = stage3_4;
   assign dst5 = stage3_5;
   assign dst6 = stage3_6;
   assign dst7 = stage3_7;
   assign dst8 = stage3_8;
   assign dst9 = stage3_9;
   assign dst10 = stage3_10;
   assign dst11 = stage3_11;
   assign dst12 = stage3_12;
   assign dst13 = stage3_13;
   assign dst14 = stage3_14;
   assign dst15 = stage3_15;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1325_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10]},
      {stage0_1[0], stage0_1[1]},
      {stage0_2[6], stage0_2[7], stage0_2[8]},
      {stage0_3[0]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7]},
      {stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6]},
      {stage1_5[0],stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2]}
   );
   gpc606_5 gpc3 (
      {stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[1],stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3]}
   );
   gpc606_5 gpc4 (
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[2],stage1_4[4],stage1_3[4],stage1_2[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_4[6], stage0_4[7], stage0_4[8]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage0_6[0]},
      {stage0_7[0]},
      {stage1_8[0],stage1_7[0],stage1_6[1],stage1_5[3],stage1_4[5]}
   );
   gpc606_5 gpc6 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6]},
      {stage1_9[0],stage1_8[1],stage1_7[1],stage1_6[2],stage1_5[4]}
   );
   gpc615_5 gpc7 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], 1'b0},
      {stage0_6[1]},
      {stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11], stage0_7[12]},
      {stage1_9[1],stage1_8[2],stage1_7[2],stage1_6[3],stage1_5[5]}
   );
   gpc606_5 gpc8 (
      {stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6], stage0_6[7]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[2],stage1_8[3],stage1_7[3],stage1_6[4]}
   );
   gpc615_5 gpc9 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10]},
      {stage0_9[0]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[1],stage1_9[3],stage1_8[4]}
   );
   gpc615_5 gpc10 (
      {stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage0_9[1]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[2],stage1_9[4],stage1_8[5]}
   );
   gpc606_5 gpc11 (
      {stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[2],stage1_11[2],stage1_10[3],stage1_9[5]}
   );
   gpc606_5 gpc12 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[3],stage1_11[3],stage1_10[4],stage1_9[6]}
   );
   gpc1_1 gpc13 (
      {stage0_0[11]},
      {stage1_0[2]}
   );
   gpc1_1 gpc14 (
      {stage0_0[12]},
      {stage1_0[3]}
   );
   gpc1_1 gpc15 (
      {stage0_0[13]},
      {stage1_0[4]}
   );
   gpc1_1 gpc16 (
      {stage0_0[14]},
      {stage1_0[5]}
   );
   gpc1_1 gpc17 (
      {stage0_0[15]},
      {stage1_0[6]}
   );
   gpc1_1 gpc18 (
      {stage0_1[14]},
      {stage1_1[4]}
   );
   gpc1_1 gpc19 (
      {stage0_1[15]},
      {stage1_1[5]}
   );
   gpc1_1 gpc20 (
      {stage0_2[15]},
      {stage1_2[5]}
   );
   gpc1_1 gpc21 (
      {stage0_3[13]},
      {stage1_3[5]}
   );
   gpc1_1 gpc22 (
      {stage0_3[14]},
      {stage1_3[6]}
   );
   gpc1_1 gpc23 (
      {stage0_3[15]},
      {stage1_3[7]}
   );
   gpc1_1 gpc24 (
      {stage0_4[9]},
      {stage1_4[6]}
   );
   gpc1_1 gpc25 (
      {stage0_4[10]},
      {stage1_4[7]}
   );
   gpc1_1 gpc26 (
      {stage0_4[11]},
      {stage1_4[8]}
   );
   gpc1_1 gpc27 (
      {stage0_4[12]},
      {stage1_4[9]}
   );
   gpc1_1 gpc28 (
      {stage0_4[13]},
      {stage1_4[10]}
   );
   gpc1_1 gpc29 (
      {stage0_4[14]},
      {stage1_4[11]}
   );
   gpc1_1 gpc30 (
      {stage0_4[15]},
      {stage1_4[12]}
   );
   gpc1_1 gpc31 (
      {stage0_6[8]},
      {stage1_6[5]}
   );
   gpc1_1 gpc32 (
      {stage0_6[9]},
      {stage1_6[6]}
   );
   gpc1_1 gpc33 (
      {stage0_6[10]},
      {stage1_6[7]}
   );
   gpc1_1 gpc34 (
      {stage0_6[11]},
      {stage1_6[8]}
   );
   gpc1_1 gpc35 (
      {stage0_6[12]},
      {stage1_6[9]}
   );
   gpc1_1 gpc36 (
      {stage0_6[13]},
      {stage1_6[10]}
   );
   gpc1_1 gpc37 (
      {stage0_6[14]},
      {stage1_6[11]}
   );
   gpc1_1 gpc38 (
      {stage0_6[15]},
      {stage1_6[12]}
   );
   gpc1_1 gpc39 (
      {stage0_7[13]},
      {stage1_7[4]}
   );
   gpc1_1 gpc40 (
      {stage0_7[14]},
      {stage1_7[5]}
   );
   gpc1_1 gpc41 (
      {stage0_7[15]},
      {stage1_7[6]}
   );
   gpc1_1 gpc42 (
      {stage0_9[14]},
      {stage1_9[7]}
   );
   gpc1_1 gpc43 (
      {stage0_9[15]},
      {stage1_9[8]}
   );
   gpc1_1 gpc44 (
      {stage0_10[12]},
      {stage1_10[5]}
   );
   gpc1_1 gpc45 (
      {stage0_10[13]},
      {stage1_10[6]}
   );
   gpc1_1 gpc46 (
      {stage0_10[14]},
      {stage1_10[7]}
   );
   gpc1_1 gpc47 (
      {stage0_10[15]},
      {stage1_10[8]}
   );
   gpc1_1 gpc48 (
      {stage0_11[12]},
      {stage1_11[4]}
   );
   gpc1_1 gpc49 (
      {stage0_11[13]},
      {stage1_11[5]}
   );
   gpc1_1 gpc50 (
      {stage0_11[14]},
      {stage1_11[6]}
   );
   gpc1_1 gpc51 (
      {stage0_11[15]},
      {stage1_11[7]}
   );
   gpc606_5 gpc52 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc53 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[1]}
   );
   gpc606_5 gpc54 (
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[2]}
   );
   gpc606_5 gpc55 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[2],stage2_7[2],stage2_6[2],stage2_5[2]}
   );
   gpc615_5 gpc56 (
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4]},
      {stage1_9[0]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[0],stage2_10[0],stage2_9[1],stage2_8[3]}
   );
   gpc606_5 gpc57 (
      {stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5], stage1_9[6]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[1],stage2_11[1],stage2_10[1],stage2_9[2]}
   );
   gpc1343_5 gpc58 (
      {stage1_10[6], stage1_10[7], stage1_10[8]},
      {stage1_11[6], stage1_11[7], 1'b0, 1'b0},
      {stage1_12[0], stage1_12[1], stage1_12[2]},
      {stage1_13[0]},
      {stage2_14[0],stage2_13[1],stage2_12[2],stage2_11[2],stage2_10[2]}
   );
   gpc1_1 gpc59 (
      {stage1_0[6]},
      {stage2_0[1]}
   );
   gpc1_1 gpc60 (
      {stage1_1[0]},
      {stage2_1[1]}
   );
   gpc1_1 gpc61 (
      {stage1_1[1]},
      {stage2_1[2]}
   );
   gpc1_1 gpc62 (
      {stage1_1[2]},
      {stage2_1[3]}
   );
   gpc1_1 gpc63 (
      {stage1_1[3]},
      {stage2_1[4]}
   );
   gpc1_1 gpc64 (
      {stage1_1[4]},
      {stage2_1[5]}
   );
   gpc1_1 gpc65 (
      {stage1_1[5]},
      {stage2_1[6]}
   );
   gpc1_1 gpc66 (
      {stage1_3[0]},
      {stage2_3[1]}
   );
   gpc1_1 gpc67 (
      {stage1_3[1]},
      {stage2_3[2]}
   );
   gpc1_1 gpc68 (
      {stage1_3[2]},
      {stage2_3[3]}
   );
   gpc1_1 gpc69 (
      {stage1_3[3]},
      {stage2_3[4]}
   );
   gpc1_1 gpc70 (
      {stage1_3[4]},
      {stage2_3[5]}
   );
   gpc1_1 gpc71 (
      {stage1_3[5]},
      {stage2_3[6]}
   );
   gpc1_1 gpc72 (
      {stage1_3[6]},
      {stage2_3[7]}
   );
   gpc1_1 gpc73 (
      {stage1_3[7]},
      {stage2_3[8]}
   );
   gpc1_1 gpc74 (
      {stage1_4[12]},
      {stage2_4[3]}
   );
   gpc1_1 gpc75 (
      {stage1_6[12]},
      {stage2_6[3]}
   );
   gpc1_1 gpc76 (
      {stage1_7[6]},
      {stage2_7[3]}
   );
   gpc1_1 gpc77 (
      {stage1_8[5]},
      {stage2_8[4]}
   );
   gpc1_1 gpc78 (
      {stage1_9[7]},
      {stage2_9[3]}
   );
   gpc1_1 gpc79 (
      {stage1_9[8]},
      {stage2_9[4]}
   );
   gpc1_1 gpc80 (
      {stage1_12[3]},
      {stage2_12[3]}
   );
   gpc1_1 gpc81 (
      {stage1_13[1]},
      {stage2_13[2]}
   );
   gpc606_5 gpc82 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc1343_5 gpc83 (
      {stage2_3[6], stage2_3[7], stage2_3[8]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3]},
      {stage2_5[0], stage2_5[1], stage2_5[2]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1]}
   );
   gpc1343_5 gpc84 (
      {stage2_6[1], stage2_6[2], stage2_6[3]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3]},
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0]},
      {stage3_10[0],stage3_9[0],stage3_8[0],stage3_7[1],stage3_6[1]}
   );
   gpc1343_5 gpc85 (
      {stage2_8[3], stage2_8[4], 1'b0},
      {stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4]},
      {stage2_10[0], stage2_10[1], stage2_10[2]},
      {stage2_11[0]},
      {stage3_12[0],stage3_11[0],stage3_10[1],stage3_9[1],stage3_8[1]}
   );
   gpc1343_5 gpc86 (
      {stage2_11[1], stage2_11[2], 1'b0},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3]},
      {stage2_13[0], stage2_13[1], stage2_13[2]},
      {stage2_14[0]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[1],stage3_11[1]}
   );
   gpc1_1 gpc87 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc88 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc89 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc90 (
      {stage2_2[0]},
      {stage3_2[1]}
   );
endmodule

module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [15:0] srcsum;
    wire [15:0] dstsum;
    wire test;
    compressor_CLA16_12 compressor_CLA16_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hdb6d60ec0e2d140a3a5ca87fbd093b06e2d6494c0d544fcf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc33e4bab5d236272be87f097af4a0d63d4128edd278fd29f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h2d5479f57983123344d5e1dc7f7fcff0128c9bb69046aab4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h1281df5d0c71da354642f70eda63f9683b304448073b9928;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4336d834a357970b4149ab4d6fc6da1154c70a918de97adf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h7c838cebe8320633ec98036c23c449a078c9814dce43b9df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h8e26101e1663a50056beffe769c01760bf632864ce6cbe81;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h3aa6906150c9bdfe18ec70cbcd1334669cf84b621b81d9e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h42c5daf1a293d35107230ad62cebe454709a2d46ddf59524;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd096b5634ad6d4364b2fe6b17d0017a131a2d00c450d413b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h478430c7f4357cd96133834580ac66aaf24de4fe65c65d31;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hfb95a3c247c8bac1d7b8f75e1eb0a8f69396269e80c42239;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd87f8736cb8a0f5335ea5c5a6c898dc0a2645b49bb35fb6d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6450cc1759b7fa98b36fcd440a8fc52ae42c0797872f1537;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hdc3f8c9de20904d70f64cf30f123161de597806ba4bbdc3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h5a0c0a28c9dbc9ac9e3a787aa96718cad4b1d01715019227;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hecd1408bc582723e299573e1d542b5857236a1a4b77e2f62;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6f9649eee6109ac13e8d735dd8283d04285959e46425e9d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h539006664041e0e1c66c252fd33629f508b0034c8c13a19d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hafb4039f101801087eafbbf37952bad3d7c241dd5592c82c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hc8d9e0abf1548528898e62f6dd27475ccc9c9c7039ef51f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4f23677aa1a4d291c468fed9f8046db84214c3c7d5bc5aec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h68c702235dd4f0ddf157741f4ccfe47366c95b4139929942;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h51aafeb26e94758992a5407119a281b7dba566f9514bd786;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha15e15fc934a77530ade5112999ba08ca0eba9a1ea90ed69;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h9d631296f4bd5748db19f45f48126b0291804fae3fee07d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h25e6994d4dd4cd4c7f47bc2ece369617bfe92fc683976176;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4ed1cf6d24605a3bcb65f010ccfcd9d6db776a0300c8af2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h948cc42b446d638cf6520c4b756e1a2a2d0d5849b29eb8f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hb1dbc9d7306feca479e6c87553106c3293d5368c2aa082c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h3ce4c2c82ddc0cad97247cc0cf2db6c7104688453e342915;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h208fe44ecb38196de2bfaa50a7eed9c2cf376fd0cfdb754;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h42e837e748bcf1501c139662dd8eae365631b5a913d63b4e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hbe36ee1c11bc0db3a207a1ecfce5563d12e10fe870be37fa;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h7bc5f58d9a53d0c35e2a322b68c60804b1eb7d48003e4636;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h95888421496ca284b05002b6e8c9328a4ef47f05015a89bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h32869f35f9995d88b135a2263e6bd5d692688d8183d46e4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h9afb579d2aade91ebfe5c5fed8edccae401ddc935b295f2c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h25483ff9e03e2128bad7cbc2c3130ecf4d5335c83ec50cfc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h18879b98d66044c6232557293261a55b9cadd85fcc417ee5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hec77b3e15b14dfe194bb28fa00766523bb18a329505150ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h5e7f6987816a3e7e5e9ef315e384cbcbb3d6396960af6fa6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hdd2b2ba4b542209799a57ee0f97cd4cbb62875a7caa2bcc9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h2336525c9568199a0256ffebb59ed7d696357360d093140e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h1fd77aaaca08488cc7873647f62622e929c548e91a1124f0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h2fdc74fbc5df6a22582c761b96ca5f1464a71ab19cee27b5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha3f2d2d03498f992ab699f85220c2948bfd20c0c49308322;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h9a2d4a1713a66c05a6eb2c3bd3dc7eec1418de70a3b4519c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hdbf457dc37cf75c436c2bc684c05bdcfea87e692deb0f62e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h199d59df2e7e3a621a9bea2d7d18efc68e0d0cdec193340;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h29b59a7108edf1da61825312a66ad03c1abe47f90e039325;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd5b1111037193bab2ff9a08bd1e25f98c1cad8742cfe32fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hca76b972a40e094b099dcef24f3b8bf451961a86c656035e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6d488acfb432726b89cb7277038030a0715fa1899c8e3033;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hdd18cee9298b6cbf9a47d617d95866deab84657c1f3cb51d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hcfcc4243d373d16514722df4a14b58550036319e566b1343;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h675f02661a557437b355c169688edcf286f3f513a592805a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hb4f05ddf0e56612ebc4f9d57f06dea85c4c2d105790f53da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h8dd95f24d833326e5d1725c440a1621481a016879ced7590;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6e638f8e5641ef51e571e64ea0536be9ad2a5fd24eef3876;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4299923c38a397496fa09521f1ec46d9bbecc2ba8e0ca4f8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h7dfdd770db05bce87b6fc2455a859ef2ba691d6a036f4966;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h68d4863c2f5a7ee8f23590302deed7a53cef35412dbc51d7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd4b7582bd20fd6c0f8a8776131d7d7a9a1799d8cf55684ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6b9557467e7cf9b1d5fa0caf233891512a6cef2bf71590d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'he7c30d0563cbcde6aca221a504206847fedd25bf55e3566d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hae13fa50e6c66e66b3d9605aa06777d2fb7d7707e652bb96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4d22410e6624f4cb3cbbe9f63577aa34b075183182238d68;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'had10dca9956fa64cd368e99daa9a4f3b19893e6cb10c9c56;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h8f61078e35fb0f2fb5f07bf53afa246f27f1cf51580322f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h99fab0e1d798f684aa7a8234003d56cba934e45894f70bad;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hb5f9c55971838048c4ad0b53c8f55e3eec959bdcb6d41409;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h9833b2611f85a6a92a55a1c68db6e17f61de4dd039abfc5d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h480b8962ee2386e8baf3cd697746612016344821f953ce96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hfa44524df9141c458fe02d05c300350d13977a83c6299b3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h620e7af2653c8d47295cfcd1ad9391a25c7d77852cc5b679;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'he436a4579112f9d72b2e3d8e465a7ed2ba4b77a741a6d91d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h26a67c1a0ad0983330bcdecaa245648f3008aa05b9516995;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h9ab983aa179c68f688c6945c3b89d9eb039ca61ed54b90ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h7220a22c4d11f8b878da9f1a76a45011644f728cd0c60773;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h626066e46ede4594e0f104c58c7740412040a4f7a98fc0d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h93b3c5881fe3c5474dc6e60ac756c4d3be58e0b5d0e3a303;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h441e83a96f645dc11a3473064cc01fe64d804c0874391d20;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hea4393c84ed1f5b30278a87868fe14b4eb187edf9fed35ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hff3fcfb487fdcc2340b2eb9dd5dc39ffd426f274d2bc1454;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h9ce85c794a942a935cea28ce479b60bea04f50c1fe7cf5c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h968782f537618f2b2a844892fe0c72a3c384478d947b8e34;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'he35608aaf1b38139cd15eddd7585660cb805bfecf03ffdcd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h4279ed2ae1f626d8104e6bb25d9e2e5f8e59afbfc6520e6a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'he262c33adfc4cbb508289b5fc8cd6771750f82976a947d37;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'ha2d183445b54d2518d9a1a8f78b488a2876b7fc9ee810494;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h59fd1b4eab371d7499bae26bb869ab3ad21640978bb52f5e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h1daa4cd66fe1125910aa9b8904cee100d145483b0cff526c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6c8fde20112dfd050ec4dd0e5b09a8b9be3aa5f8cbed38ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h6095e0df685cce2b702e656312682ac49029a1f23560aca5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hd3b9297becfa23f43b88bea800358b1c0cd1ee60cd060478;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'hdb0899e23c9b504f746e35a4ab401d95844fb2f1c0cf1751;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h1b33b06af0204a0d67a62a78535a264090f59530d9ccdcc9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'he1a7299d484cdbd69ef77c2248e2831c750f3b0289286c33;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 192'h67ad34c199773a9607e3e399c03fec0c34d32a4667b801a6;
        #1
        $finish();
    end
endmodule
