module testbench();
    reg [27:0] src0;
    reg [27:0] src1;
    reg [27:0] src2;
    reg [27:0] src3;
    reg [27:0] src4;
    reg [27:0] src5;
    reg [27:0] src6;
    reg [27:0] src7;
    reg [27:0] src8;
    reg [27:0] src9;
    reg [27:0] src10;
    reg [27:0] src11;
    reg [27:0] src12;
    reg [27:0] src13;
    reg [27:0] src14;
    reg [27:0] src15;
    reg [27:0] src16;
    reg [27:0] src17;
    reg [27:0] src18;
    reg [27:0] src19;
    reg [27:0] src20;
    reg [27:0] src21;
    reg [27:0] src22;
    reg [27:0] src23;
    reg [27:0] src24;
    reg [27:0] src25;
    reg [27:0] src26;
    reg [27:0] src27;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [32:0] srcsum;
    wire [32:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f93f9e355ab8aed9a67c35578368b87812d117fad4676d759dd27eb654c070ff7e5e3622b76a8692db92e5470551e0ebde73f61aab836ad60e50352ac720a9ff5639fb65b5e2073dc24286b7443cff73120f0beb61eedaa7e055fcf8eddb760ab51;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93fb540b11577555be5436b1ffce6995ec740693aee99375b623870bc3fddbef534eebeb0809f9ea26b819d7fb0a55bd6e6f5806c2dca57d44de3ea32515d8a7aa6436c99ec70d37382c14d6debe1bdb3e1a2f1ae4e037dee89d7f9fb210eee79d8d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hccb0c12ba62e882ec7724450e9a728c4c32252bf930a159c4dbaf255abacf18df5e5ffaaea9c3a9e91e436f92acbed01c2d4603093997d99ee06c5b8db6fde35697f2b6e665fc8c1521235878ee272624cc0fdda8a1650f8c881eee17d8ad9314878;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha99b3c216ddf50c1b5ae5a98260b9ee38cc80ee032d1bd1683e0c62698c8f905a997dd6efa2c24e1288be2a43076783b893cfdbc63ad5922654308bdf04747407f9863ea6f618ae833237ef3b5dc1db822a9ac40918c5061a87998efdfed7daa401b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d417dd39bcc2fe8d0b338c2a1ca6b171cadd7998962ab1c10c5ed35f032e0a72ebc74681fd42d73399fb799eebd8156378943b9432b61c992fd53a4f57972e435ac2f2478d596f17eb1cf1af9adc2ca6ccdacdc7c9336b771367a0123d49b6610fe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87ff91d3eed42d1cbabb6104bcf974b32d56cee9bb14c87eba973688801613a7b355a251b9cd1f04c2e4c87133cc25c681d2465209da4c63d0aafda922c5efc8342c8a4c429716d459990c9e47b51c6bda44beea90d82273e3d12422dc54cdb21182;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22687417a366714ae2f55dfce41ffdee7e9cce33f88d7a0d10f0042d721d06b238886c57c5c0846177acfb666fea1c1a95362141a1a082e553dca9a37a297fbb4ca1c27a7fc75cd199615de419ef1795593b19208d26e32bc220aad9df9e0eb3c747;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8145f1c40c84eed1b3430665be41a32b9a63180d0cbe461ca4bb210a3085fad77e2cd58dc35d85f8ecc5b67938c8e238fa2161f1330cd71a3caac5f7adabde1fcc0c137ebc4dede6a1059b53bb6ecbc156d5048a2bbb26a60b374ff93e3af5dac86;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4b5344e865b1d740cbc79f245e590892c3dd4d6f99793405c8e2b6368e39c8e091df3dd6a9fa5a387ca8aca50873c9b11d5f50b43e9f865f93f97297a3e42bc0b3ad5b0e78bab7f82b7b1f80217d00beb2a963a9cfb08710b0cccfe85102a6d68c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hace41a5de091e33be3f95c521c4c944af2aca9fdbc55c5bd8c0d9c9869963e74a40edd7e627ab277e991e6ad41700f282419396a8731f989bf65847a3ff0f20102ad3272f02b24d69d10091bdf886bd8faeda37ff7f9f6436d2b32fd756d3cb73864;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8cbc49f150444eb71c86a0b27988d41e6cf52a82c267f2927a866df90283b5539dda64b4195309354768097934b11d4bd437d73c341731e78c07773bddfde823240a9296bda343fcabdc0ad0f58121697a29e3664752b6de2c6d018090580cedfc5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b01e7d0767b84b581a4b04aab81419991cc44aa70ca20f88baef0f4425ffbd224393b40c6c3200880b1270137162603b3aecf424c8c455378537c253e44f4b3402724ad0ea786aafd1df7bfdfb88d62397852f087142842d2b8703cd896561a4243;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a5fcd2fae650b84dcc97e1253cd8ae3d51be1b9ecf935f4db6e2912aafd84015f00288ee13685555349153791035b2ff315d88f63a0e1a3ef7e8a5a8349c855a61042c137e19c443cf5c62a67c9cf61bbd5a4025dbc3458a6840e78dc66a6557bd8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1adf8eb1c34144b2d86a77606008b2ec0aadeb84eebec24e70a577dfbc11df34b33c31c4c2c88722729cd254ceeae2fda90d61190fc6f9269c04dfc4012e132166216285bec2d63d96249bfd4797a4ff077360054e26c374fc45873ec2309fa79e19;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e391f015f6065bd4cb147c955ea099164b3a1ee1652f6e7432a81a0ffdf8b1103afadbbf469d5ad97fb3a4ab0c2083cbc696d13eb502d8eac844ffa3a8a282a3e9f70ed94b54aa4614b56fc089262ec25d89df6dfaeb285f28dec885d504865face;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha653cd6d88c239411dbac65d3418c6eba413c86f08d0114d61c7a8a1afd9f73b0c3bde0c4c01fdca1732aa4e9e7ee533bd743edd8531e439324e93fe01a1265a11592e1f61daa06120f3092765d8131bc1836ef6fa05e2197d36f0af4a985c2a2ea6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5775691df27d5c9a24a4295c543b5a6ad87b4958c998dde5a641fed983bf8057dad140899575aba5f47553880d9593dd7f8d082b5c5aa359c4230d457bf2999da29c2254cf9e1d7f8d6278f4db401e992716854f76b2a51143d4833657e84f0b5ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bec5272de8f12187bba3120441f708437bbfa2c1bc32535e5a7ecc0794e338ce34a471488ffd21f30a3bb215ed906f36a5706ff02a41e426f5e27db4f6c94315f9b99566721c3ee4ca4d325e73ba1b865a63a3071b643bdb8a82e5e7655e7c1c92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a4fb688333465a0cf826893164337bdaf0806331208e75dc8e493488d94d5b437f3a1fd8a89bf37680c504b3e7c6ceb72e01f3822095f6b8810ec44ed57ebfe96398538a4bee50cdb27cb8af6c831cbd455f9fe189b503e526506886957bc41e50c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf16d984bcba99ee556c001abf90f7d2d0f6b5ba5692c3a3f4e84655e7f9e49abff922ad2a7cdece4a19536993d381e2e12dd26a583ba33c488c9672ea83c09d3963d278f27530c08425be753b43d8941af1a2f9f7912cb9a59c922c28d9f030cde1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha62f6f144a8fae8e84ee85956c7ee5b494b9041556fb6ff59dc1cd4fcaf0fd75d4f87531d8fea57425294a89c8e375898155b7213ea89db1c548b6342d99c5d4b9dc04a58d58d0427bc939dbef1ad4f0c6fc84fb0c71ecdd9ec6547948751a222cf9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h528fed219fc943b4624e11fb42b8103b24be09dd3a5cd0b77deb090e1d7221edd24222465e7b005cf17f0e88f7dccee2560bee0c8196c71450b9fd42ee26021082a05cb1a8ef758401b7c69de43b4536cc0c0ab8c539af29c4ce75f0a9305cad0fb1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfd61cc9509632df5961c3f9947e771f81fc01d5de7a28c5bd08c1adb1222e9ca5814bf5e9acdf92c3ef25ca664484b969afea6ea18ee24efe115568dce32191cf3ff78966dfc6e4f64d4ac344f6f88be4fd357ecd2cff499c89371be42e176568ac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdea6f76c31bfcf59b341a52709f938d41a53395cbb76d2b929061f6601d885394a2ccfd320eb0882158e85b765c4311be985de03a32ca14b9f8fab28471121911e32afa5ff6c3f97133303c55a73f55f8ab9936d84a082d2eea8512a8e1cfad5d174;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39600e2d6b2f6333588a2edae3e2b671f5cb03fdfc403eb6d896e5f8efc95617d2e4b608807dd2d477f9c1ab6d52dbb09238f3088a2a0cef49da5c1d136935a3885c225d84d1e8f510f7e177748cabf97a68860fd87640c8faa25028e1cd51a60153;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd23c710491e23a229a480965e55ecbb13f4a73e7655747d3b0372b9aa576a6c7eb376a894e828619eca4a0b0b0484f746e415614ea5ba272d124acc503cfe251ac544912c2a7cef71a43a747211d82e0e3bb93cb114903fefed1caa398d63b8a803e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde5698b6f350d946e314961e513ea5e4c711046ceeb37b2930cb436e9d543cae2ce28a081c6fdc2b875ab1da2c18378619e78be82e2eb805cc9304e2635e3a6e014f2e5305769fb1bb2c414237d7dfcb38887b126e20796d3e1cf3adda7ea7be44f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbdbcf4816344bc78b8ecce3393ce4742ad9d116ba009b84e1bdce7e8a71777f828b757e12b8b3ab260fc09f7e18d4d1a8d817856bae3e2f0451d9c485e7310577ee932db48ed166767acd6d57f90147c7b4b4d8cce409199e58702c36cae2f18df6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd79ac7088c33f3b60768f7f79808ae19fa75dcae57e68291287ba0f37cf3c1f4085b8d2b6509cf652800d5016026f13fd47dbe3b469dd7363fd99bd805821e2c5bfdeb928527633d85974c4edccc1e4071a51e94f0daad6f4f83e8bc1d853a0359f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d25d241ae7b0f06b1960a4d67a00f6625979a20e671687d8aa317dd25ada757bd536df7d8fd1088654c306ce7b2e18076a1b52cbf5a06964a8dc1f78db14b7438fe26d2d7033037413c408f69b81e9a71833f070d8e9815759460ac3d7b5ed30041;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h446230acc91d6622421610e1db585a7e6a4b71f2d7c98233affbd2c862c8ce9d0ef72ca161ef573a1c57cadb450843755bb258337b61b1a58ea63c9b18761cea515dd4dd8abce8f939eaf2893b3760c105af0330a4fbb63aa95df91bd39b0d1736c2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e519183157328311b43dc1ff6946a87a25c5dad3a59383a98c1424edcbbbdc482ca088fdc3b52eb885f42435adad5016d5bc5eebd3cd5217bf97953ea15b398837d9efee4e1a06c561f3d7497eec3abd6f768b4f2b5c1ba9ac16dda73049ee39fd8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddd6e99a91d719883beaa6704a8d6ba7e67bc3b729240b9a160423082d78845b2edf315c85b1055e8c2819d62ffedf8111542c112f50983fb52b697d9a0c6dae735c3bf20eeeae46247ee019f2e8e6618a75656cff4bd55153ff78c77eb999b6e010;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1be1510aa57bf4f116a7604727e59339561d44fbf462b9d0d39f50cee6a3a0a6e93719f205b94557045e8a8520eaf2c90642670c178f44640d85a9c5498dd6e26e3ee33d6331b8607121903a2ec3e5f6eb6ca9df751a8dc6fe58804626aad8a120;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63cf46ca5df9a69db5c59c557045ec234dc38403f507bdf38eab08bae5a993575190d9689a1ce2285c28e3dac641b868cf65e8beb0b0c0d4ca3e33d5fb40caa5bcb780771b21325797fc53aa801401fce85af88e1a028ea3fc35f226555b17e80920;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a09faac8484af8f6d7e1fb7f9241318f099a7cb433dc98d7096fa9487ff11d0bc9b7329364b86fea3c0298624ad93846f70cc2d76f1a46f98cabd51df07022b93c4c951cdf6a8a8e16d738497d401d7fb154827feebabade52d2af14b50d1e6a5f3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3bcc3e04a5d029b020c9b623f6d6a99a44004dcc5aee6ab6deb8982293b538ac818aaca3ed4ec3a6474d5f04be42d2c5c79aaaa5a453df8f249a9e4edb8fb6650b31c4ae0f567e84c7720b5f672d0878b19c2cf87e9152e2e2c5b56a8dad95cf54f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b9aa8670f150c2ad717600a1ef992e4209956b859053be7c7ca96c29e861e386c2583fd2a3456d00b78be25e792d31010fe691e300013f3ceeabff519f0a3f97cf62b647753beec02fdb1af2179d665e8d951d82c7601c86478ecea7f32925d778a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4bc0dcaf260c1c81d48d1453ddf1735f6c4c864b613258bd447a6746e5d100964048997b2e8bd9e06ab43cff2a7231a2576b4ee594c1e5425056032ac22c25db3ddf57f23c76c381d534a872466c131f9db8074985da2444757b6552b464817a52b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h161d2db7c2c441219fb45fb7461d22000710521d543234b8042c528040be0dafa05ed6636c14411a7146414a0054122cebdfa597d86259004436fdd32b3c6416c231277b67821e255eebf60960198a58f210274626a289f1000365068c4e925d7e1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a474d026d76f66ebe63201e09bba9060c82cd660e01c8dbf23bd71969257501a99117f5db0fd694e49e5a710d55da86ce0b0ad9783abecfde4257d06cb1ca4108baf63b8af00ab9d890f617fd4c40d6d622912fff769043da61bedb0713113fbb78;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e710b020c2d423337977cf9800ad7246a4ba5f2faa051d8f55a994a033549f49d3a06f800003742b2bf377e32f66ea4bb9b593cd94a9c19320778393ec0d1f39ac65a18f8fcc78ed32e5ad8ef18bff7d6a947333a94ceef6feb4fd5a9cf6a88979a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0fdd1652393aee7dc6d9a72f34488146e6b7e36b5fe34708971b2546e3280a7173a088bf587deed04170411bf6794b4b0276a9fb78a986309f0301482483ccdd78a5a9ff063a8754276a463c9c1a8e7e4da5943edfe5c693526109fe35df8dc7cbd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd15961492943fcd1d81db1184043f9b61cd0a617266a7a5eab4187eae82e297e7605b1d8a617a420bf090799961ff63df6e612a2a8fa289e62f65e68c1a7ef2466c05b76ca44e335a2e4ca592d770a4ca40242ca5543c134d8e67c086c07c151f8d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a2cef60af9361fd870f7d4bd95ca2aabca44302dfc82a86cb39ff7328f69538294cdc89e20e01f8a6c266d0653c49e7bf5ce16e744955f40047805852a449a02c9441e49ad873fbd9964be1187e3c2d824ec9ecd90003cf50bbe315efb32b300ec6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ab3ac5cb3d22d69028be3469327988e31a7169be7eecd9da38542f3f6b78a846988725c742ee44dff301db79a1a0995f322c23e143e6221b3b419c88fb1ee06e3e48ba9d042b0f49a6ad27927ba8157ce829f9b697beef63d28e689d9c7f6c211a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a6daf3c73f363c43bb44e287cd7716cfcfb4a47f9b9901f736501422f4f28e799d3856c7f52a6a24f64cadad7ac051674c5b1386238acf1f4ec7016ead182c49963cbe2f26e9c6acba2b0c1f94fcb8c4ebf912eb9d5c4d7d7dd5778e81a65965899;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a2ad9ba7e6655bd97a7f52ff1089ded91559a4bc5a75c97c0dadba7a2026683dfc3e91d9fbddc1f378c6d7df0aeab758d947652b932547d45698079694136a21f0dd23948bc56e6a4ee7d7e8a301b3a8ed8b297fd16b3136c5b1630782042086a4d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f58f360d293b4fbcb1f6db88d971192c525452c701a57530c5e594b2de305bfd49e67efe4f1a2b8ca1063a0de1419925527dfad909fa4560133f675bfc33e9756e33b50ef6c6ac268eede43429861450a402de94b0acafa33a78185517a93753331;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8e52204edaec9404ccb9270f333ef2239ea61f27f0252e59dad9e8b67b13e62bcc097d80b3a3c9613ba00250746d357dfde5af988d6cd89cd95cc34ddb919480c0aec52d6c922bf54ce9173cef544afbcd72b02dcdbfc5d45370bc7993014fd0717;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h349447fd962dcc58582e58a9a0c98fff43734a1e761fcae8d8229656cd24afb7a5d079fa5de9653fd35086661878867bd367c0ac833d4eb3e9841d0d4085d11d49ae92253f920ab7c3d5bf5273748178b836641113117361fdb6ca59332f026bbe64;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c892905bcfa0dc2b534b61a5ad0c9b3ea5341d9871f4309d3e63b8978d60fb18471e09a309680738252f56c6515fabd139a5fde6698d3c369f805426fd5df336431304fe5361b7cc6144c66f23d4e36ad099813aa2de29c6b7255c933b2796388ec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h446ac9d816d461e0dcddc638055b972af0b6d673d9623f8bdc2f0c80e1a60814d5ba5bb36fb9ef1b255c30371cfc4e72e4b210c24fa72b0ef4f61cf7d6441b511bd99fae97413513fd4c5bc443fa9173bb473e3b7639089a5407e7c598b48b26ce12;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b993b8d06998735b12362339820434ea43b46a6e92d7f01af3984ed455b1f52da0d9e4443267dd33a57b1d2b4acaa38056d0b2e31db7dc941ff0f82a732b2db0126230f7ac1fdc5071835f25d5813e14b0e385c65f2b37b683d329ccaff4278e8e4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2bdaa26f1b32770c2a89ad3890450ebffd25a857a31a3787a550fda1880e4e37eb62c1f7f97163cf71a5b34a4dfc015f9fe31d247728c2791c165131983a814e0f69e10a79c7a34f0e882b3a1fb25009601dbec4e55a095a66ef4b7083f0853cc91;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9bea7ae80011a556aad83c855c1424e50b5e4788c598d160184435dfb8d9eeb06433143eb1586bbcb771dfa035067e11684da77b603bf1c0135e3f1af73c9e93ce18144e292423704177693d1394d5142a4df29587436c42e213bd7f393b8f6f033;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc315ec24b87f9a47cadfcaaea9efdc79d1e6ce6c9ba43a47c7f3d8b1de1c883fe81dd1453917dc845ec5e12197c556c86d7c939e5c1943ef015f844ce7bfc7bfeaa245c083493a1048ab56a9c689ebed520f346ed8f6946ad85fab4b36f6dee5ec6f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa2a560c80eb8ca05664b86362fbc8aa0701ca3f278532c61df6dbfed61b84beb9ba7dc43898ee2b3e0aa2e05a97838c42e6ccb2d9316563ac9afddd9b8cb09056a48a3985f6792b956941f675b218c9b86af7ece74621a1e5945403f9f417de34fb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0053ee9d9ab4841d651abc551b3abe5d30e5f825d1f6d373161c04659fd1e5146f9a5d0e9d5930a0bf804ecc1aeb70cccb67c9052dd9c82f43aa5f49e9ad630107cc22309e2df65f825827c9126a1e2612034768e151a434cdcb4cb9035a5ba46f1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1bce68d0a1c3ab7e85e68c68f92dac7ca75e3a2fab6dc17e28d1e3bcc2b14874023edb68e9afa2ee030abcb0a77afd07e53ce92d39440af2303b9b534167194d12ba6170f0c8efb49b8b0f405fdb4d461e9a98916d438cfa1d46f91943a66de2e5b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74fb6739e44ae41890540309b98342b0b52ba7aed5e768f062509ab7e14f0f7ac69516a3506a311d4ce8cd2e334790f37343f14935e864a599d226a95ab48d606a592548a730ada69189625952cdff70962caf65b5f882fdb55e0c695166345f0653;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf466eae2a3efac23072a78d68e0ee59686cb5290c18b708996d9560915b5694aabf515840e82aa4ac72b47cf93fee5e077f440cfc74e1090926ad387e8481752956672d2feb7d9c480e2d512a3e415583cc8046b734bc94a477ff49ab8c1c8059625;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87e1a8fae7ef7714e2f8f402842ed4216e84858113f5f4ad38ffd94bb7a7fea9273db789ce97fdb65bc501e2c5be2269a1a97664a78786874adac65c77970b1aca114c0c37afdd6806f262fc87871d31310dd0d9a622b25130a4e40a8be6f25ad580;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9dc9d22ba96f0c262d41ce770efc429c0fb962dd4dcb70fed6f9a5e156f3b15cf16c22e5ec1212e884b54a7ae7e0365e29b8337b2f1cac2ab2b9d8e72f131fc46892f2f013f7bc707e2be8a0d7a1d53e16a4422e4b339a95a70f53f40dacfbd92e74;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a1bbc72835a3ede85319a6efbac8a5d2e3ebf68c9ede5542703ceef4337a7d2aeaa9b05e529c4eb3c33671be08550cf1fee4857919f822607f2c20f15bb364598de193da119af4ad51ce1a5c1d8e172ed76e96b7ad96beeb3c5eb37de7c763dc538;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h894ab155ad6ee04ae1b317f63fe5565816d6e7c0875d1498ef4461d2ab87a205857aa955b172fde8b35bf10e4c2880ea38af4800c081a05686f25213da270fc7e8dfafc3331348e1d7872c5824c36ab2f4d583dcdc8196bac1584dbc936c99a1ed61;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde8e80e5e027ea9d066eb11f760950bba1940a60a2185649f3ecae265564bb0a501e820b46c9e76f687303c969f50a7fc242d78fe88a3ece291a45f8736326b408df58d05c87a0387403ce779bfc5779fe11bf8ff5be92181dd25d330a10519dbc86;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h411621b857428ff1bb32f33f9c4913faefab21ced2fc657b4087e44547b1dcb73b729723b3f26e6f11c8f1165edb434672ca2b2093acd06ebdc721ac7fe3ec71c60c600508dceeaebb9b5559478c1ea07de6eb671f44d1e54dcb0d0513829200817f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea6d15f7569bb58b138cfeaf9e834a79e0e2ff892ef8d334b14b0589778168bb66edb4588853f1c6da19904f4cd0ac29ceb37c115ba7ac0f2914cbca79ba966c488182c85c9877fd92e4ca0a2d3631a4c3b146cf68c006632efacffa042d31c23644;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h697dd54a216546032d8ba12ccd0041ca7fe181ab4966f753cf38aab7b0eb74d6a1113f919a91ee460032d5f60eacff73dcdc1cf49696a949d82ffe2cee3cbd8e69d79ed8350fd2297db5845d47d2cda82517cd1f4ab60522fa29cf1f5f96667df1b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c2fc0ca5681b373a36da86138b1c88240e713f11f5a6e3db683072ddae6750741b103bdd16a6799232129146683acf7fe2a78419d67754b58f6d8285a8f04719b16b5f655e5166a928bc234d45e3f3412ebf10c46e80871678d87cdb2fd2ea7659c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f885e0fa154c4da9dfe78bfbcb958401bd556b96fb65f3d75486f8b2c538e39139e7eff4285aa9406f018e1039a6c37f818a41fa46bce57001523e311e4caaf16c63e776a1eb0ce5eacb608b4a8e26403f16e1fcf9c04ef9601b9e50a2756d8dacf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc615e4c9018af419ceda13386b06be411b8e599e85abd8a7e9ce9ba2ad5520e810cdeedeca0f6a5603be2de06b48231aa03b680cc85df080e5e17031f94a1b8577e1435b6fcdf6ca6dcc44c3da11fe3a496d4e96cf2ceff2e3b19727b75a6dd9f57e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h645b76f2bd99fca5a6d2a532d49832c27f47c8ee494a3eb43a24fb68fd668d96c42d6986487086b7d2cc4f8184c6d5fe290d2ef6ed1c2a75ee692619db4191c051543fe0cd1a75a0b3970e2dfafb0b739029cab1cb63e10fa8e2841aa62fc282c8dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4d64087bede193c2702ce0f03f3c02d803c0573b490ed80dc83a44e80faa18718a3e8a46719706043b89ea4f822d58b47090cb6d6c10b139806918ae906f3774274cbafbf65e0507261d625b9a44d8c9893c16a6d356ff71a35ee63f92efaec6005;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb68cdedadebbfdcd84a3f19fed5065a114e2b29c94a35c7690ac893af101b275b41cc56aae6f244d76fa99b1dbeeee8d83a58e6634a91c734dcb381e907def86becf997a296a2905e69ab92340ed138799f7f1f24d22f3ae9bd6de76df20dac56936;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he42d23c67bfb62cf8366479dd9287735dc4092f84a0cde446e0e91c7d53c4eb9c5811603b0d1d9cd34c7fb3be5bdc5b1951fb9a7bcfc8d73991451c4a5a7cad178ed0adaf3758787d98b4a5a6546d0bd5e94ae5ad7290456f90515c00c7aada270a8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5482a840fb278aa354484aed43cd3c595992d91a6956da2793d6de3752e31cc06282c33b90e28e5b0b12f4d11d92ec5cc3139c702de06ef0f56df00c07304c049ad1d817c58b0d92b4ffd221f40e61d5c9f9c34cd0bb4747d4538b4c93a67e8f2cc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5758d690330fee55214d923305b1ab4c9e0bc97a246f742d8b1ad981ad1f86b99168a33bf1e740fdc8780c33241da65c8fb1d7b0bbcdc105c6049835f151b6fa809904c26b3928a15da294dca121b0c4b139ba379b35d78b00e21ad49ff291c41ec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1598711dc56fb6c41846c18e5814d44014569ac56d6a6ce3b2ce59ea4542021189675905487265bdda81a6731d4e98b7d287e6cb036952862f132102ade58448bc4bf25c279671eff360becc687843b9c1d7cec4b9d66911562f8f5d3b7cb0744dd3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c1967572da982d44939515b770cb3c2fd88b2fe636b30c751c823e6d6be4c02190be424f49be3d5637de36ed669d5b218eb310811a0b7e124e61cba36e9fc4ac1ab1c54ee93794405768460ec560c71ba827f4d0998e3d096762d62c007afca0aac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29ba22d62057f4f9687bf85f7f884a22dce4e1e4a918d655a883e281f73214f1df12701b7916da1358f4debc5921165d42de45969472f490f9525e599c5442773931df898645eb95333b2ded3d5441967077bfc20d495d901c0d757981e067d8acc7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h341a47545b5cad01bb1807420c31d8e1b4e1e092d88b8cbb4968d342b1ddd9bbc0ecb2ac19cae207695c405473f9c6f7db1967daaa3c80680cb1c3f24aaf3bdbf360f3e3777fa7c15d7c9691a5fb501297fb8d1919fa5b8309979a6a0acb20a464ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a42db4fa42289fb3dfdc0bb74f94ee98dc29510a672810d560922a4e4ace3ae1b46c282bd7d2e91afee23df0df0fa010b3d22ea9d6ea962f6c0e76a9b4019bd22ac80647b40124a6c97138a112bc36a0ee3ed6a30bb240a2c4b7b38576720a71e9a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb491462a3b7fd509158d169b1f8161311bc6d667eb694ef96785ccd4310b384cf3822d0a95f43664dd9fba08bf6576405147ea9183b591e564a53adc2bd74fe843c262043f1ce1f1b5dcfb46e562207f7c7d1c083eba34d6f1e93bc4b682f54e273;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h753408d49e316bae2676173e33498f443b5cd4f8e0935d09ac3b9e427eb3c6a730a5e9dfd81ba7c927d16ed0de573f8552469b139510ce7bdf9e6a205d57fd7beb039f3d1222d2172bc0baf5610773d82d8260dda699da6116b52b73bb811b47c0bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f450f0a14876096f179aa8db130507de092be9f5691310850a540881c0bbcbadc60392c09507a5f3c3ce32ee377b56f0a5279ba65482a9ccdf83290cb990030c3968512c85eaa41ee80182c89c738e933ab12d8f6acd19558ab8ff42e1303b925b7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84aa274ea64f93f1289deaffb428c24d192ac00a7ba80305fa7dd533fbba4e8356e16911787e6ff9211f79452c97831d7628c8c643bf45e56c698bc455e9b5ced94c2204d455e597ee63a9c6af8f5e28d1d09d5054bc7f08930b88954396595878dd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f39bc8c2de2860c13c8a873dff937f243d823f273555b62aa27e16a37edb7e589468983d6ff0aa6ca0138e04630c52e3e6a45447dc5fa95c9a4adf06046ad708b9cb565b0659185e0bde816864959eab719acda9dd71b030076aa1471b88aa5659;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92811f435636c16c528b2b956d7d45480edbbe746312916a6d1cf153f4cabc0a19501b827764a032507b2bdf52a16b0e3b4b5999b40363e65188060ff8fa7ac6e23618f4ef289af8b81b213df271abd3c9f4b89b514c4bb9c8dc46d307a411daee8f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb313ba61e2b4cf7725dea6c6d243a3f8a52b380941525fcbbd805d3e1407e635b7df1bf9b16287a7fc8f6feabd984dc1727d8c6797ce7f8d2a6f026b3ba12a4d428a049dac862e0a4a3859ff65daf5a61886cf4a231fe373f02d617682878c59dd36;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7f565e63ab6de2b6bcd8ff3c4fd9feec4eb810b4120a3cb2439f84cb072ee1ba9123c5f2287a37bbf978c99c4d1fbc91a1808fec99020eff2127f510156f22b3946071df2cfc60ee17ce3b6a1c00cd48d4d1dbe57d3170032d6aecd32e3a251b01d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae6b06a4ce591dab1a052d611d0e834c25f941e9ac0cbef27c1b59a8ca21b2f01cad93e44324fa162fa57c09c4c5e6fc10241139c62e9c8634afdfdc809b861b4f7b708042246dd6eb8f90467ea953c1dc85931b95153cf8335dc6bd08942b05cf65;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7a205f143ea474dcdf7bc289aa2e217c1ed2f3e01f6b69ed2a3efea544ea23d17e908433b8d5c7f2012517f31c3ab50cfd2a8acef5e4aab8c8fced193ca73527aa67efac5068664d0b02cfea74c724ce744d8605005f399756f3af0c32917e61a34;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75b3722fa36d2467608c383b69b3304cd599d5760334dd6ede4841593409e3981bf99bf59955c75aa68e67e28212bebad076f774fa68caf46fdcfc4f9f77b38f32be7d00916ca31f119ae398fa06dbc8a0b68f8ad3a17b170f9bcfbdee0e66bf5a9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb6023e81107d353dd5cc051fc4250072aaa4c6fdd65116f698dd5c9a5648b9e243243d7454f5e325a49051d58dd2ec309feacce604ded6e0ffd2d9617b69be739be6535c320668ed28e285bb59f5220bab8e719f161f5c1d8006eb65c0fdd6ec435;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h438421ab2464e896a35779b5980f867eefe1047d4c037f89f0f43cf44f40c62e5bbd081f011214b2230cc2f4f1df95939d1ad5a7d22b14c20845528cf274e58ddfc3d164ac89461e562d5bc81d09bc18aa050672deff79db951c33a245ffc7f0148;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75256ede8a7817aa5ce9977cbd7c5a46dc3c45f6d18b02af73a4c722984eb78d8c70b7f07aa1fb305ea5a9b727f0ced604b46f4881f7ff71c47165c1b8392678ceab3af86b62a891353f07a96e01dc81188bac5d31a8f2c71718874ce9a48fe406ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcea2c428c9e949fa9be505991f1d4159c072706cc242ab8b3d472969b46e3f8a692f859995b1486c58be01b200f8d82d3c55e64a8e8ac5681087582005042f5359b9a55744d4656134a17767abc8160c93cc4cb4bf3ce815707c5967f70bfe20a34;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c85ba4f8614a9f7cc7ca5920601782301be18ef339904916a2d29463aaf1e20ddb5d98a79fb7c20435da292531b65ec30b4e73ed862826234e30874b46d82cf9f7d3f0406f2156a984075a5ff4dd47c746fb1de431240849449cec63bb88501c9a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76246b91c7788092e949e827665f726afbc6ebeecf9f0eb18e5087e30ccd76e9c7f6aa51cd0cde13df2e3688299559124eb859113fd94ecad4fd75e62555deb245a3c8da77f816b5f3f8cd0e6dcdbd63ca5c33b6299b6cd4035bbf76ca5a5af4a781;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86d493217729bef81194cf17142d2fcbac31262fa9969d8b54193e0c1ad786cd370b193230812522173c2c82f2cbd9d35e1d679c6fdf179b94c0af8b801369edd04cb8309f53629013b6a0029a59fd9b24e5e73beffcf7cee867c5b775c988476bc0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h275eb39d4dd3f8f8895008df5c2876ec643d4d6130c44636db155a3b4d9149cceb7d7f34d1497ed93d3381b764cadb4bfaf4545c36b7954d82a61902d46bbde9fc35978c817b49590d8b0bdb402beec8d204c332ab8bec2f0ef1905d9d4eb9edc9c3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68cd4b004e7ea46de5b11bfcf75c76372f7b1553e3ab09bb560af0f2f04e23ed00ad6e9cfa8e85b95f2db49b9d43efa60824ce63502459da99af8180e900dbde0e3650b86997742c2da24c8a1166312ad508f910e56456e6d23976a62e579426a715;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1278f04cd33b7fbed2a5501dac423c1b76626e6cc3c580f6a3cdf4f317d796a6c3e83e68d8499a8a7bb3fd9a7805e1ddf2d1a3e9ef51933256ea13d9954473d4c2dc1f95a7d2aeef6e728cf0ca09f87c34718367b6ae15eff9c2de6d1d3126b9bccf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80a95b8f41920de6d16f2c58e4e47c2199d193cf3b7db37cb9c74402827f79d031ff5ff566193dc9575de6a144e685425b9840e9d4d6611ab0c9098c17e00ef2a8f74803f0391fd9e09a2f63d7715831c8bb4964917c9358c9323216fc4de70ed1f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha26c5915f8a4a31cca13bb6bd2f94b3b394cc1b3b35ecfd7e27db5478fd132954bf76630220921fe0f810dbecb4a783c781010c0265e24b5d3f54e8ba0a094d386f0a3ef3fc592122498fa7dd71eb409f508099c85134743fb07f7db6ad969b04de6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8be8317ba1279fe7e0b68144c165fd8927b06eaf96d89d94fcf2c579c88b4a33427257e427dd97933a211157d39645f55528f4c083fb931807b78c809624d00462ef60bb9d32fc739b115c5cc85f9e0c1b942c3b1724d96648b7efd1e44d48090bf0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a3e08b2380287f8df530615110a27581293154cd49f79250397382bb5ed004b7a319f27ea173fc066614f0a61f6bccde447f798ba8f76ae8ff5f2f8f0123fc019de519be30c9a31081826c8dfc1722bb6253d6b5d6cf2eb82a6762a84e7dc8e89c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb4739436f5111530f2eb25affa56bcec2504f9a86407703598b05502db45e7911b7295331c138d31f70e5269bb036c8ccbea43f1d846fb28eaae6c5e76fd0c3cf6bdd54cb85ebdeb7650862e522929c0a37214e628a87e38c4c68a638f73da8df57;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a2d211c5af9ddcb8080547c1de3f535f133e31cf4a5d08280958ae9efc49eb99baecd47d5e74b7b88e73ee4ba1b05760750650540d1f6fd8f05cbdf210ede9625ded90dcad4ba063b05d610e19723a3f91c10bf5dc7212f390a3c42cce7f4ae7fed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcebc0c58fe7a3b65753a8adc48e101421e7f6ee5602e0b85396b03db380e811128988f804f05cb019c7c2af8d65f7bac327e20a48b79c7332521eba3bf977c9edffaef0794c37d84a744ee98f1e4cd1c5507098631d7789d0713ed418141768106d5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23fa1416cebc82868b71e10a494cfab96b12d7fb9b5514cfcda9d221ffad722d67000ef23112e8b294a9769934b95982b006aa0b6b371d7ee4916ed00a1a4e4694624ab289060eda46d5ac29b0fe0c66c53637ffae00c765a20d6c7c827060befb32;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e412a76b6637313d235c102872f83796d19f647767afcacb7f980ac9b9eb452b0739b7491c4768f9912c85d1a91eb50a82b260d2343c50c5a674ae6c350e5d62f424a5ae91a876e7c99b7e02ecd9dbb24439326e61c9d87d989ae208049574584ec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98a9826a0ec294b29a984990408c7f8d0c64556a15f4635d217558bd6d51b03556b1028db88b0cb9971429f338a7b4fc6286f696e7f7e025469046034f81d4a11a1b544f17df1b0bc629d69b64d9b1ada196ded22a1afe58f6fbfe75754216681de0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h934e80602402b2fab600741cb0736924c94f9a1808fb2454032c2b19039e32fe1108071e5261143b32c3dffabbd6cee85f9588bb07bb8b3ced9ad02e737f0eb955612944785c252bc3454d0a1768a753aa1444b098617b4614a4947b939bd2a3ca04;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91f06d39b0fe733c328bf26db3f70e9705bbf7de6ed777fbb141e749e6d0cafa1507079a9843dc9c20d84535370876e34167e1156ab51313290adfbb3135b626ed8487a36a948f6e7105f8afd4658f580ea43e11335cd2cb0f937be44340eea2cd17;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56224066e629552f245156b3647b1a623179bf233ea3fd5ab872ac7f7aa76e583c58accdb8cc74ea9a327b3caa709ea563ffa1d6971b567e1bd316e9ad6af5d00b4d7dad9cb6007c87294d5358f8df56540596420c457ca7c8f994a3cffd28466c54;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d9f0935e095cc74e5af9a4ea374be2b71ab4c1115e3e24b5dcecc149e7435f629bbbf9c94c545a521f22b0df37a06ca122c259018eb9738b1cb95b522621917da7ec01fba0c023ce466988003a5da7ab591b42dfe48a3dc7be2fcdb449a77514199;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa783b303bae245f5db736ab0a04fb687d36838bcdb05efccfd263ba873100f0514d6a6d97ad961e46a8630c7f3d1909b08af446bd080e2eff6052d70a9627f72cf49052b87a9c5ea83e3b2376738b4e876655b9efa964bf084155e94dda30ae62aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a397505285895722b85c1f64f664047bbd44bb58140d18ff636db2c349a5cb37e54bc58b467e097372a3af211b56ed86ec48fe71390b956960ca86d67724e046bdbbefa65432b5940950b2298e85dd02d5f7d616a239331077d40cc5f48013b5543;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h539c153cedbca1348926815f5a6b9b352433e7a8f41e2de8cabf1b1762c55d6d9d70ebbdefcbf900353acef9dc12beab5276b3669a3bae0c0cd812fbcfb9091b2845aea888fd76d61c51b852c99e96982658f73c2a08de2d40aa8a3912fe5b8cd38;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32eb8e19569bf24d271d666dceeae872f839938265a6ac8c211328ff1ae5b3694b5bc4067387be2b375ddefef8eb18a4a639a79f1cb98b3ddcb2d6b3776fb51e3c736f5c3ea7017a63e5686be79b33f9e1603d28ef667e9a135888e4ccd60ffec866;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h270bc4c6f7187acdbe38e39cf203f73400916283a7d42e1da96865606c6528a69443dcc025fb87be2649ca2a48e8f3b93a5b58b97e3d3891ed6eeb24b30fa2663486999834ebf99ceefc704fa49cd64651ad4348e89a81306dedcb6646892febfdf1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf9757f9beac9b5fb9cb5b7ec177b9794e4d6a01bdf1e4fe8228d63c1efac0f24134df33f423c18c84fd7bdcdde894556ac548174176abc603d1f5c5a547cb6be7a838d284b0bc1517e06db23e53e5dd8fb510ff06a1124a1d069169914a9319785ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1af9d9ffb4960e127e4db81b189332263e58f274a5c1f5dda3a13db6afe3cd992f96e58157545a025fcf34093919a26e57464112debc283770a839435c550d7e9ac634671a1055148ca783c66da572106ffbf17da608e613a8c929db724f4dc244c4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdcfea7ee86c631c96a3223038297d8926eee0eb78bdc6622b365385484a2539e782a0c3978146726cdbb99b1a7375cc5b8d1563c6b9ff09c59f05099ba16ba10bf65a697e7118f41810f82aa481ee7debfb7eff90f1ffdae1d7c09a9e7a8e121a7f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76488921d088dc173eed058de09819ea6586fa8f30773d1488b6d8436c656da98970e73fdc62b9acb9c2a4b41ad1419dd5d2320c06a6073ba03b74f57d38c0d13d531362b9cd24564be782b6ba846f88a7aca68b72b976529f58d63829c6dbb08194;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddd824e3c210f014eb6f73081949bdbb6c3b21f9d8722095eebf78c06ffe2f51e03e9b4757960848eca2842635effa11a3fc0a6e10b4b26654a04b2bf41be279157c0cc07fc15409a3567d651dbc56d844fe3794cb8f2a58455e87072b16381a542;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e56b1a3968219da8024fbf61e79b4d76088f9a300508817b87a0769db372f30991c22d793af9628d0824bcb0cd13e14231fe05f1d396af0388ab55e7a6f686e649e35ffd786033de7bfb4a49a893b418372bce866ed392813c7378467b293fbf148;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfda02e460b5e9b97a50f00bc59382f29104a7a02b918337c08def414f087d30e0fa3a96dac22373ad40ed07af67d5497e0d135a77e6c2a311ebfbdfd9b529686f5d3086e9c0071bd22dda5dc2155762605912072b2976517b3a308c86e62952bd9ca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71aa8f751a7b9eec0d7c0206bd9a7190e3ceb723a2d76f5acb3fb285e833ea654d5f5774946b6bb5665db81a8935955faf75edb729badc85578810a12f098834e69ad0c15f2ee6b218fd47bc3c966577ad686d03e5e85bd16bb0ee698f96033e989d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbeace9f739cf4de21fec46860f50c862f232023a9481e1362d079b5e59c9538bb1ac668000a49a9fc0f17937d4307d85221936f2086c6449783af6c3c9a2116cf8a256aab88d30ed72a84576af837354f42de251775e017497621d48bd875776c6ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2887adb04a48ac3060e470b0d5886735cf17c6120e80f507a9e0b7d97e581597edb40221676c4de11798cef834ca49048c8b4d489a840b8b8f98b5eaae6134bc171889513d35423d7cee177792e3eb7ea45b4a0369522f4a66396a3c7898d1b7179a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6157d399e7154da003b59e16bd0022164dc0002eb513a25d8a8bb86fe199ab79bd16765f94f8dbf12ede592323db9eb6b66955ce11935380194ed7afa25062ca3af260755b8e8da66b9926bb45f692dcdce312dcdc43afa476d74ffc7ea340a30a7c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22934b267f038b7303cf7f0dc8ebce8e66e658e328ed21712a7b92b75054a9935e3944d0d370c1627361a5394b509b2e75ab237350ea4b9244f2cde3fe03b135e5fec152a3a702102b1bb389806b59d254daafb5f6e08d392cc21e75d0aa18dce8f5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e2751b02d3fae5bf4ef55128189d6e7ce56138f3c07fce9cc75488142e41981f352e28f3ceaf5946c8beb14e6ae6deac444fa2779e111e67feafcdb8c18792f0bdd3c8f4db8798044ecdea0e3f4ac4ca16b28d35b821594bc0ca00835e15d38bd36;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3dc8a3ad7237ecc9eab681dfc2cd327c96495760dfca34138597d34fadbcc30402060bf9b3e36a8ef628d09f221c2e122ea1b82f82cc70eb3228d1a9bc0317e51c013e7fb103c2fd85bcbc40426081844a94dd17d431bf118522534d908ffe8a6ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26a5dc93f210da86071204a49fa147f43db9c54cd9b56113f558d7905dc374482715a7bc5f7fe09e2396eb87eabb5e2c3a41f10bfafa521abc7767a87be2e45485f826df06c80856af775c64c32244aa2e4114ef016e4c5a8660bb781a02eac738e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf964d9e95b1a083dfe53a2d15ce4f8b6af40ce1c3c5b759d6b51ee500b830aaecefcd345647bae2237bed2d7718f833212ac39b27d8f9b45b2fcf84bb1ba6b05d7855ab6b4f011056443d7ee462f55d814105bd0a964489edb87fac00a65f4c2855b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h535446373cd7b7c55117d6bd8da66b57a2409a334b4df476e36de05a4563ec9b84ed738b7f5f98c02432b37a9886d02b625b9c83933f13e600856529be2f33a1bc317d565c322770c1356abc8a0bf580ef7b3063af016c43151655d533c40dfefcac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67a45bee858ad7a22839f01ba7bf01a4e04caf0a57cb1df0fb4bbc51a1315f0f4b77ccc653404c433e6f7ac3c08f5db9c8fa746f8149cfb83cd34fe6c649796a26288e115035bafd8fc687db760269ccc602a35937ea2a068abf99d34418c0e4d49f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1fc17dda9091b1d5e9d69712ed476f0f1c119ae4fc0b360130a0147312ad16ec9aa5038805ef751e20b0484447b2dd88a0397ea2ccb72adeeae0ef2d007c93f68a57cbfb8bae9b456f88740a164d036375a25d5bc64b6d02e0e6a985c8ea30861f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf11a483e3ad6e3ce2967addd843e7a05336b14cce55f859b7faf44f293cc9da2699c86e3d18d73ec092a08ec28a37867f761a14e531255e57735651df05f3f17edd1fdd4baac57e1483c138d67f40c1e912aef24567c5e64a0f69c0fd671d8076230;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81ea7429b857a7cc4a37f152c41875d545316f79b4ac93f60df0a7eae1d01eb15da73c89c7df7e35933285e0e558334fcb4bccb1d9a3a6b823c18b1da08bdf6e2cd8110c11e15b14fd4ce54819acc19a1a7d4af00bfe53cee65b5e289685b6d609ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h307959d171518f7adaf7f6cc89ce4d500b5486088001be0bf39c2d7edc176ab8c9ed9d29b8cfb759dd3edce5420b326e7ef144d27b436bed019d4ee2d9fca44f1019bedbae5315f05231e7e9d63086d3056ee5fc6c8fa6eefb1501150a858582a9d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf695cefb0041acafd86dadb8ac47d62b8f36fe1307e16928471a9839e94fb0b622aa439e0536a169c959b0641043e76b0194f05ffaf7d6600d28e476264de90e1b531f6e65164864d23fd849451de949bbbccc320da4bd156b5d4e2d2214c3f18712;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34124a8369e81e33e4857e54438650edecaf10a4b041cb8d7902b5a0ef569ae9aeb8de52fa2b9be2330f7a80afa9f044a174c3800f40a32fdd28e12fd751da872fcce09192006e83a05a6166f76a815c11c8991b2ed62de2188417a9c360c8c4f0c9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca5e3a9cec8d23fcfab07a292d63fd86961e72e09d9bfaa6d92d466bf52d70c95b6a4a2d32cf6a565396e0b6a066ad1710fd2ea75a8dca2dcbe0dc57d02b86f3c79db4f19802f4406959d3eb285cf57aa4871c1ae567cf7cfbbab0fd6849dfae6bcb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f27d1e15e9cebb2223baae130f32c033f23c4f5605c8ca4ff89123ad2ffc9a1bf90158293480beb7e86b4faaf8f1e02897e9f607b9d913bd3e6365b224480afa4f53e53a8771ce0f94ab32105caddb3ddbc6b74fcb7f98f7303d373ac4a12249a06;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8372377e5ce988c8756a2c23aa2c07e8e2e655a375975f85c315754075591e532394fd608bbd6751376f765b2d04f5d9ea7a0f2e80d272f501c1472f3abf0a0d693fd37299d5e5ac5f07cb831e86b31584466e0d1175eaba360e004826e408653ba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h807ed8ad23652d1a316498c97ea2da9f22937f035a5a5af394646a8ebd4c5355704009b58e4477ffe0dbcda3f2acd41aecc8e04515c1507b33330bdcb3968d8adf788bb799ab43f9effba544ffe987f2fbcd6c594bf36da6c932cde3d1e96ad4a38f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31f5ffd99c536bbe1c41e726a066664564e7337d2a15bc33724c5a41487cac05f7445fc018287d556a6b3591a9a66da0901e427d931d99389eb4f29f1dd2fcb109e09bfb1a4be882d9ac06c90155567d94930d579b12574a1b730e1443443dc2706b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d135e2fedf163b2b0b27afa1c39e58e0200510be7bf9c3aee9b9a399fb5db411e90b7a41832ff0ab9eb5dc3c49353f5d744a7b005c59fa4b531e1df9735f0ee5f17bf8285655657efc5f98188dcfeab305e20418b864c740600b39e5f06809d4bb7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2596d3a4d5960128769ac8bf58568673f67004ed404a30a880df671b72fa829bf5c2d059cd66da18f03f82776de83e7e786b1fe0e4296f595febdd18b470f8ba8b4bc7de26db185f7334825559194670e9aedc7a6d204bee06c745ddcb2137ff701;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52a1bb2c2606e24487a16b181c55f8eb9573f0d256b39114e66a9f82a0d50a62179556fb9a9812b8268d441cf773046cdd0faa17b4d51d2c7acdbe9f95074d0369d8b4fad5e41cca6a3b5e353d29d4e9e7d0c70e34fb098b08f4bbf69ca426cf6cea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he59b63872339ed062bbc3594f17d6fbb8733b11215d6d9afe62ee28427788a386976b509676d5e0b50dc837df89651946cebcd26316c59c1d44046c2f0b7e73f0e70e80b4ec7b998736f4424c5b572bb48e9f5352fa0f95fe7a16999ca6c150dcf26;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2715213f414c7fbf914c3f6797baf05a79de4139d0f71533cdf0342b56669888adb2b2629cab01f0588b474ad40551e1aaff105ee530b9e34a6e76e8c3c43a7a3cc66a641433b6e644bb5f0dd4ce4069e59d6b38545ad2b953e66259d700374f087a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h318b7f1ab0c4dc027fdb80bb04a092448e75d8ea873909f4f2ca7667310b4423597cb36a11ab50293841ee08a61ce0d84895a7056cc694eaf8f2213d919ffb63738c61394a286af8c1997f4d8aca682a66753e021b84cafa64f083a047bcdd33c49a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef2e6e333ce1b0223fca4f66657715d14582b8a7f17c10d05512a0e44dff464cfc95af5c6baea8befc8833397e4494b4ab687df633e2ad00a00d29708929fc36fb6adf08e3d8082de6b1f2ef92cd1feb721b1cc0cfbef5246d17783dff88be83ed42;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h312854eb1e0b62e24237f4f391eb4cb2d12bf341cd32dc23893ea846befcfd213b77eee6e9e1d3d9badfde1ce3c1bb71eb723aac51a1feb0441ab2a17e47d1b89e207a61e6cece33302cdc7596d825dd1f3635191d681edbd4129e4d8c769c4283d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haba37808281027f91c5247408c8baf09e4d884e3a47efba7c22fc0e8e625e08c0e2aa9c28d682cb83a815213ed2da81761158169aa471cdd373f011b143f551d03b9c16e3b7b80aaacf08117249bd19f9270d4406e5f469d94d516b5757d1737a148;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cf928e1479e2af0206f4c0686dc629c2923210094998266ca5b0a1fa663aa4f4d85fe214ce0322841b48e94382f2f9c2049af936c2852830da681bbad07b6d4be312a37b7a8db7616112ecb167241e1fae6b1f07982dca4b9c6ef1ed6bdc73fee2c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48f989beeee94c88ed23f25c045d1bfe128b1fbfb83c260297b37b64554ee3257947b580cd4cef041cf95ecb9fe4ebf33d1b80ea07ad9053a18c974d88bded455c9eff5e44aec658af11078e3a99e34a58304ab78fdfd58faa84e3649e2330bc5379;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50837285af9733922c93dcfd5d1b6a2c2ae4d7b2447f68e1d556d1981a1376c4c496af86bc48e8d028d464edb26885a64b33d1fae905fda56f5a4db276abfb541f248d9b968f8e8ef01827a54487b8b233e9030e20cb27fb6e39efce1932122bbea6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1dec1112190a2478f38422f248df07d64df5d33a4d0ac1da6a4ce56e4e6def8645a01fb453b9a28ebef6ec75e5d56520080272097806992361ab4af947e8a623d9b93131e4362ef95c50e9d5e0764eeed3d138df8bc2cbff1479277f9f63964bb14d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55bfb257b57585e77f00de6bdcb7a79a7c7f51c3efba5375abbae48bc1e3d854d9851589f6d3f00e38f4735167b8e51a65af7738a4cc52d852210907441adffbb2dfb14aa90ba68d3c9a5c8693d7a1dca1246af231fdd2cf0baee6c4aadc0d4cb5ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79402c53f1fb1d2b649458245fe80b98ec07b6725d7665395718cf78eb0e73a204bc53b2c4e69829a98996dfc081d3a73265e2a21200372806d2c4e5e1ea687408537e68633a70db1a9acc17331174d483d37fcac0eaa68c6787a085abc5e71bd4ee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha91a6c92900ed11938fba954505ffb61f71228a4dc9604fda5530e8f3e7f1ed0fa12e7ca749fd3b14da6f8e3f5bbdba9a6730169be61e6bb6815e6f0bcfbb8cdb641f3dabc4caae354f4c7a57ef9fdbb3532afe24393351a980f03b842901a19316;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5dbfdd4fe570f8cab2d75f9d2d2573786b2f8ce16601886ed228c3ec5a641956b669a0d18ebf4d83038ae435e9badd318940986d25a5be94678505e1d7023c6b313952ff3013b9f8e7207f2a1818d90f1c4050c70f47185d771087af57560d29fb7f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h932290d16fd78024b6da0be6578fca4eaa171cd85d1b01cab5d0a467c34b30d5186283068e8696a577601b7458e7718cb77de906907593f70908b00bd9119134501c6f384ce110a9150f39724110c96ee9a3f832290727e6df3da53cdda81d076bf8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9eaad3cce3fd54b282e63925483299a4d07b9a3c436e790bfdf8bb40e06ef4281f058966bff2e8751c54eba342104ea536d9249a10fce44abf41802ddbfed44256180158e6af158b4bb24027fb71bf3202de08e75e3ed1919742d289da5f0680c52e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb66116eb6b0f2e39b9c403a7f6dd1f499fd2e313c78eac754a113bd928fa73169acb1c68788956ecdda7770f5b19a157c8a7fe1aef634762b92107c4db8982a6deb7b917dc5fcb8c27eebffa877fa0702488064c15bbcb6e187142b2090be7d2846;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h893c161438b2c9c3119af2295c009660d3e90ae530bc382f2869fea89fc340f3a9372a1cb333a5874d3d047ca1b0572ac43d8a6fa81d29875a67bd18624281f62fab7e8f1f0572027f4c6da63e44dd3b11b0c985641604850a101490d50f14b96722;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h642466b42230cf6f54fc4ef511477700b2b3c52fa278f3b34ea3a357d03e9d7c546ceff88b42365da7955d946dcde51a2efaf76b3a0b99e4172040f8b7d0d64d5a01c5efb99e654b043ff079b3ddfa3201081f31e5052c6cfbdf3062f8b1c85271dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h955f689e5b9618d1e93c71faaf706e89e41cbdc2df0f319719160ca1d1dde562847a8320408f9dd5d78bb8a35e82acb7b807754eaebd9fb5f37aedbf6216f0421af9fc41341f233b1e408c9a7b4ed4c2e0f33ef9b2803ad37f5caac9065cb6485e5e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43385ad5fbbe3eeca0cc396f65d190b06800d14bb2068f2f6ef1e5f83e9171876a674ac3e855a0d6826956750e4ac9bf8ba4ac2aca5b2b1b82a1ba4007a1b6629c96b166a7903ca1b1c946cde5df104eee36991aaac23d068518fb72b131c5f86d8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77f97d5c468a6e00fd7a084deba962019083ff9add91dba12a218d6cbe5b771b60df257cbc6111b97a32df542b8098d72551352772fcb35e583343f2b8601a971fc6d45e4a905cfb720bec93ccf19b0685a018974924fbefc41d1c870f604ded1bd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21d7722588e266e5a9f298a58e823e5ceb72a6c979a2f9d33e374233b0ff02319075c04715ec5347de4b4b1b9e7b84b9276468d07c059134d71a37c826a51adf934c2ceed2d2f6753704e3e0c6a1b491ca0b2e8272b8e637a2d94467682a683b5220;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7e9ebec0260321d1dcf57c0873730cc4a3017c452d9f37bb66ea82c5cdaddacb158941a1f946ee07d7dc2af8a0920a17f0f9729647dfb4f8e5ecd6e3877ba4c381396dbb5c39e7ba2f13aa3eb90b03b7c86b5d6489a6f3ac473a1707b9a4904792e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8a2017955c9df0177d6ee749a77daabed14a942de8efd04e76717e51965fbc51b438905c287f4af306a70c620e90e55840e47b38f6b8a1f0ef41aa3c8a806a3e7f239042b6846590dbb4af014fef6a35ce764ab6307dd66fbff4c7de7107d6242c5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf30421692d1e98332a00bb383a06a4702d49f01647091b2301938df143ce0889953ebe86d22ae67e66d60b6fd9b09a7ca04077ba2ec533bf5d09d7a203b3663e9bc4092b73c2842e3926e070463bc70fea7dcf479a353aeedecd1f7751e3cf9341a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce9e7b055e7b1629dfdb77de49c7604c7fa3c80743ac6f658523b92ba9e0ac1bb3d3f1511b2dfcf0cf4cf4fabb2288892323c312674c06b7cb5c8e698fa4fb381d060f67fb2f03190713e872f7788cd5f646a05079ee076e031a73db94dc8caa50eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40d2581239224a7ec2c7d1c92df5ab975c4d9a64d5df43b4bf7306e99a7c953b14fb364fe5b0d9476b42608e8fb601141a5a1631b5063eb5a02a10657b478a2f1428b6c056bf1c92b4af4728997898216f1e5dadd86b9a26dd8d27d61491ddd87ff8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h220633183052286a58aa622693ff25d21671141e6ed355f0484cb227f0fae75aad1adf031b010de0b718c175b0663ee7608bd1c24fb36525ae9862360158d3a328def92bc51d28ab55b384e4458d500d237df8cc030fea2dc769000acc21f59175a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8cda321204440481fadbbe49066c65c46585ff6d02211a85d0b4c457b7f3175a3b7d15a483dfb0596a0232386d6c477c0db922b45a8cd30ccceaba7af7d52022d6d5c7722ef68754ff18f009afd9287d0830a6310a30da4b1a78b1f804e9633fde47;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfb4ee62c60ac6b378a8be83b959029dd5255390cfd42ebb3f6c776ee995e73b0bd2be2ea5a68c30d47cf09e7b5cbee9fa8b7821f0bf246014d73890720ea9b4565b49b0d5a04f4321c09010fabd9bb1c87e9886d7c7ab51f47a8f1fce90cad8243c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c61f08ddbf9d47bad88cfe62cadb513965b198fb18903c0f4e6144fb6596d8d4bab52dcb3da365372607226b75f2bbf9e3cbb2a6058017c28bb6d74c69163c9518eb7de8739b95fa829955273005a296bd6beb8de9e02cdf1f20c764d15c3d0fd70;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94a044a1243438e4ff499fd2dcbb35b4e4ec4d337d0462aba164b442ada525f76af4505ce95cbd66588594489ebf427d9da8b25ab8c20e5b2c98a8ba4a8092e5b242c657f6636e2eb47dd18d0f602b0a0bb5b5e7c9e07416e9dd7fc54a637da01822;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b092a7dae51ebe25f39c0fedfcfa6646119982609ca32f67828a53ce7775d8bfb230d910b3f53fc2a108edf1920a79a0c0014a6ab4d7c7f1193f325010fa86bf5f91c3d143bd83f4548b21089f9091b2dd12a18b5fc9fad0ec2219529c462cef28d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78c9c6fcd13458d36612508a1e01ca9f11ab52d536c3525ddadb3d21e04561aa2d67941accea0db1ae7eb7ecc1d8253cc8fa0c1e358791c4da0b402b3e8404d3cd4c4ada64aee5730048cf56c91bdc7fa0a4bbe2a9d6aa3d76656155fe41653e7567;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96915cdd7f58801f02fe86dd79b1038e5def11a7b9547d72a340ebe4768ae76e7093ce5c679153f824133bc5946d05f68729a563f4db9c259b7d0da13334bc365acf282c3d01b25886bedffeaedd4326614941db59a1b1f77eefe6c6cb0c0d076635;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79acb05d6d1e6f26ce1f1090cecce9d172bdfa79e5dc8eacfe337d96f93411fcd43b3d2b0f89e8e5e4913d8848dfa290a273ca10f367d4e6b8e54b27a69b5974e1298ed87701ec5dee304bbe6af84bf30a9086472dd90b2718d5204ec4ad323843fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84430975b1d76969cc99f3ac11af35354bb1ad88abdbc52ba89c5ecbe99ab3b06464314a3881a56f1eef42a060ce49977d45efef837eb967e1ce9e7931c9f2586e93cf24a55b714dd16a04d6f00841dbf6d720056bec83b3aebd9d26bf3a25b89fd8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7201fba24ab364e1a982cf04dc9d9669d3c4b011ce3e307b71bd2a992cfb451f2d657c5c6bf96281e53571730a1f3cafd1f0389332e3692b262b006d6191a20666006e60d62fbc4d83a72af1941c49c5bd36cf4818e546541b1a27967a601a3af47b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a788b442fe28be7b3c02407c92c509aa6532d235dd2adceee08dcf735371bca958a52d8a4702bdcc2b683990cac4612b202f9152e9c9d987d6e785c6cf8a8c114b9570032aacfd4a9ca8d9916c94d4ab45962f12c8e61e2110ab1387bf1c0de3237;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc03b5bcd0a5ca56e394aaf9f393151945f85a2f1bf238b2197c3df8ca3b631c09c7d17a3a24fa8a5de166534eed7bbc6009cb36b7dd6a9b7d2af79235fb8017c14d9d8d0dc135e05f740fee74a43e12577f02a4a76888be22e0ac05f95c7c230304;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cfea0e5f2de47672da0447f2bf09cbd5c4b87931c6f3df3d921d27134c08fa1ade95cd95f11384b45b6f4b6fcd1c70a44ba5f3dba058609c02ddc702ce904b365f37c4e1cf350414141cc586f47785f02fe84ed5ad44b6d0dd2645a99ed04425b51;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e81e17805890d9ee7803772781d5ac7e9d36dda601c0c6ce877063ac6de1178fb5712360b2b06ff51a55138ba713f1c339e84b3a5943cc9fed8bbd450cc408e68198c57a0419f162689e446b14ed4fdae4ef91b02d3a7c78a5aae7ccefcd09f033b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5302519f5e72d095311a07d567cf7c7fa2a313219407fa62878a301476f09f72c52d5a9b4fe2f1c1b9dd92d9ee98ea79434c641c2a7288c55bb1f46bbbfdbbaa5e99bc0bc226d1c4f6b861eba38b8faf014f9f973e269f39e27d7cc46694b5c84c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77cb957f8efeaa5f9287668cf7fbcc28ef4daf02035205b970818c9eb7ae44e398ee736bd1938837a6a973fc6697a2a9c40e3d11b57b0a3d1baee8a99bcb38555779f27d7104479da16c0521ea369f224d2d01dbdfd4d9b5d0d4532264bc470c8fdd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ead3f633da8d58132ecee542bcb93577dbb63ace155b7c093beb37c9f7fd10924deb1305868170643cefe284f4a83d2d23e7447b2a777141fa2ec6e6c80192f96b7d348af7a036b4fc345eac0ac031d0d60613704a0ef7d60ad1de1ef78edfbe51e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h281df369e98fcc801b5e8022b84fa7dc9b703bee237600675e9e9e69364fde5e8a15d60562bbe0d1e3c375b3bd50952883a5357b9d33b138650bd966dbb0dbd5001936b6e73b3680eb759083b58a405bd6952aa513fcf426351cd68e6b8cefc050cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h483f7e89351fba711c1ee937ede185e2cf231ce4b5b25bd87742e409623220a82a353c1644f7b97df071ab30582cbcc1ab255924de2dda3aee5feea30b4b156acc80fb7c92519393068b4fcd63f98213528281fc1721b957b283336d83146df24c52;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b1a9c6787f08643895bd421efa14bc59c677f5dbd40c38d8087ce07013c6781ee4a9d510b98c11885c9a173d81e619ce0ecca7cdd4d3215a98ca56d1f15e4214ce6cf4c66c25b6ef49dcc209938b4916c31e342328ce372e217645d0b34f0b07356;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1b746798a984ca3216a1fd0abbd2dd5120cc243cdd4a1df4d6f9061e990365ea4a63cfa5088175db60e229f2070938e8da12e47964c3b74b70360b45ffd8378d6f9177f208bc1d7e61d35a0fa7448e4c9f7fb0a58868db69b22735aab107df07f1c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c1664bfaab9fab5e1e9d5397e013798a33496911505d8ba0a6d0b7cb8e8d56fce7105f49630e2cf5291c6c24e0e6a7fb86565974b23edcfe7af007f8f17b970d416b19e406ca89ab2d3171035401ded86cdde78ba0e536b3b0fa6953adb276d7cf2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35c906c993ff1f8f77fb6a03be467b874bb72dcaef8478254d4aa4cb9211a89e490f2c3c70f1b55ae5031961f29f3bfce4ae624158b38793845113e5f12a4cd1ef36f9aec0018afce95185acc498ad3c2cc20e3877cab7bf17fec2731a6c5cc0390a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17ab2cec6f5b387e7ed779d7ed54e35c550f5da98a7d0128f1edfe7b9ad42380e491524a2fa70708e0005c34916d8a6e0f6dfc19af2a78cdeee79548068e61a4c98ec8b6e4febc5f547dedbee0faeec87eb21268fd33d298b132bc93fdd0e9169cce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ff2b99c798d55f8d7b90f830558dbe07faa56a749cd008ea97543d1ecdd5356fe3f960db989dfb95361063409309892a44cf8f1c622c96acd515aa50f5b38afe169e19cc54a49ae85f7546c6cf1936ce20484bece55fcce2e50c1de4808ac4a8a99;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ce58eb85f8708e574722a3a4621ed7d63412c3467459846b6b2626bd2636162779730e06e32c94f2578ef134c2a88f503bb738503f46df0e399ce12817cc1e1a413b134ee703f2c7b6d6525fab1d744a1119a3154b29762805b7e327cb187480155;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd49fc6ab95f7d6cf85b2f5dacf14bb14de3990aaa9c5847c816c538119071c35c559525fc857a4ede7be9563b2d788571503f872742000e255c7d9e9da2ab9d59afbe4421208095aa330282ab5dbb1925aaa37d6490a0ef4b31e8be25fb9387b11f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85f3ded40fe606146519740de30036327681f91b2cda96a8f4c70e3031af4b04de8d736ffd190b8f374b1b184b84e7a1c0196bd1420bb1c7c9d4238413ecc15e66fdfffa12c9207c7a448ee1c4c45f79b5a7d654a949199eff323fc5c75fb5d190b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f4d8e7480e3d90de54ae0be6e4a046ee396b8b774ec3f029ba4ed339deca8b9dc7ee9a8c16cb406721fc909c1ad910111ed0ebcacf738584e3a4d590f436139b5413e2652904556422674110e48934b15ce4a3f6b7e664854892bf8857e29c1e03;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha50514ac81d93c35392bf3c81ded4b0e3ba14ce68e5fdbe2cf93ce45dd579e866d50529e5798ef6bfbda85606734763d03fde1355e8c89bc514efd025506a338f109029463ecdfa8660ed64be522a7e5f1c42b13043558908e20b7d5a69b977f5c97;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4021a92a70157d7f28b349fb8c3634041d9f094d45ad4cfa718a4ff9e113203b642e8fcad9d1c4d79354ab0e995a699658f29307b71077faa35f061b2561b42d20d489ba9207569c40465ac15312a34c33c6e178f6aa3c3c7a078da3efd21f7b1b6f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7113088e408c02fb191faedd5a868b6724f27a5de839c6594b6ca6758a392c6d5dfbc493f138fb7fff8ae625eea483c3c9fd4d3d5135d07dd5899b9bc993289186d4490c564136ceaf081369ec0a682538055ce8dd64f86d8ff2db0c73af94ad5f0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8852c9ca9596075517fa8cb7236b66bc19d7fef475017b2ff68bd35e877cbeee0e9f53ce61467f0552d67485a1c890c4d7a4d889b8a4c3e6f082014482287405c05899e471de90f8235b02468878542d8e35562e9d1ca13cc679436b890e322a3873;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90d705c154266a39f08c4586f8a217ab8e4bee80acccb10ab2210989ac01c543ad4564c5f16034cba8879b7665b8379f8cd892b6fac6347b1d80052ff7425c8ffc1d559eb41a6cdc85a54e03bff135044099de00cea851355bad8587ea6641e52dc3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d1cec3ff9f2650283753ecdb0c2aee1fc3f9e2bbd57b39b35d3b43b7438f1fcbbc703396699519adbcbfdd193e79afb141e7c277b9f034659be5406295aeef805e8e93ea9faa1a9cbd4dd21856e60a06e80e50bf59d50a10a4de8f0ced557dfcc42;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3730b997003afd9432150e542b8614fabef51b24fd2328d96cfdf5e286326572f45adc2015160cd267dcfefe7a0b425c0fa67883dfe7afd68108b9b53b3bfc071c402aafd0c87f0954d17c49f81ef27b12b5876f104e16a159c3973edc388aec8a67;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f97c1ab649ffd5523cb52c721e5d9deea2fff2f2890c8c4840a9628f21a7db377e99b93fff471128f56c38be755f8089e41b740082a45017e5f499a1c8165cbf01ccf0bc56c8a58b7c125399074ab4e8d02d19cf6a2d49266579cb67ed1b13fb414;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cbb8495090ef610b3d2c46ab400b100930ec844243522cf6b5564dd87b58f95eb88ad45ebdbd39c1362996ff7a9537950bde182574b9f05c8e67673eb0dae7ae29946c8132e2b00b80034f1c1939ddd869f894594178cc41e731ea600efa0594fa7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha92732fedfe3b060faa47b08042dfe26b12bd892d1ec14c62c3bd37dc4576fe33af6d0a5e7f9cea217e3301729e53e9c70cbef3f69edc72058f23336b53a38e765055009500216a1436db8deeca6bdd891749cdec430947c443c6c01aba001f97164;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3312899571473934c3b0847db12321a51d04ecc66bdaabbab1c256cc4458aadb9f108b07ec7d46d6e706abe3aa1d91ed9335784fc6ec8f44cdfd262dc6fae79199d8474de7c1f225daa0550c64e8b53d73ec49203ea515ef507d362c90a5925fef80;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5191ae37fd1ff46ad2a413bae62b58540c2d2ee8f82db3a36d5fc1b6628ba7026d4e3ac0775028fbc5618cae2f7a169c1cf4b3077ed3fedc1b1039ee958728e4e76bb5cbcd180d04c387e0bf6de3adfae15cfa6e4cd3fa07b449657bb288d057f8ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f13ae8d5c03008674be41a701e8403e44e7f0f29835bc4af999989af277815a800cc05540843fe32b3f74c5339f596449690c3cd4b3765292c3f00ffb920188f52c491e7ba10002ee77bd5bc735c38c9ef382deefbf6976692588882442196f9d1d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9436ca992e57d9012376be9722af03dd358b03fbc0f1c8b921eab320ecc7cff7f87735181e51acb4bd8f1b4a8080cc1fafdbb06bc6bbd0da3d1c5549adc38dbb7a7722b4db6b1370ad8a9700a035487b5bbbb67768e33b4bfc2f31d29c6feaa9731;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86b004f0d3cb1544958296c0da97c8c8f9ceeb2a15661f0bde4aee6e3634f27a048fbe653f068d8c375619a7d4d332f38cf61c3da3744bd15d43600ec1abe2d62960af3a62ec603ea06be5246f73d40a269133097633dcdffbae71f503a66e09eaf3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d04f655f981035d48301ee93d79272c686126735c438c4bb566714e0016057c392ca4b872e99f8aeb665561c185f772e44b40dc0c8b78979de091cdd1edd1c5726dab06c2491c676eef649ff19733debda28a83c04c018667bd7cffc280585d300d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h931348c48431bd893a88137b6877b5488c665ecda38701bcc1e06c4701500dd970d5615e7f95aeb32e222fab8469b65e5141fb7668a3e28b2180cc004aa69bd1ed76e06a7c27a9114732e5dab62f5caa8b1d85d62af0968bf0eaf5da14e27d64b4e0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5920a071a3dbdc3193a17de141cbb95e4abf23ce2feffa9e12887b965444abf3618612925a41ceb905f9c5d091b50fdf4dc9c4b7f0f94415f9c33cf0177d219cee6f6141cfb2210a2ff9f7c7a5aed63f6408651edf34e411bde3e6c68cd7c081c174;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cdff099f56ce075ceeda5b0a0740bcb6096277a53fcc856e2c3ad335632c59ef0f8e69408408f4658facbf7cd6dbce09fe841e3a283e49367308e90fa527726ecd033f741c0f06dfd6098d1fafd8c806d4b22e94a638f3cf1ed08fe87f7953da246;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89266c3e500f7133d91f0d72ce1f941d256c66713326ac0c90f1fbb2a8f4daf291bc208b00c4a434677b47a0cdac9e5261a60069c5a0998f28d8d65a88bf137860134f47e8a9e71c67b3f33348da1fb2b5c6912843fbffb9c161472a2b975c5225aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d52cd80f14e9df12540f967c969e010218112adfd6eafcb1ea40c605daaa60993ea9972ffa42c30e598a5812153295683e4d9178c017a6aee17bf96764e8a0b034a110033db56da904a813617508f448544d37d8eaf07254d4f15d57de857ea51f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4a27616ab8378ebd154b6a52ea7c4fe8e368a3e222d6a80132f4e825e4614ad7778f82c6b093fab13773d9624da7eee0b90cd18ecfb5f3269e6deb61dedf1de834ea2636c3b0ab433ad130d08d829d2e0577db763ad37d874aec955195bdc4f7337;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2eecf178ed4d04af62b9aa982133adc2b1b9a4e02a5a66a3619096a11b589a6aba919c657bef04615b98e4b065a292de6cbfe7e8447945e3919878908d060734dfd512ae246a76636695ca1ed30dea55d94a43ea6099cfe12717129cbd09ff295f8f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3768ecf4c1cc797c9175fa3307d1d83045ef58831074dd90ce4310a9e6fd70ef7207d6be310c0266de2a4f754a4c10a85087c34c36bcd559c338426f490dc52c38e53ac0be2acc9218d2e881f364c0b03cc8661d75dcf0481258008c373c080d8be5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd4f5ef9a54b7cf2bc4000368caef99b50f4ef84f7da6d4d09045724dc109dd917b39c74cb674882ffecd813dceed1f78bcb94bf64fc517814c0162ae0a075d8fb2bad0599b7460001f5750e1cb6cbe04e6e0a58dbfed0c59ca4e7c716832b8790b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1322b931f9bd105c35a117ebce51271e5cc2933ea2805cae96943087e13bedd5a4dc2c217230e5e6cc18406d1fff9fa78b82b3bd9dbdd5700eff2abf00686f853b839e03c86e255f666347655ca82614f91747dc5bbf7e295fec005ec457f6ca3d27;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed824ebcb96469b1cac68c16b5ee8158d3cb10d64df247c4eb397b0b63a2c6438269083fd191a2086d16820c8bce6dfbe3d2b4aa65e3fe66dbd78c5a6069b23dd70c81116a7cfca7a411594670f78b46399b3da2aacf04369dde31d91ce8ecd1ed5a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd075b7d233f984830b4b14219a74e73196574a5d53a9fe17069cacb2c321e65414112a2b80babd2c04eb4a02f7f9a1e7026aa4c4ca181a47dce132716d15623f7e201edc4202e8ab29c3ae813c227b910dbf5051622fed1a312cf5ab01d699c04796;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46363328702cec960dcc2e0b4db84c06984f0ae4b54f7c96f3724f01df63a986734cd66c7e0af07bf4ef73456d2f70e614628d1bdceb3157a85d890c26454242d9afe729e50a735b88baae95a2607776a59d83613228420db8e1d4b84349b788f7a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ca77dbc2614719dc1837e99b88db840b9c88f08cda755f1930e43ac94e51f69699786140c9e755a8c36b949a7f7053dd7586caf83e2037e8b5bd78b675dfc332fb670e39d85bf36a56b0d30faee84a15fea3d738d7970e1475f81dd1eb46c5f42e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86d20d2f9355b0578af16f118ce912e03e54d5e3705581bf49f776744dbe740018aecf68e7024b14d95fe7481149ca097dd6330e4f42f3a620dffe70cf62df357924f78f7d32a04e262e342b4019a986e555cbbf7171e3ed77165c7313fca1677a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe02aabe3a35ed5ce4c762a9f0d0791987a109a80ad820ccc5d97183e713a4a29f643af2275336a31eea9dd954f6c6929424107d85c52137435df816c70b54fb120497c63622ab40bf9c1e189c9b34f62fe1337a4b15fef62870ba95ea6b5a47df0f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd84a09fbef38d4e99aa7d123f97afc9177f6d4c953f03266b8af45a0ec229e242bbf30a2c1261876fc83f711883987391f0e6d2e049efd8047199977f9837efd16a1c9f7ff889b181478008a1a8d6b681bc30c3f789e398952fd78e8a9d2a76d0303;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf0095ccbe9b2e4427db29cc63f9a910e8bbac05399cacc2fc4d983e99cae5003f5151d8835d317a13c0aec2a0fbb6d2053d6b920b625f9633c96e3932aa7802bcb2735f9bc8a71b664da74612d7a94855e48d79877b2124fea5f51d8c139e78c2f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8663d90982cb63e2376c734ca79590312bcb0b7688f9d5ade339832c705b774a6ef253cffe94c96aa9bc5c79cd5bef176b78b5e810523bbe5a22716344884b70a12013c3cf9b8ee6aa000f8217d036cf794f29d4e445eb486a4d48910677bacc4374;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h449cb2ca9fd713546043102f2999fed21f09d608414e9a70ddd7fff069d7af7450fef3ac1a644c0812a72b02b6714fc2b73e4e92524f079b592432f0efd9fd50d4d92d8d0b0cbfba90d26d4902e0701ff22b71d8b14514759e283c63cfb67c083545;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h845bf4df8b5a2b0e84777d7fa4f338d95a3888bf103c3b844c3e172bd51da90e3604c0840d5eab528861a16cdbe8c45f84b122b6a249992e4d5754db2bd62a5be732ad4da71fd8939ddf23d59db0ece821d80ee40976d94a1db56cc0d743e5095c18;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf971c5f8510c2bb7b403804b9ba8344de3236583852fb2f5cb8642a106bc75e6ab92fe0be9919da421bd644d81e4bb5c66a47cd71731d0d5f4d75e6d8d8c09e536796ad4e7bd10ff48629b52ff862f4680ed59148f313cf9b97171e842c7e1490795;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacd6a94a4f09b274577e272c9406b2f5357edb088c7f2965402bc946c7090ee301eafdebdfc1a6b7b5e6810a23c69f2c2262b74d29b84e4f7e0db1b5f84c988de5a51a1539e75286af2f4efbd2fcb674a0b6a34fa133896e20a7077fc7a3bf10a1af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82ef506173e6e19b0f9cd5c9f04f2d3414aa146f7d45561ea4f8d73d26f57f2a4edc27327f6f8579bb7203572e8bfeed5373f5b600b35d147f4d67db1af7bb074e384a420efbac3fcec2fd7b67a1d8de1ea3c34b71e61332aab36f88d5d2ba60b44a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4875a814ef0fbdf23ec57aa81b9b9df5868c3f11d402cc5e156a090d2c28a29f92ebe77583107a1f839ffeac7f650d5cd3a7ab5cc7fc7f65c3ee3bf7cccf8ca2af5db254a093a20e06e1356105d57710aab48b3e40fdf5beab52d6889257db095b64;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57b2148e8f7a37acbbc4ad8b21d8ccad1040996a28c813490b3a5554ea8efff1ea3b45f73b16a5acd05a556e9c1c9fec227fd52bd2058a4e4fc52c54bd6ddd0047feeebc4292668e6f1b5d50b07aa036df9b35ec6bf4dba003c1d346052f911ba1b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9754fbe41fdffe9637e6d8b753e688ca1b881b1c2d2708bef4bee9a1c4a2ce17fe6dab6233562aa408fc834d65e0a54c309028a949fd28abd9a30eb64ac8486d6a87223539918860b370c18c217768e7629918db7045b98f35cae8e47da028b8757d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ffbb95e9e6a6a43dedc78576ad3fa7ece25fea2430a5e04dafc04e7db0ef9e227318f25c2a2758554bf7ce3529782f54917f2ae14857297d18b46fded76dd031e8ffb96387e8639c357473f219cb771ea20923b196fb7dddd0ad474bce00fac3a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b7dcbb6c4099998fee8ff690f76aa4a67a9e99593bfa591eb4ef74de7d97761a60d69e27e01a9b54bf4d8769b7ac412fac40825b660352df18030d1cc5e7686858038a44f43451e1d0b751bdb4bd283aeb2abfd0b1c2f27bcdf06fe594d81a7cc7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h167d3eb6ce8ab52c7da012d0c8103a531e4ccbfe232000f2e6e69d6907b1c68e1cf7460e946288eb22b0e53e4ea6b257d2e6b1856c70427b1c06e1c6a2a5a7a38bf86f0ee971b0ac7ae23ca6e1f6657b3fcecd59cf0fe5831c0703ef0e7f5868f07f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h700bb7be8d255f31f495b67e9fb3d86e04e0363f0d5922634e42a3be785f2c0c5f0ccea7057ae97a0551be9fc63156eddae06adb9ef7d2bac15662e5f592b906e4a6c70810870aed02045698632316bcb7a4c43d1bab0e0f55ac99b723f47d100a28;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha257d7b377d7fd3022dd7dfec402a1f3cb731af388196e8f0c670a8dfdce761cc4d6c8fb2ba3e6342db876878a398d2ef080178ee1127ab92eb2c954b3003be7da498c5d3952e4aa8e52286b13e7057c3f0e1925b02cbe66ba6fa21b0537e1cc7e94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecc18a759de7dabcf7c69b2aa77d0b707f35782b1504eab449d35cf1bf0725f4d9b5dd33b922342c0c6e4d6fa3470cb86cf3193fc629d29cc03172ec436b736d76dd0c878039c092ef7fd864a6c3c4e5b83d94af7ca9231565455c18adfd7698c6ac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc881659c05bf94a0c59c477fa404adee2833cb270ea57caa4a56d458ed1936030738546bf89ef47d013b7354d4f287e6690dbba9fa71fa66b711b9a8bf0ad2aa134650c008c72a5cc991181d45cf667147c45840afbffe4c7b883e3ad26165fc247;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18e23456408ac52c8ad0d17d311389ef3bab5c139f546cf71192d7613827b10844dc8c7fe52d26ebd5e0b9e27b1745d6add4df2c17950d0178d47bfac85eec79f0a2b1520a770f2b76f0c0fbca9f2547fe672672dd30616425ae85ae61a2d479d292;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd5035a65968d8dd20b499e3065cb0a47d38975f872e6457854d9a1dce7bfcb7d80ec427db4a17824aa38d6cb59d4497ad4f52757ee7df3e9ecf8fb17a9c44ca8d6c69c96405d407b38ca03d6e15c7e2a00034f23db5223b36bd323b25a57c2cabbf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e5fae864c5c406d3c53c120dbdd86d072fe956a36a411c71ff7ad22fcf5099d77da01f5391e5481bf9c1a35734d62a8375d580ea292399cba5aec86b54a5664a3a210e29664d44b8914307c5fcef06ba8c2860cf576a550120d6e664c7140a197ca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6828a211f695643d76cb414e567cd3590c4ddea8b58b2566e2bdc19f5ffa578e398f32309cfe8896f38f004d13dc999e99e52d965f6a7eb2873d7e7e52d3c224a4fe81863b0038705516651e2e57d1eaaa2ba7e4d88f4e3e100053eb22d11b3fa9fd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbad22e33cc2dfde60d8574d613f80aa0bd4374c96f50e8209cdaa9d818fded474f8563c2eeae99f9d2b3ccf76ce472ab44610050609cfa60070fe17d50bd609c0cdbb65da122489844a70be34de738f0b5df019c23245959b246d151cbe5641e7e39;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2716d16c7ecc913854b055d60964c8f1d63c87d7e3008336eac87e95257b5a3ef054c75420579262dd5a41b578586455fc0f16e8e6c8c316c51fb4e2a511f1758c1d88fe5035c11cd675381c5ed117e94e0d7d97c5b21ee6375cce27ff8a997ce237;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a6b1be0ea617d1de05066cff62dfe8e3fa23dd4d7b54d1a0fe0001b9cb58e73e509cf6f9f786634cea815971cdcd8e94101e54eaf4ec7fa408398c81ad8f2bd2b4e6a31e9ba870c28d74699d62b23296c80994235f7b9b10997a4b8a209cbf9c162;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c4fc0caa50bf59cb187308adad3d7557037d43c57bb5c6b6516e5e945af34e2668719fc108ca244dba803758e795243d0b28afd1734c4d3d28d614de6f4be6010cdde4fde2cbfb44bb41c390012880d773fb8bf0fda3a4ac6616724710a8289ab3f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h348516cf102ababd8ca088857c1a7588c633a56bdcdc031390c443bd08fbdf2ba18df506737224c12051f311727bbd3f171b6a59346ea77eab1830df4657636434d6e3fda2ccc897797c6730682a9a501e3f34f88cf3253611377d3a8c31c40968c5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2670577f7dc2ae840eaf04b16e499091f514417e6399457c186293832026d90c0023a92d78bf3837cc3468ab8a4f4f0f6b8d035266acedb1e6f3a06ec0c7ac1d53fd47c4feaf68f4018653e53270ea0a004adcb057d0a299b953297b2cb685fadc2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha142c2c8985738cab530b5836ca8e8d73d8d81cd17b66fb49b82231d080bd165a9a48d2466e868a7a7574c0dfb8f8e8e7ac2366f8df529810dc7d990bdddd9805ad0c1d3ee03200cf777d970690746493a1aaa419a7e0b2d4321b3d4f8f5139b1587;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d639747b5c0bb31e5a9aefa1cb8ad420acb7615ab9ec212c07160a94f20b0c47247781d8d135491134cc8b767f11c4cdd95eb08d06230d0b10082c502449a5b24d4652969597980897734bdd58f46c40665d2eca8ac4e91bcedb59bf54776d7bb3e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h405b82216191b0849f9c11f963a0dbbbc8bd27a0ade4c804949eed41150a09c4aa86b3e385b78c55f2bae081713c490df296f35a2657e1d467c29bf813f3cc8dd2878f890d13fb95561295daca50c1c56da3420446ca51f6115ac7d0ded16bcba00e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32ada0bc6e7c0cf770c582effe0796ec0ac1dd39770676515018329a1435a2ba5fad5cba4274b3e08b1e0a8df2523c541032e9c9cba12dcf510128c5208bd63c8ec83bafaf579577fc20f8e383aa7950eec8652398d84687835a1d938cbfc78d3df3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12f5a48527171683f17dd951c85d98c7494aa0f604660665b8076f23e032364c966da21f4de074c656a21d08fc2d706da8cddfaf3cd418d416703462bbc1b98b15b962c5dc5e152987c0b13a0c61cad2c3850d039bb7af12eb80a21e396413ab3934;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h762f756614bf83c93feca951324accbadc5c4e4d9f165ce0bad9dd38101438e58c4bde9de00ea3a7dbcce585363d1fc2f59c4523991d4e6444bb45ac8c72377558ab79c37fbf673386f54c82942f7911ffdc82c1dcd4d7fbf684b10cb9e0e41b6e16;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92685e5e888f89da0c3e93d7a65cf2678f0599aa581b1332e54e4970c56bccb5fbc1f1593116e57b646f52365457521118b5364dad7aceacd3191f3ae8b64e1d1d109562041be6670e2ad9448d46e620017295f94c751a8923701aa998443f0287d5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab173c02f0a24b4e8fd72e1656bde8326e1b7060d6468192b19f41808b4f6fff41d7f11d3709b369604e1b3944b7f6b7a8603843fb8a791b5d49ef973a0a1b7acff9aedb9d587dbbeff086419a0b5027ebeac7d1e3769e8046ff8cf5c90d6f9ab847;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6f9e2077779c91b4350b68b138a3e579a1035f6198d39718a040ad45a729a6feb9753fcb4a7ddab75da4a88dbaca704d9f9daa89b3e438c9fa573f9427b8137e480ef03a04b62fbd77cae8e74b2e0db997eebe5b82ca9963d3e7352b4daba2c2b8f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haeb61d9ee9734e1657102e66b8fe2e85533eeee539f255ba01d055ad8ca473c6df22e45fee64228ac3ada50b5a4e22c8783aec27d4340b086b7bc68f101ec8ab2b17a19d818cb798a5bc0a549043c68a981d5d6c3adf0b672f2aadc7011168fb6aaa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3feb9b272055877cb516c25d44f49c23fe9808f39a59cf1eff430ceb51a4ae038357eae75840220f5554952e3699fec85d7399e519905f4416a788201666292aadb0f0cd35961f99ec43e2437be790f6e904d5c18cb30238b50b38049609bc1898d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8cc18726622ed79b5b4115d2c713fe6742ad63b1e9ae4c7800428e324e25525915ef4cd55ccd5c15d25cb78f176c140f105edac966aef993084bb1b518c086fd414b4fd5efb36df24b79cd557ec5c7d4ddab0c0f28223ee61040f1bcb780be2d458f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h533f0e15a4958756414d7a164ebdcf50e37e883d888aaf671b7c69e7a1a74e136d757c3e87ba2335e5869fe782475f3aaae42d0b24703ff9d0e2cab6765461a4ed760cdec826eb13a6396bf853cf72a71e2f4f3b655df9dc5bfdd033224cf6ce3346;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbdf34136a93e679f6d38ebd5e123d58d907c19424695c4b4b02fec53b3892e3850ffd7fe213212d0f26fde9e4335f73a2c935711fdfae912b796d49e5b3f2e9d4e72a4dcf461f7ab0569ac96985daa0ac76be3cedb0989aee37da5f5d18066f887;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27888364dc0bac8cd65042c1cd36e8f1801310cff33f69509d9ba9cc2b0ee571d46176c1fb269e932a8f36243987595c8acf4a6960f32fdfa6ccec3f64375e3814f893f4cd6916f8ce6776b3e406545ef986aacc4b7253407ffcc2f2685340a85b55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b43f685454048009e7e4123132741db0f5210bfd16c57ed2a5094266ed9b125f753a4dcf27b852c5ac54110746caa366fcb03938c89006f30e4a8ebe397147ba2c370a0deccef9a1490bf153c5bc8806e2fea494ba498902db7b1c27c9e32757f7c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb949d1d3b76c9ab8d008bcbf2c26a3fe5aedfad7f6eee863c164a269abb0d7e025ae1bc496ed9ae13984a75d0c81f5f0b7608415020e86647969971464d56f5f9917a7d2427ab286c5e240581ef831af96b89ed6ddc3f4c7c6b9f0b02a712005edc8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8637de66d9899cd3ee40f73210b51126e7f0432f796551490fd2ca4665228edc4c79d07c52432365370c6f0868eb45408b1e471d51b109b13e57ebad149ae922b5dcd7095cda37d74f3a4686737b861d00225d7005e4a720b6af4cc2daaad32315e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9d7f9e0f67dd061a450d6cec0c9626f4355af0bfa056212fcef1af2006aff60ed1ee406fb98ce7e0c3ede01a13cac0c4295358eb16a4be135025f8a26d5dd023260a84c8c2c53da2b29d86cd65698ae2976008a1d946d7d82445e92c3de4c5a73f5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f169ef79b7102ca24b35cda8a2eeb64b27be7dd60c13cb0dd82abf8636efb3e2dc8a9f44a4f5e59a60b8145e10273c2c6626d201ca4f1d40fc2ca37225055f6d828a41ce12266fe586c04a192ea3e1371c6dcce15a893f4f903d93dd6c18f9bd9d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23e93316442593dc8c96c0d86ec116ee1159469c9a99d7e40292ad628c8a9b7decb8751d98e14b3aebb24078e008a3ca45799007507e80945230be28fdd2f7a32ac526c4f7c215d32c80ebfcedc624b2595001037d4777983a24ad0c5c55574106ee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3974d9e2864b3490a4d9db8284b20b11e44fa5163cab08e9333fc53361685e662b297419538c6fcc263b4058c1055f5773ff0605dfbe649ce2af074a5b0046ed901eea41f6480e17d106a6a4635dd308e98da903a812ae715f5b757014d7187b230d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebbcbb8fd5b6c7d97be9c7ec477f02a4c3c8bc3009a913caaaf24b2461b5cfc1fec7b303f21254a49cdf2e4d20e3ec4f18ae3496c4941146193523f0341d02ff92b505863cb29c64c99a9f91632e00401cef16e5ad282b4fa666fd091a487f3b3be7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a23ebdb6adc25cee7102ace167ad031b3c3b03245d2bcf44db28918a8165d96d62dfa010f4c32d642d57bc829907f4c17dca299cd4af9bbad3f73f123d04da5f88b9373b8961577418abf0f126f0973bb2432f954b8aa2c9b597d41307b44fdc2b8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0a7691a9d643829a8f34fb732e8a4119070aff03a9faa92ca396a54d2863df7370792794e10a1f20e120cf30a65df6547cbb28475b20bf3e50e30f2bc5e69793c13045a01c22a40f9a8795fd36fe78ced5fb326dbc66f0e825301ef7e3d1b0cecd0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a42af08351f0a62479e4df4d3783d847cf99210d8acac0ad55167477ae967e2c5932f8e2c08f7e36ce7e18ca4391c9d8cc7763f7d4986f744073f7dece47cb5be6efdc7101a4cf0d0f983d64998028255cba580ea3b56feafc7d2ea80b71871e895;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h160902b3cfb471f466ab7cdbbd06802218a609ac8108e03f620908c99885f547843778ab2272ad3b16f4440ffec45b7389edfefd9c0858e2a86f46fe94d85b42c33fae5e4ff7b1144edea4b1b7ff1bb40dd44d8ef2cb1e0a585ae0137a6825c29b19;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19108080a912021bdaf738c27a4172da7f9939e6ad083266e15c79bd7955d02f7afc91456651a9f60c902fb95e3c9a2931d75a919bef710df59a5c0f957e799f7db866904c33c39c2622fe0dacee6918e5fb0cc7cce2226de03231eac07120739154;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fa92b41e4e8bab30efe19b5e1664742d3c10bc11c0f35a67cfc489cbc68d0470084da94fa9760835c665061f58d3cf5dbdaaa5ad7149cc4dff46978e3f04c2b58f13f5229d3eeac23d5d8ebcb1a0b5075e3b90bd6a471a09d8965e5d416d6a32c78;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58288e861bce2070b73f831cd163685404b2f421474d838380cb0fe29e9acd5fe1c7b6fe3cdbe31a0c7a19b136fd989e3bfe83c2dfbecf59d8e0d38cfd6c8815cbe44d663018313c07b432a456793a505406478da880b5cb0dde60a34cca7e1b3e8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcb659ff38848d9b9b38674720b954ad0164239dd31e50c835ecf5560cb9a2b1d7d0eeca97be4059d8d576286b8421fa0deadc8ace04d25cce111b24d9243278a4aec6e85b2e7b0aced8a5a9292fcd5dd5ede7ff96d4220059c9448caf106d92df6b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h419d7c533724992f2aae1b51f0aa1ad46643a5acf9314b02f216a040761391a8ad64d5337fd09b44604903b433ca5020690ca2aa0c01188252c73547106f07f92a3d02110bfd4c22f64bbf9bb3631d4e872d6edaa0c8364cac1c6d17a7a9fc34b8ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bc502f4ee96d324877ba5e24a0f8b2d734bd67dec64dcc2d4486371b63955b7d6c08839e5dbb41e35129030570e6c7aaf524e1194c06e20d38f8d3376496e11f43a8ed8a2926a3c4e183acdd81d6a2da2acce0642f6ee3186caef7e4b52a62cef2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f993a827485e0943cffcfb1cf9d1e17db1fdb94a42a783977fdc6c5c0baf34c54d987311df7c6add56795d1c574a2aced5189a1abb7af7748062f774b0188d2e822846c642481c5135138f0b997c96644507afacb393d114913d9f83a4f53f89ade;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83695f4c802f85768a645f130bd8ae5b660da55c8d4bd54594f77a351cc7a4e431548363d957aa5b26e5bd09e8b0b4fc858cef3e4c010cb0670c2c6d6a11b32b580e81a67816fce3cf7f8097410ade0dc2e7cfaaa0ff1392371051177c39c50c3fea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2191f8cb8e0c257b095e0d59f25151655fb160bd5877ee8d0f75483ee0d132ea6edfe00c9b5cfa2ff0a24bb51f57fbd966ef6d5be4ef521e5176b619fb1eba0d6593a9a745c367e0e162d2c1d605ff560d90214322dc6ca7509f1dffa5a44bedac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he02690f99b5ac574560054b76c3224f0a6a07014cefb162fe86a5314557928de7786be25f0b7db82f282d27ab5bb6d1f9f925803f26556fede7b5da8eda0f55afde583160673a308f95e7f6304525e87befa7dfdb03629bfec6381a95a114154149a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c4b2135fbf34ac2dec392f0f16d3b3866f39b1749967810094713d4c9998f43f8d44d4aef626941eb17ffbd2ebf604f3bd8cd07a2ba083dfcdbe52e99a8b77147c9e38ab8ebd1a2e36a074012b9a10334ff41055dbb3190ebed37d271306fa84979;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65717aaef537a03213f36dfecabf7ddf2469e2f824d0b1b5a627f995868592cfcd0e4a3c511c668f81b45b985d879b497dc2d956c12725418d1acb74341dd015ace3016cb7e29a9d5eb21cf14a8c78434f06712b83e0331382d1a1bc8f89278bc463;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d389da3d516d2dd6e321ccacb30659a0557aab1fbdf28a2bc90bbb60d4b4121da0ef0748ebb3beb44d603fd76336d705570cdc9fbfd7c79feae554fbeb313f2e12199da51d61eb498f0df8c5e383a4d20f8d8727a138e64af84281c8025a6cd056;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h477bd5540a50319c9b47c2546ef2ac990d98d29356545d4341f77445852f5d19646103e3b5a052775bb90c42281a316ee4913381875228eebd00d5c8e2777cf01159d30070ffe44a1b48238755f7bc925a8483e26025a65d6a150d1b852b80bcd95d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbaa72a6a0b501dcb907bb202f8fd50c5eeb37b33d0919bfc0033484063cc883575830b701787e7fc8b2fafc01a5e8f0e7781f0a989e34e035176332a84fff4eed2acc88bb7543f9c82f45ae88008673a081f9c2e65f8d649ce1573c83dc87053a808;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5a5583949377d4d5605a240103c6c56c54773a2bb89f802fcf16a3b4f586a80ab6a5fdc86d5dbd3eb9bbc0a78cccb5d3d67cc87446b5fa1cb31eea03a27b1c000c4a501aa69daa46039cb5a0bf8deba484617360ed4413976658f9374665760b0d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56984d08fcd3a9313de0b28cdbaa05fa0e87870ca4e418977d07573e46936b2cf3352c619c0cd8347f9006626106845908c5095c6495782c515de00c3092abdb43718f69c81e8608f120eedef51eb4d8474e50dd77243785d5ae7ff2fb52ac0c986d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25e749a86c562da8fff7455795239b1ee6f689dfa9618ec0c7f606963e9b3b5c066272658d70cb61b986f5604a647ac79db75960b58239813c4d8dd18e581a2d4d2db59da3c89cddb300d83d50599b7d7fe25165a9f4895e672085a78d17eac50d41;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9c2ba823fd720377a1f1e576700aea1c2fb4b2bc5c2ef7cf11594d976f405af8993854efff7c257bd865340aba8f7ed6bc143ed3bfe68110ef38b373f57c9da11ca5cdd3652e392f33e776d02b409e066761087c36f983ef1785b165fe7572ac1cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc95c7e80bed927f256e6676c8538d372ff5079cee7ca9ff977151d8cfc6e14e0c27dac28a3d1e03942bc8f893f65d14c3e8cef1e4f3e835c511eda69c2a32131c0d1678637b8e1c99995408111d4738bbe0997ff116507b3ca44ad5d367db2823ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30bb6dedadb011f7842800b7b3f4590581f682af2db0ccf738cedc7d224c1dcff7bdf338cdf5b1a7e585b236f748484832f4aa536835ffeb0ee462806c4a5a40fc222c27e0ec177b318d4fc9611e4b1d036bbbefc64b34331dd0052d5b3c19dae8fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54169f31bb4714928d69794952697abdc0bcfffb5cd9657eb28df0550e451cd17d60a1288d1021257f97b3ea948caa616df7b2e2261fb01e07466dd054b2f980bbfddf9ef2ba15beb87bf55a04955fe1af62847004bde7435c2beb675e7177e311e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9780b76b84179103f8a7866f50f13097105447371c64eedd45add5111baef31d29b1799a281bc478bd19c15f79d91730a691fa132fd5aead94d1aa0bae20093754c9ec628729f79041a21b5d3e36a5fef0a7fea2de7e17e48b0880a50e806f25f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h269fd51ee9532c96fe00304085a5737abcaea25a82277304fb58aaef696747517c03601c4ca01b3d3e77025def903fbb2220bdcd96ecab005d234445a76f02c61aecc03baf85839f8a9491927b11d92e199d8132bb7f2650194900041573fa032a35;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc14597ded9b092594cb278cb771bed40c0b00644036e27beda1c921a19bd0f19eb947fc826ad71cdba469c0b871b1b04836c742293999911e1e752476c4fe57f42ea3e9e465d55d6068b3b9e323c9865d624e901c39ed39d81aded373cf998b5d16a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4742d31b88d36f985dbf23239308cea1e83f4d6985de2454c18bbf11e0c7567a8e6062b7361262995e9eda03c84aebead177218d36e0fcd05bbebbbd2633ef447295ce1bef138fef0b4f8ab71e19e7ed8dcefda52c61772260611bb9e8061d19051;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62e500cfb57779d7ced73341e8eebc88cb4e09ebf1cc6342ab3e67a8deaf7bc3989d0d01dff74dd59fa7e8a8ef78e8ab494eca9b5fb7863d9a13a958604deb088e5ea529c0d0367308a22329a0bfe84e1ac14bc27a5084c7ff4a94527d02290ccb45;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b2380541ef7986a750d55edfb3412e478419d6ea0bba347e9caae69507c73e1e5db8228ef655d2c4bb99eb4a9def2da8de32ddb6f5543173f92caf6fca9402a440910191b30a074744b1fe7247e0a2093bcdca07ad636b0cf6e1a132e4be94632f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf21b2f33c289467ff86b782dcbd130af07316b81303ddc787eee33910aa8ab42387e6217f68e8eb280bb67b45419b3853fddf984862fd58b622219908ee4b4f6b1649a21d45824f09800e14f888de897aa081c621124d3c758d79288bfa6625c6864;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96b9adc547bf6b6f084ac121034314729bdbe022a74f07ff74dc4801557243cec91bfb60f79d4bf8a7a56973d1404c02c7167cca19de7b2a966e9f299a5bb3487ed7ff679f59c52af5ec886a245ff33418fdef0f470902f6ff9ac66eea103bb0461e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4d44ced5a626535e1ba64b3bd19e7427ee5329f4a293b642f65be8b7600e32697feff05425d89ea2e5282944a4ab5f2b872fecdd0332628f46ca386c247e5c1bb4a21d47d915282568e8404e7841a4deb6348bc7e8ccfc19f14be9757f775a09cc3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46a1bdac7addb03eabe6f2ee3bbe4af75758f393d5e61448019b98442f5b60482a5cceec2f55c6e8eb2ff2e7c044e83fb03663840fbe5320bfb1aae18b9c1f404fbec1f2425e817152829716a75434b7d0b049ccb73c3f49a3c779258a9739a11e85;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc16a7483dd20f8cfc9f23fbaf25a7fb2e1e41d97ed66ab69f80fe8cd4ecd9923ee7d808cd12c57d10090617f4ffcc8392798698d8e378160d542386db4a081ba47bcc7dd4df8e9512660c7bec06d962fef3af21baef0ca095c5a5f6f124112f425c3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hadac048d6d02de264f68d441e92e8f13f0e91d91314a074e51e4f819839f9eed88023dc8effe1197b1077262aa28687a5b11e195e4549e255c0de0195b3b9a057f739d5aa357f201835d0a19401113b9ef4e2e561de5817d63800adf54a0e1501796;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4ed3661f5da1fdbc2309e961fde2efd74a7ca10d7d4e51ff7e77f36aba6585c28b4ece990309780f243e79fc88d24b851b4ac94907bd062c04ae97f159bb39518f3c989eab354d131b9049f18815de7a50fb02ba679d4b91384b816e25b2d981631;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he67679f78253fe8e46c7b13604546937ad81b9b3f0136e432cd343e99e84824c169d76699f9ecc417bb7f1078705bedede6eaae36b0119f8e03624e7279c4cece8ec019da34eab8441fb241aa18d3200e3fa6498db07c2dbdc023c95f7e48484360b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2345e659c5082e3ea1c15c090e045fcec5bd3caba505791437e0e81e0daadfeb80e11f570a1db021268dfc3fe3d6bb0fc2c3181e73a3b8d455133d9e2049ce0f5b9f74c81cdcd3fd34ceadeda6c6aed8401c9272b2606b51a0f002197f8424a8251e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcda7adcbc7dbeebd26678255842904bf98204f5156700a657e684c9140ee876bf41044f8234382ba55414021eb4bdc700fe12c5a5ac0e4786bd03d65d37a10060d95c5869959c2696e13d440b629fe5b1b2d209698493f0cd30b1ae11f6f7623fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb83ea610545e8abab1136ee035968c7e884dcc39ec55a2d088c2fa08202e6714517c033b370dce77f98d0ebd0a5b8dafec719db8a9e39fe90a9ddd8e09a95a440b57c5c5f02baa237a4914d5ebd167cbac837d5765d2fa0fbc74ef29356a852c9f47;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdce5eb2fb4f23a8c7f037b41bb52a72c1c4b8e361368655fa8a735ddca3fc6d029da6bcd462ccac3b8de444fecd6f2124bb0eccbd50bdef8ae8251935c3f5ec1263a5df5ef9169aa6d7bf38fbeea394031788938a42055b0d76e920ac499f3975670;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h937d7883011a9b37edc438f183bc8fb9681fcf64f01413daa25c4ee1c919f4f294d1f8299ac25b9ea9e75aaf947c445db6fb5b7e46f25234f1561c1d8dcbad31ca207ecc80f0f743cc87ec0905570b4838729c3cdd8995bc483e15574a6332bab2a8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd84b9f648559e1538d3955b90e94b7a2464eb577363c7cd7b790d904ecdee4dedb8f6cbcdde812c19967e0d5d54870728c4794201c63c6fc4fe7c62c3bbaacbf539050b3c1199bcb091ff11428bc960280395d1a270869f0b17087459eebdc1b6158;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee44f10950c2905151fc1117fa7f831bf6951a7636e2b315206d208832c6ba1704e483ead7ea518589a6e4220928b8296a30ee95ecf03a430518c40819a15cdc443d480c282a3d57e728e901cd9ee8f6b993a51aa4c3442c5bebb78367cf34aa2c1c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7fc25acbbd4f7df94ebda7cb216438302cdd3081ccd444c02993ecfdc3c89d8148681bc7bf866dddf4fae6ee6d79d75fecc2275b1adff2f9de2f5a4c8742ebae40ef213d905f2fd393636723ed96b47cbf14943630843776f6272bc49d2962372608;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd1dd8690a9c47703d603e83c9c85988843a0e92f316e7dedec05d10e4022e19c95862085e045d398af9c9dbb9950243eb5fe0b34b1ebeb6108f8537fc87031cf6e377097f44925b06e2fdf786096b2c5f0d564438a5b30dcd7438c15d00b14b9850;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc209211a708ff640fc6305385675c40a40197ea9da7448bdd61d2189309215a42ccd1bd8d372f88465786bafa7bf2972af7a8c0c33f1b1e972433bb72fd526d128a60d2401697f1bdf24ba4c67fbc2d08e8db42cce2dd481fcbc41e885a8142ac90;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7528ce65f35fd0bab67cc0329e232223f55948d7cb4eb6a852548463449fd3eface798bf59cadc59e8b02f708dcf53689d6373a543120f281187aae8d2cb586e22a4d897c86c4f9a4031bd0fc08637bc18e8b2fac21ad47489fbbb3b4a67f16049a3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47c9836dfea65a01ebb4d2c365f542c4adfec92ce05d3e198ad659a25e12b72106cec28c721c93e32a0acae2801ceb4ec5e588a761a93f3cb4a3d9407c3fcdf56647a678fd30ecc65d47417c4c65f5f30af468bc6e50d1f8d3ae361e0a162659aa29;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1359a505569be3b3954ccdd740e661586a59ddcdbf6444b3cb5960eed2d136ec1e4af9c6da5acfd891b87630f785ea58a1e03b264bb420b3bd346791ab0d18e0c8c84474715b573ca6f7bd1637efef3f19a87bda15fe125fbbd23ca2f522393db95;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha091e01076d6db1f78fbcb843b25324050967551dc420fe86fa3b7c9d562065c1e8ff19fc9f6072b87af815b5f03673455aaab71dffd1fda1a14e9e2ff365676cbe92c410438ac1d65667bf12feb37ede8a19702b0801a3dd4ccac0ab6571378c1bf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdddfff35758b027be16a9805664a80fbfcd340dd5dc3c5d475435386a512998ddf21707523e8e2c666c02e9c90311dcf1bc3c6e8cefda5a72204f7dfa5d4fdd597d27300c0f1ed90c5cab7b87e281d7e55c984b48a9104bb2915785c30a1cfa833b5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd71ca2f7a3a9fd003bf1e76118c2ebe972ca3f3b99128d2847f8d0598f3d2887c8488c70ed3c753765c139cfd9175431fd42d40220a5e2543eb84112537a5fb270fb70bdf87b07e1205ee65cc0d26c0df1f4637663f9e1d24447eee7db9f169390fb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d88cdd1f8189d047fec4aabd80f5c09b49c8d00bbd36211d3ffffef29a63a7d5777bf22bddf99b5df95d547791bc3f95c0281db154ec51e7c5ca4bb517134cec6b881ee4a5e80fb3c413921c1a9c41ccaaf70688a7a66ea97f80130bdbdace1b958;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h281a75bc710bce3ecfc7e9489c4ca952d476567c994b4ca49724222d2be6f23c67b040d0ba085abbb5fd391ba1a00b91f907ecef7a6800737f673c89df318b0a1bba1cac9ad5c3dc572e6f90ffda6df2a02e1312ee215f57e5e602dd7b78fec6dd59;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23314fe98fe09c9e76eac89d32bb7028ba4c3db392930971ca95539eff383f87d939beb0dcba0fa046d6c5d4ce114a4a5ed5ff8b6ccc94f2ecb6044daee4c4e5201267a52974dca461924c625d680049601641b5ab6d0439bc06757e2cf1d5096274;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc69cfd69e19a282897828e7f326e36337ba1509c1aba391077e30a4f1583ecb8559d483e3eb5d047f79d0744a1b95faded46b2e7d7e76d76963d978413f3cb2736b8da9e07d88df757dce5c8623c26a7c6926076ff841f5d1cf49f217a501769975b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53012161ef6598d81efe46ea01979e02c193936a4605304150d095f0bf58f2b7d1c4336ea12acbb47cdc8450601e88ebd9a74a247037075996dea7dbaa179b041aff059c076793cf3610dc47bc30b0c46bf8635c4a89a6afd20efda8fe371e70efea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9626c5d707f7273aca6edc795e2ed0a84576b04bedf55adfb5e0ace9f481a16f0961901b2155677b60afbabc287e07ea0f371f945508e8bfe83db7ef0004db7d4660c1f3eeffb79b23e0b7d01a7c155773fd7aea08a7bfdb4b8d3f42caf4aee28157;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h386083758d3e501a43cc0e2bd227100b03dbce596b0f4f289717861b6ba61a5d88cd8ad059ed9927c677ff1937c932f5c8f6e656c3f60bc767c8204974e71254e15d136ff026a4de15ba9da3ef2872a576b2ede51dd459dd0cc8675855630a39651a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c9a7c9838b8d724b00a9fc78f3354d41eec710ff9362496fd6f296140052af06535715102f16416385a653c41cb9037283af7908ad8b68317d4ca113eb6914ed11d2792c2ff67decf28e42a9e54f8c28690a0c44ac63fa92f4f0d6f5dc9d9215334;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he47a0a6b4b5047b5633703c04cecadc0b610fd7caa57319fa55ecfa285cab4932a658583f84ef01ab94feff05b29330a96524589d95c0b571b628f96350c6cb6a0b926a7d2e85e04b5533e547bf18901e36377f55fb89111cd783518eb7e3863a1f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcad4237602009e71061453e0c7d04e3725e95192419c5b08a972e192eb95447a803c4a941e78e7b9cd2c42b241b3769187f7914fcdabf88e544fa81ffea59354d7de8f3064fa35779a6a16713089d4f251c000b5ca7c26fa0f5b091360fe9e69b0e9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfd40fd14b900cfd51841c2024fd1305eac4ab319e405c2a45cb7204e33b9fcf544f5daa953267ddc379d6211ed9535ec293c2558fac55dd359ab5f7ea84839522e0ef63f7a544063564c26625fb08ae9ddec6f906e79051ed6a1aff5df06bbce47d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha522a83150a1ddc3a8c8ace05607b0ff651eed7319680047ee2b2a14e0b3d3a38e54ede967428e8a0ced43257c832e9814ff02a8801e84b067299061e4940a86dddf93eab796a91387480baa52d9bd3ee8fd0cae22b9458cbacffd0066a2b01bb345;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6061f1cfd23a65c64b9d1647129b8546830ee56ecb77cdfec11ddf075d03905493537f96f7935e8786f3d9f1761a64cb60a1268f4fb87d210b302bb96dfac5d88b735c4840f5319a26e0a620cc91c1f14419c473db6b145d25a8788a8ea87499010a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdedff2d02b5d1ddffa54a50d8b36be80a184b98a773feda0ab217988d76a5520ad28bf7a989909ecb42ebf0266ad8053e37e4f0a63e36976d82ef0c8582d979e205809d012eed301caac58a79a87c046eff265feaf10950cfc59817b4ad584faba21;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a208165b7571cd142c1d824a7910b62cf450d6bb08115262dd3c3055d0685fb50db78eb57b31befac10eac55a918a11a0a87c5b3e89b2a84b6dc3dad9426700b6f2df0230b59d91e697805b02f8b7f37cd15baa651c132e31376cd09e4037cc1d07;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94e1276c02984709430cd4f40d9cab00a104d1e32ebdaa29df6f611fb647022d65fdaf769edd091371f205a27b78cfa4488e2d684afc15a97dc5945c92e731bef7e5c6415eb2d3dba0c6ab845d98bc7b283c532dbf79043b7969a6f632b9fc900e44;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28dcc89bee12f53b8a029bbb5f845952d16d9ac0134a72c06588f9c33f41cfe7cb5559cd5abb65089c541be8eb7b86a379eacf84b59c91d348521d5c2711adf3f3eb90bc9911cc0356722e1110f8a80d2067ecb30f574f45d1ee80086264b6a4f3f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ca0e41d5c0e0fd7ae0cac6e3abc6f9c848d9c3e42b7160e9b37e845154c561cc583bfa91a44ae723c2317d6af01142eebf07cb672f533a754f8ed260f54a8a790c240ecd79c8f766a81f9c3b1b1cdf7cdbbc1dd9a4b7a733e5e6ab5e260d50fe54f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1eb943d8b3a9a9b749a3dd28aec6018672c62171be6117bea6101ab908091864a022a6bcbcd7424414021bc50db6beae4c169dda490f611d95720973a0e2c8c7ddd191b8f9c62e5a2ad38098cbea139ab7c1d07dc8ea824d65e50698a597c6903fb8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h380edf1f7759ffb2b4463828bc7a5606a1f749fcd1a58ec13bc4e423b8c932d481fc740358a1d7601f4437ff3f88da303071e5734479df6bdca47cf535caaad58367045d9b7bafd934a18d5734c8e73fb48f0cd95f73524f3b8232cd038e6af3734;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefbc46229850a190cc8b14ab1ec3b3008181e2e8b5b4a9ef59bd9b774c10fa6af5f0ae9b022707e25c36a1c51989bc8bb0200f0e44507bad8c29c86d61ef3097590e74e77974f2bf03477adc28e506f2c97b8252cdeb74ef7143fb7e4052b811d9f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h823f1e26f3ed137607ef0622741ef00e52739a12fd04348e5f154653a78fbee80bddcd83ac2c3e64343a7c4cb4acbaac6912832d8cd05a9955a441528a461c35b72e149b9d7f6a3dfd0c3618c9a19335a254dd9830616ed3c4c60a1ac3a32dd81839;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he671e1c0eb54c94510677329328e16a3133636f23e06dd684b646592927800881449c260bd5152e15419477b46482dad4a1270782689e7023cf1588088d61bc80a28fbb920a05564d1dfc245b0ad8a648c1b133300db19602dd6486b7574a43ce003;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d994e854812a18331f0acbd3967ec5a0bb3ae035dabd7c075ae0131e380e13c388ead31be9508b224d0313a741d69d0d632f75d97f41e52c7fef8f7006fd9136c2887e19528c46293412682f881c420307e03b2ee7d81f2c46c9c89768c932da014;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0d96b221f7f0e737b761f14d081cc8e274581785d89ad7a081360fa6e6ddd488e6401597dc65e0c7f79d02a9aca4a8fafd664f9fa22cc5ee1f3d526a6d0d143257ba90a5b71e5d1b3fdffc5d8ff62cc8674bc1c320fa8ddba75a82b331358284e5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffbedab6d042f87505725efbc486927d1655dc5ba4849dfecc6f64475e254e09ccaf084d281cf03ea017560ae4c5285e3c03c7fd37d5ea20d3c6ecaa4b080009d0b223e822ab469af9a746ebc2c01bc811196e85a04af2d1ec02b9b910222e8c8cd5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc34c63e2ca53025c2c4e4eec42bb1f839f5b8bcd082e6f782d7ff827670c3300a64c1362073419d6a5aaf325e282e7899c02596702cfc1bf896169ec1544ae7e63c970d74a374a3800cdc75007c5d7d3a8768b51525691b9b26e4ee9d0e949ec61;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73bcafc962d25c4063a5f970e85f07ba0c1e2369ff06cdaf07488a6b2b61ffb7baa3b5885778db931599e5d95c9ccaa1f3d09927f45aca8a2cbd613ce5ccfa52fc13cdb8e5b73535117e4bc00370c624c6c845d8d26d434f8a545f391fa1f48c79a8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78721fcfbb810e6edfbb577ab05041e31ceaf797a7fc94d995796e01fa24f29e92b4117f666ba44ffadb6f1cdedb7a2cfcae4bbc4156af087338abf80adadd679462f88480bbb50a3125d46f229de8503129d91296225718d538cdd693c8694a8d3e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h687f08648060b1696178aec2bfaf3f9b6e4aaf0ef8ada832375d92618502eba6c4ababa8ec0a16695a8cd9c71645246b73029d49ea43b75f43937e1d773a0bc762b8067238e124c60e26853565fc1af5a7a5e8d293d8602384d4fecf318feb739e66;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4b559f9be9536b376b70bebd4ca28c495c5de9a0e96d4d6e4e9eacd7205e628fb81ffd65be702aa62697e36a55d1d1265606025e0d766630702fcc83da59b1c74d55247d58291c5288cecefa0cf67b852a41f4a56d666959c51f4404054f70bba81;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99180d8650e849d09a4b41d23c30e4d7c56e51d63528317679e829c441cc19ee165d4d9c3f33f4889c37435082aa3b9f4b1bd86c6950f9d1e2f835ad9f26d121c2e35baf75b07f70cf89c77b6de69567db2d08d98c5c175e85c749ad8fc3671dcd3b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e56d2cac7bc67efd42746cee0ed863882fae656096e0662d6c6f0b5b9083520391d9c0db23483b9da2b08bf35d0f356cc373af9f02837006af7a7ee7b12835416e7bf77c73439a57b2c56b48a3f3662e810e8b2855e18c01cf6c29e6d65f1499858;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h212fea215d45ac6f368dca64e1155799a2fd234915fe034d896f2f447242e67acac5a6a855f8dbc952e5cbe4615783a892aa54e591106a6fc1824acb036a999d21b55dc37de4127e6c8159d06a95fdf373402c4c378f1b46538f58040f27c987c24f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e0cb01274ec3513d7cebcc25227a339d684bea14edae0cc9ab4eb671d98f4a3bf3ff3410ccede35a704c059682d24ce671cfbc2847895e924b11b18bf72e75a24128283b82cea34b9b6d865d2e2b833bd7bdfb878c09639059791fd6b3d042707f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe98057b784d266399877aeed98b9a3e791b84032806c70d926d369f70babe8dc4bd7dd1deb89b66da944b57c10f4d0f877213ea1d853f6a97152bcbbb222b2c3a5092d3e1ce1030e451bb2a6eb7c9a24f1b8b84f06e2a2e3ba3d9b81f3b7582468e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habab8c7f3d8c81260337c9f93be7958d4fe6c6f1ddb16167f442a580710fdd526d272c4fe7548cc44536c8b2c371826b8b6c5652580f46b0a229958a312f3a933f28620ee65e012cb7e18c2e8dcdc598e20b3500385ef201e4096bbc164654c7ea2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3268af4817d2dcaa71e8f0d4f0ded7a6ade7eec5206c421ba90b8f5b32992449584e90cf4b2428998fbe2917e43f27b46a2ea998e6ba0d5958f1a51cf0dffc4f887f9bf0cff3dcbd9bc1104a1ef8196ec06c7bd87be504f424f6c5ece81f563036fb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79c111892fea9e8f3814f90c51867855ba617fc6d24fcc2245fddf76388cba62b6786278d79be171377dfd54dd7070213c50e84d818d319c79ab207430080abdb621df8897804b31be131658f98596b458068a0476d293ceab944491213abad197d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86171f10ffecfe7efc409d03e5f58d74306f69958c2909c056c3ca9bade67699f5b00ae0222f4ade96b67b819ae3773cfee2b10047fe811749774a40992aa34820e99694fcb4146b8df5dc8ec3660f66e491f0615c1cdda88f9f68e615d41636eb33;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8abd3151234e2badb88a3d4f1fb3c7788ba9f4c22c7fd767601e296fa1729973b465f5f33a5dc27a138d41fa4e2af5688bad5760b9af6f194af67744c1cd4576de16f5da296bd9c4210b63de522ca0d8a5da55f6e48de759541300bb9b383d6c655;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7445fb114abd0d78aea1cea2e46a63248f8311aecf124613e18d6fe0f7101e38489d4e23339ec1e9967fb79245b0114206bc1982957a40659700088422ee838ffec3565fa113776209e2fa0d91ceacb0a808d72ffe303daade37bfbc7a6661849c9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha898466d49e5319e768faf814851b4f3bfacc2c13d7873c35e0bb12840cf3d27c28c267ee196dc2825ed36087573fa44391b0ab86f545e11ec5c1bfa9d58ebcc2ac057af6507773d71adb1f10ad252c971da6da65248a991f7f64f9135729f3fbafc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffa9eb047443356ec4ad283bf8de8289f23ff4065442f8928860b6d498f00abb0caf5ee1c43f6f9b2983fe46635a435ad258a7eb6fd87a31ad5e2f014f3d276829d991e0579b36053fc3ac235192e71cece4b2a4dfe5509dec311c4884c50910239f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbad4b593a2fe8ffcd6511fb051e05b3a6538c6dd8970f7e66b56590b5ebd3d9ad0701a25feaac55f037ce9f1863d33d93f5b7898f419dc504ed09cd27420f00da9d97f27f2cf1a66d6dd5ce3fb8d727d4b0d25a976db03bfcec188cbb7a9140fb5e6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0713c128494291d29f49cb4090d05e002ed18c838a9b9ca63da6981c3fbb6c50b3a6b47f8e41e79146ce59f17980e717a73b25fefc8ee3848f99a60d0bf6db4d4260a15a8101c0f7a9c7ccb2cd1d41bafb7fe87ec06597fe246caf7c6e5e9bfcdd3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79222cb241f675127fdc869e878ab3dd926f03eeae756dacc062ed4ee4f631a9553bbb2ba31651464f9ef6d2557a2622ddc2cb8631e1bd513b84d68ecb0ca33b9e8e4abe4c9ebdce4a15338ae77117d56ccf281b1d431cc37f71c0ec3f74341d8e9e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84c6979f4dd430d09e683ec2cdcaaebffe96c2e6a04bd88d16b365b85793f8eca1bd0aaf692162eb6823b9dfb12d6cd7c75c304b8b87454644b128deb6b54ec12b74dfb2ac2fdacba9324b2aabf9b1e290bf8238f9088b5accb33d5d07a7271f6ee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd95a846b24839e3f196c9ac75605ce259f63b3b42fa775dcdc2d8b00fafee1a75066d464f9a5e7f2849eadfbc8bdf6722c4fd403e6f57367b5e642b237c12e09c1c27b5f542e13aae1e6629fe5314827a9d0c83fba81d6fee9493f3e7695e86fa259;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h936c5f3a35efa6764d2f66a6c8eafde6d540a86965c7f088fc9040538dd9dccea7cb0824d6d6d270d3eba0ce146ff4b6a46a5880c4c27df0801104c4661b8a1ae8cd7093ddbe97b581ea86254e1c34229e4c6fe02c7fd80364dfa7da7ec80f98dc25;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8789faac69116ec67ee57de55cb9d94babfcd64b1251109051cf34735134c51581ec5326029c86300fe51e62768a07092c796234201dcf58c567321a5d35e09cd65384522efaf3ac97012432f27dcd8f55899be002fed6a4a4f4b11034f84596735f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha55dbf7a157d1cc031f10b078918d1480db66c9442922213cff305eb4334858a122f6ceea5f5951a9329414ace7cddffb4485a669c0caaaa168face797df48ed13f242770191c64b4915f8b1ccfa759bf24dc2d5c5571b2c46b39f1fbeafb753cd68;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he20ebce999ecea65bd1a3bca72fd7b440d17520f66bd10368b3f09f7d08ff766e3ce5f5539ee0a6b2e1a00e519a684dbc2470bea705f894816cf464e8c192adad2e913cb0b8954e40678a229f266e91f24860b5a166e6566b15282ee16ed6475b202;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2de46b15d34358b196e85f2c12e9fba054c471fb896e267e4350af5b96a6e2e57c4bc64faa89e234d5d8d58f0063a2ab24e915aa89b14c91318e95857f49ab44c83e2658fdd8e3a420f2c08cf2316ff57002f59d59b4307e56f370f23f63dfc597a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb4c20728380686d28569a979cbc71b7cb8da07906380f56895ef89f34ee72dcddfacb74a8201a823ede34080c6b44cdb4c7f14f032bf50e7324517db8c315cd3fdbf49fbeb117b2b82680445f27d54b716b1d07dfff972f59540073a49ee2a42374;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf31be93fb52163bccc69aaed8240d93c5bb702e271978670ce6f171a8150d7146a02947acc9c408d188060c87b525868d2ba239cc8e601cec670280a0b4f8935eca7d62761114794333ce6eb6415be25f5af518a348137c7862416d2be29e8c0f7b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71154ce54c0eecd9dcce669b0b7cb96b4cf12cda4f443d62492cff66d4e68b81981ed55ad56f83e13cb7dfd83284d89919a006edf56e66627061104456be97765fbd77cee7d565b1394d4759abbb6b523f336fad2478139c080cdcf035ed6b9a2d6c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fd379e958cf2abd306759e42024dfc96e6a379a9a90d10ae182e56a6fe337a91761496a4bacb50ede4284d2793ef0e6af4688d843372316eff5847b8d8f8030a0bc10e77fe8533014174c6215810c63f59f8714f980d1975b7cf24792cc9bce780a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a0c79fbfb5b6d8bf8b7d6ffc9ce659ba24355842cae782c38c4e51092cae9f3ed7ef36148ba52d1aa14813e88be5f1ee314ff7ee9b116c9ac2ec7509b78cc2d7a37aa8c2648029591338c881fee5a305c557b3f9a9b0a55c54a469fa5daf73e4c52;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf40e8e46edea6b9722ece3e4b7076e15d8adb99b135548d54df445dbb63d1265727b76ac8212eca4ca8f06ae5d28e5bcdf940b0e562d4a65c1759ccb61b969e417e74c415f29911c7be8c661875cb157369b1f8c13604caebbf8a3568ebc758758fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf41312feb2225bd6bd9829d0beac42230205428b7c2a111c8bac7b70cbd43c37ca70750360ddd47cd3accccd0a3473716072ad80543a94203b70f6612142eda8a93d44e51b695b8f48f851b6c47788d01a98cd4dfd80d6035913b31a21f256bbc63;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7537bae2cc2df6463efeee5b0c5470da419d381de69469975dc1876e1048c62f3ea28ae6083bd8dcd4639af9b1afd82e597269a6713f465b1d60f36bd87a85510c1cd1278bb64a606f0edcb2dcd08c94ed904cbb79e7e0b8eaf28a5a01e81056f02a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf347db8baf94f22dd5e34da5c44d92c954354ea972aafb2891ab06bbc15380bb40de1e097a8adadd5de67715a53f26d1c32126456a3228ecceff8b5fcb67b38b7733f4e2faf83b2dc8b43693a7c41f3fb9f05d80776b618c23972d1416180375e013;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4066e5b5a7f2a1138e2aae68cdfa3613bbd9efb32d8f170895c42ee6742995bee3a7998a5307285f279ad7d3eb9734c1245035b09ab2ca69ddc75c907848d522a6c4daaad5cb76aa056bb529542e2d8a73835e53fcac2e262469ad1ff2f3addffba7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52a97077bab7a9de78db5fbaafc2f59eda5478d5ffa61538ba148f6b4dfb9e1ff70ec6cef6d13cd3c391db6f436529cc5bde074355df522a456551798e8737ac133995d719ef123c4c50b89f3d6e263665a6ef601cbe6b605d88c61f1f7ac73dc1e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dd8a730d0d53f25bac2b39a92463751542ada8e11d7e67a68bcc3becf8969bccb90334b4f81d34495fef927e8db9b367480caf8c3af6cd01678fd8d699106cca5a5b43836d30b19c6ca3aab5ee2d3206d810ffa5972084d67bd42e418ed133350a7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb50d25a25223aadbcba9779aeab66f3f56d6bcf57b0afd74fbb43105d3cc01d7cc6b96e387494c51658e123c3e60c432553c3b605667b5576f19954406afe17dfe4eb0987aed7b055d91d6fc9092a60c1a98dc133e16e50d6bb4877ccd58a06e9671;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9d032d1fe5213cc3f878e7bee1e045e661758f29575ef5a3ee79597922555a47213422d6b9fe239f6e5c37290d6e9afb2fe2a3c0cce750f992b36d43a67410173ff621a1a2d64dcfba13b70c9db0c35b8121bcb4b17237497a85a8ea5848139c90;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62213e39dad2a442df3afce8b468af007e205ee30ee86521027792335c5f0cef1247426ade04d247caecb18b52d123b4539a70d7eb607d3d96bd9922069e298bf4464bff0d103cd113f7bff4cec2eac6a243d4a9a2ebf05cd5a2ef7f45ac526c922f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70025253b701dc158d8b7f8d5b2b9d9b0be85e8201ba1ff674f538c777999e7caddffc88fd93a5c23608eb8527081c94657ca704743a09fc6387965ab84934ecf0ba737055827d81cb46e18ad6f35e1b3b8184d7fbcb4906e3dc15cf05e5ece0493b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78ef8ed4fdd6590332ae04d3083b0bd0cd00f9eeeb3b11a6304170c8ff1560d3f9a36ad3c709c1007fe3a080f5a8c2a8969c17550c39e24f20f9c31e83a15ced3bb5bb3464ffc1deb574ed7142e04f39b8cc016f834fda47cd26016310fe59f45785;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3816fad0ab65f012f6728a9c5cfeb2c5a886043d0ac58a96ee6f1dd06e8622e6cb6dce739912cac1153bc1700426bba7abbf9ca80fd0926aaf17b49efe7e6e91e6d41d01c46c99a3daa2ea8c9446b853014d50bf6a3fddf6578de8f0b41e8b3da54;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hedd2b40a6cf610b61800cc4b74ff4605432cf066a02ccd766ab581f95acdf915d88e8c494240bf0d2216e8cc57836ceb82748648148c0c77db15f1b479384b934314e87957ce0d12b26499a85ff0d490ec219e709f2f9f584e27143fb1867822df4b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heddd937c21a1031fb8c8402c95e422748f7971213a50374cb52dcc3170b2fc589932501854541d244f6e1aea58358d4cce22c9e1818f1cf5731370005c5efa957bbf5f344d8299abfe86f353d786fd9016db422f256fdd404f433c2aea45c74af363;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14796ac903d4e910273ef2f10ea988560355c05f68859b1a85d417dbe856defe316f3f45b06962bffcfa1f2a4f06a6e21ab98e7e8c155939641dccea80b0df5f0c73a87050150c7dfcd116946d65fae5642d61a7dcb37dede0f5a5a94f69d0dbe0ca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h452c1520cda075cfcdd7eff5e662c161f633c564ad253b8427fa8b20ec291629f5e96ae5c2ac68c87642aff65a7ffb70dfe1943dc593080ea7fc0a7cdb7d420fad00a28df424ac19c039f714c7a7b96a451cda0cbe70b6360e131f2af06454c5b70c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5203e5c22afdd977897a5afe9a716a121bb5e636a1808da43b9e41abee427402288830dfde4e13dc3d93304399523ed9b3afd395252da29eef7a171525afc2e56c17ef16b4baa7612fccd3f2e4fd84b370953cfb2ba5ead32813b56815b60e25bd10;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0d56eead9e95f375a3320cfca65b70180978951d3614cdb4327d7cf59ab4d04c572ceaaac7a0c2b9eb8596d1a0d13fbd08f6b07611f53568c1da060ee3dab4b71f105b1768b2876392ae14fdedd42d8c8ab56c27cf8c5274a67793475aa7ec89387;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a712153b77fb39fb2063dfee5d0949ba1e0e1aa6bf220c396b004152e11cd896e8ac89d1d53757032d5ff5627bc441dd0ce1d67baacbb176447086d5823d67ad01ee11252e1d6f52cf9c740669c4968184475a8135dfcc042bb01499ff7a5978007;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ad0c4127f7f5db8fc695ba1d3e759e8f5b11f2c9d9f2430b119e39db94a034d6b2e4a7ffe80576062613ae453069e06e0100ed51e15416eae5cafd5074f748e77b9149a634b34134f390371d14eb60dc8344207334f514eecf04b4816dd7c0271a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc22114beb35cce3d8745f6aef06f7e756b5bdcffa6001a49021e80f10f4f7c0effb8dc8882566ef8b8946dfd2515dac78a74d9ce36b71b498f84546dce2e7d4f325b4875684350a7d0aac21e35315fb16849475c735989cc94eab383dda3c2d7837e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h232f854e7c897ea1d7d82835dc4ffcbfc2c3f1b2421b3b13f74c02f7f3ac8c31166ebdc0c130ada756bc25f07b31e780e61ce7e25880543fa8ec44a1f6f489c42200e02c2fd8cdf2870840a855b37bd59bb2099a56a74a9b61341f3f2e43da9037af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7477d59cc22f1ce28b8a0bfd04718298e10ebf83795704cd0f9fb8c9214f3da2a96bdf972c8d01c3548977b0b9cc83daa462b65009ed577dd2966fb80c17139c570acf29b9b6f0fa474273a7af20568c3ac9b1e14e6ff4310ea26323b401973ac38;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c234abf3495ccab44b211c04242b49043d9a502c03159f64713dec4aa0a3cf433c759395884d4cb91431ad0ded2d17326f1eeeca8e720101201f19f324091b377db58f4e6e630105b1dfbb2486ee059658fd3b196ef9e227072e983cc380e13f9e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c9c1473c478e76530fa71fac2478d7e612501f8d8e488d1fb3070c1a60f5c3a154e4231741cd4d14d430487114a25111239b0082fb5b4729d4815b0664c3da1bd6cf447dbc8e3f432c308b0c0ae1fc0f8a2cde304f3af629fd8e7b8f801d0320ef6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h857236142524b42762b50e6ba81492e02e3578963f84498ea2c7c7f29405c1bd56b4ede681eaf5e3a52bbd78e3189c3dfef6851457a0aef52b4dd01c05f7a1a6fe7b881afa967c29a4de0f6df4fbc0f04550dc30712cdd3e02934f0e8550f6abdc50;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdca615a783849c2cadfe13615f4d9cb67cba4fe32652b6a2a133e5b2e8420941f4703cb8b0e07c7d3f925638c50948c3b72f3aa131a21314a515576b9da76427646093e4caa9b503e0b01315369de36d27765e8bb945a4c18d4b4638772442d8ab3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6267d4fc81fe1889e5316afb0ffed3e58ed1abcc641d528915aaa7de38330a2af8647d86f998622d50d6ff8a5bddc4cbbd51355ae1390cae33157df0e5dcbfb896e4e8c188c805cb7447b8d0db670cc6dc5763c47a6ac2c31dc2878f446df9683f64;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67b23262f0c4ab0b0060c4089ea88d06addce50936388ea5cb3a7199305c585a173b55c70645b4f42ecc0fcc36f25ea7850d94609c55ba47e552b115c105577c7b711bd2f30ccdbc377b0fb8d84d9bfbd455c4b023d3b30ad864a8e0afa6eb73c6b4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf6dbe0ae6d305bdad1e380f9be560561966cbcfa6d5c62b498777082ef6cd46a2f7877a400304272a8ee1e7ee0da3471038524bfabdf5c19b6513993726cbe809f5c012ed2dd34bea4df6d66fc8afef592705a39e847b6f65cbc52e69604b6c9cd9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha90bf3f87253ec2e4be81182c4dc9bf97ca24a117ee18de3445f3ac3fba4c23e6f6251a60bb4d477abe260f80d32741ae5a8c9949e0595104f351beb74ca38cf52b26b5a734f260e0d50ce2d22a3dfe1c745d6e39c9842bbf135d909255fc84340c4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4c63d2982b68895bf46af7888c7b149c8e2a72ca1c014d504c8fa78716543e91673a7a939e3e0bb4b4d61a7ef7f4c0a89c8591a789ab6b9e79ec7372bca9b03fe6207339280e64fc8971f03738073cd110daff6f9975958732d3f3a062ab6067b25;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55b3228a4ce66f0999d6d108f106d4266c6e7072a3869b3169ea689c02a3516564b4646132f71db00281cc67294615924e871bfbe8efb96db50b9b19ca64308a6b8ba7c454a3ed74c2f8434614205227ad2d394f29b00dcf69279c4210e9fd21ebfe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc01008c197d603e0ddca1d25baa6a21a39657c256f11601c183ef093d6f6263a803b13c0432e4024dec316c907b92024d40c1dcc2644ca17735855098c11b86c92efcf2d54a8a8bad32f1e7d0c2472741a3ebe0474f73270dbd0413e121ca3dada8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb96909b09d8ebc0f4a603969b9c3636b28a3686fe310195eed219016b7b7afc14c819804d985471a561d3eccfab33abe140a5442b7bbe8d80663e49c9833c61ad0cb40e2d61a9ff7ba6bb4c9b87d85aaecc972869c932e77c48adfa1320b3a1c197;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11852fd122f29ff8bae995eed8ef57901e50ed5d80d9b1f573478a5297300f986d2934768da53d3d22c19c38a06f5d81803de75461969c2262f18fca6b92a66cc9958385f5bf6ab2961b6325123231deea3322e1f4e2c46b55084a1576bbad7a5f3e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf320e8bea6ff1cdaad744c1d42973b12f68a2a593d1662472b15a357f61b5c8f1eea7c1e873931de56e707f6035143d3b40ddbef66281d9eac8887eab04be081dedbf3f4ae39a17ccd46c4791d13f41fd3f0c76422f66e9159896d84a3802570d466;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62a30b6a285fdb7c06ed5c2404924a9c39588eab7f4a96335cbff5554554b4c6c4724d8b81983f2dd314cf28eb4615e335b6e4b61a355b1eb40fe2e653f9d5c5bb72b9b89cc4481398ce34d8e270af90bfba1f7907a7e22ed5492d42e60f878de50b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7172d9ff206a6b66fd60752f38f16fc34491cfba7bb76dad07af9e6c1dcffac156e66ce141b79bd6600b34d1a6bb242cb0505240efdaecfca80507ae4c0f489cd268e1377ac0b5a8cfe1dab20233f29280d6c047e698c9da96ff4a99e93a209c74e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha27c8e122af2ef47ed62f7a40d5783c842a5a7f6cad8ccb9c4358b770bc92ab39385a0b8afb9b3caa520c421b839f19699d60ee0e77ce9454f064b36d66a0b3ea812f88469774bd19728b23d5445430ce8e4592a473f3db268b922167f998817a7f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd77733e8a85acb979fd63742daa5ca8254824c9630943d6c8960985b3b2a9a66a69580b882d9bd14a93832f717ff8b9a33adbfce022f1efb174e6de4823c9ab9327a57e56692e527070fb4c9e30da4de45bab492dd92c7ec6eb23b555c461e4544dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18361d31633223c2636a9cbcc58cfdfb8819854d6384b1d66e686785e2f65d210a87e5a65747cd64075b03548220453d5351a814865884d52e5f6632d8b5d55c306aaaef84146fe46d1bdc35fc315ef6350168dd22272546d9cbb0cae3ea096c91fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbd2aefab9ce4e20de891af98068fcbdcb6f8dd2b3ff20f55c3c838a404d482d59108c08da9927e41f6ecab13fd31596e3e289ab20a90e513ad8743da5e9081a796d3f4dcca2ac0179aa10bd677ed1214372a4c449425510173afd8909536baa68c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b1a23f75e97dba588b0d4678598dca016883eafdc1c3044de20658a8bef4a452d2d80d558c4af63a7fd2e8f04825881de4102a57ca082eb059a29fc9d5d21f1cfa84c04bf44cfed687b555b656718f0afb188409f634d57a8d0e80b518667c9961e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72569c3b31f49023d15da3c012f1e36d065b02acdf5e91a9abcc6d547055f2fbbfd87ef6b5f34b036a8ef2c23195f18f52720df7c89a611406ad578964c1ec31a9171f2537c171ad1be6af77779942ba5171c7816b7419f6444d9177b97b270c6d51;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ac7065a40e60dc6ff9fe15935f1c88b94a82b888fc9d9850e4372bb312b11245867bdb45eec7ba1ac5c94258732bb07ec8e9606220bae7f6a9c4f9afbf4fea908940b37aca3e80bf88ffd89bf5849075ba1fa43ac97d4375617b629fce2e2207752;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1f658da91b6bfc3551404345fcc221e7381e1f24105b6ab4a463484e14f37b9c78b8f9b3e378ea1604a104bc6821f7bb75fc771f021100f7e910e1ce71d311a46aa1bbdedd454b610e9e63994e1ec018a13c9c6617a50b61f0aad8ff77ed6d11fb7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3f8303e3bae12b768f486068228135c94dcd13f67425af508d526701e0363b835232ecc2b8e578a871a59f8d88a7ba07c12b54ef81357bec6fc0589c4128e99e8a45473a89ce4dc3599d3703e86dbb90102eb11c784ba2ae9754fe9695c8343cc6f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67773e6acc1664162a828f46af4744e87c79be21a5b94042394677179ccda30c72aee529fc716c26b15fbb09172459930ff4e9e1da3674243ba86b6a2f4306fe9b409a9ff8eb1efec33ab73b04982465ac7f598cce536428fac4a623ba97a66c5404;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddf124d9f52a45fafa5446afdc2924f437abfcdf42e2486e650ef62f05d9804aee84c07961bb5cea1eb1f1476b9c733378d75795f1a5f4543303912500465dff75ff35567e14a9509b1849d573b1725b86bc7dac4de9153c74c7a409ce74f011f099;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcdf43edd484f223a9281ebf90e4b0011acdb8e53d48cdbac047bdfc1f98e48541006f094bfe598c14bc0644e753a5f7161a2cfb884bf8cd2a509ddd05c4cf080b4effe5d7f14ac38f1500baecddd74b8a8acf24669dc13e73029e848c32351be7531;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18f813061cddae32f076a015a366911fd09055005066af7ca8ff1f8144d3b79ea7352ff84377e51605d0c89a3c8b10e8e67107f4abba648c5e66ada6abdf1698d87433ce158112e875ea30be12b799c849a00711d6ed9228612423fb17870eaf2c6d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3e10080698beb61a4b0541fe13000a7d818906164564c9fdf2c0a0ba69a13b623820daa1a39075e7bf17719680dea9aaa88ed8e3f2e053145f83a3e76669900197646f48f0b8138859c8a8d84f28ad7ffd7099af41e46f49336ac0778442e55b5c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f29a20ea0cfad8a7d3952e670145f9bb8c17cb7d1127f2c0856a6cad8369cd6f81a5a3b48f5a6baa6e7f67bbaf6178abbd1aca36ada558d45e6d9eef3dd4c701eb1902d89638edf5378ad758a8cb46ca1b196462a98abbd7f4fe5cb4dc8d18f7372;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4d12d0c843b1b19aa84450494941dc68f1dc4ee600682ca9d3c558a744ec064bd7ea2a80af4a3361b2f03803292114432ce1313438f30d6edba6e45236d6272d851182d6930997172aed20f9a35e011fff08bb93727275ab9c60ede04308efb17d5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f6dd91689eba1eedad0b9d409ad24d513fa2522bfb80f9848dabccdf5ceba04c7f5184a4a8e5fd99e6bcc245eea5e8d967e366e1250a3b3a87dcc92df6a383e138b28337fc499d269c7f46fbc270761cbd563eeec2a720cd81a0603f0c71766a290;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0e788d2c667735d3fbd24cf83495614512e7f0038f67477953a3614cbcc95013a132a8cced65fd0fd6b1560637da62eadcc8e6d482517bfb5537da69941f5619ef38bfda2bf7987f60cb8dcd353f22c30e3ec256f070672ce5ddb0230c419912e6e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2ea1cd3b892727e11ce8df16d322d161a1867eb1e9537b838e16185dbd671c8197b7a47a06e06d27eca3e6ea32d798d952414e93be38b6a5df44a102e4dfbfc83964130546e42a3d97726c49b40024201ac620e7c98424ba09e5031323db3cd32d6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2010780bae271e36e2e676d0a871f6c0664f6558ac5222ecbb663a66029199a5446e49b577b9e411981a2723739ed496da18f8d31b8a9f9b4874bc2e7f5ba7cc537d0fe5c5b826d14a6ed3a6b6d3afd800a4ed77892a0f36a5e3d17374d5df148ada;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b56a00e9cc35fa93eaca640c0158b3b2e01469d5327414522a9e8e7ab79d966ae600e8cdebc63998ab7f0df687f4e14327526c74eaf79bd83f65cfcddae87076ff1e7b5f13bc88abad2736f8231857bad0e01ebd19b74ae85c60ed34624a5bb953f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa205dbb019bef5e50e2e7520e15aa2e7c690aa66ecc2a932a5a1c22814db83858b464cc634721c61979014fe720ce43e804dd90e048511008f90275f1e29e137caf8f065b2fcee462a7a98858c94a11ba1da8ffb9e06a883b4f8e83a3d5d97d67d1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b6c59a1f2307d73d4b26b1eaac19b15dabb700f289b1ea8671de8240710aadd1999723292683febcb862716764e2a920c4d06d4b347ef308fec396982e75a7243accaec553f7fb550892b167ba71179088d1fcce8b89b0891c91cb3f65d110cd762;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hace2944bf0082a7f7275e73f0c59fec901f16b1cbee690dd6d4110dc341024d27e706a43ac3acf75e2c0e9436e3f8ed80b205a70e394d422421596b0ab260fc056f239149371bd8f702f2ef8fa484dc1f1daf549709b009f1182bbab24e65815075b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeae02608a895e89d6fb416c096cccec050fbcb799191062c0e788ad50134488d3bc6bf40334ec7d3b6e513a063863836ecfe7b514c8c69888b3757b7cbdca07baee8a0c00671011332305b5a3561e1cfd961ed56ea23fa9b1b43143c8637e855205;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77d8adcd92ab93c5940be7799e5682277ab06640107afec64e226d9f3694195835312d0c3d6c67502c24b4126f1dcc30b299265e52f3879a81a7e5c1acd0437d82bb0d45a88155941a6cd92e1ddee2c35034eb3f3b3019e36d88570bc661864a6523;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf40a61b02d2da9ca65bf405c44e8a9659d3a1c0edd20ec1e56cbdcce944376aaf5e072a42b5940e509915d9214e303acdff083749327f9df5baaccb098e7a00739de9e3c0bc60ce3724cdd3a38dccfc97960a3cf1f6fd7bf1c750ed42fab27420db3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c8eb258af149d2877c889ec97b92f06e01fc1858aeba204d9ae979ba96ab3f7ccc87800e4d29e1bdccd83b45e4751f8ee0e92d991957ebb8de840f3e29387e37932f7203437616063b5431489dda9473a34d1be608400d0e351a31aaa1a3711674c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd1f5aba40cb45b50cc3e257347ca276ac924764024dd83e155a1d8d8d019a83f2d90a08684e7adb5fa072a948c4fa78f624a86c29b48c45e6c12a3ba5e7642baf14cf4c9e9f8cf575fa99ba4531a3dbec58e7405cbe395a7ac7f11cde36a6900f04;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fd44e3362feaf4a19accfb679b04e8fe764f8179eff7b2e1e0a14185f82b1119b9c02111073f054aa5279aed64af50d5981abac1c3bf6121928ed61aea27e32518b07f8ae7b8f848e48311487161bc3aed0edc45c995b12e10f7dbdb123989b228;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37c2a9c7223528730a13dc8c0178e3f436a605f89d1902b67c60c440e20621ce468cfede34037294b994566eab437b7f902e09792d400c3cf8b9ce2e185fffeea1ded88b9f4a1a0fb3040d7e31b552a0d618fa62ab4a5f76e1e55257b8fc1c2ac589;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67a7d0f9c2348c41de91119b79c3f66de47cef0d5f85e99e6871e124147d843d30fd19a9d51390b52a482959eb93239052e708f330925ec5e4fe36cdff2e6157b2257b7156bfdbcdccc33ce6580131e47466cdb8f34cd4a1ad03dbd546e20aa26b8f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6c81614a5f6380277d759e99485679965c6f94ff75f40c9c3ae71155f922f6acd1ddbe88352b51fd522f3b38cbdb9de762534c0952dfb49a73829b80c4f79581636c2459d92f31bfc91677563938a8e5153305467d5a2c2f965987f614f44e9aa30;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c074c83909e1810d9e86fa4d8dcfa61e0f57adeb97b5a4f3b837d73826332e306900416ac7259eec0f5be6272237b1e65593f091792c2d2478b09e0f5caaa04ec8d0afdea2e555fb1295a469b7553a60f505ef3d4b79ba930236a6f1be5426ea810;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7ca5e711a8847f010685cd5e8483d88d40ecaeb570ba147ce09b4f2dcff3e86049ec7f1233ff483d115379de0462d8292e921518d12295b201054d937723569cecac4cbd8b5e2fb09b30caabc692a6798c734ae213312115ed01622283b46f03ae4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3386d9ae69bb4770d193b1f86c39ed2dd473ebca3b6427418755edd209fc0bc694b981ebe068b050e720cf923e2220fc180b7a433e34599b6eafab4a15488befe21df25a3168973fddf3da04bc7f9f9c554425cd7def6ef457d4fa5ec66dbf481042;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80baf2cd3054a2fd95e9e990e6eca205542d8b8695dce24a4812823722e3ffd710406955763d7579d92bc3f8db7bc145caa0f48859675a80342ef26a3bc6385421ec0544eb708c8987d39ac9336ac6620cbe095e06527bc67fafd3f2a53a65f2789d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2ff8b7f48e66b589b18e6bce3b74f11833a72360fb8df4c9f9d1b1c51d52127a39a10c13160baba06cb91a8139d96843e7a4af170fb43d1d829232dc431d43636e7e42f562406894ed378aa1456886248bf09494ca84ee56c61cf353c35efb8ec1d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87528a4a7050bbeb5c023552b241c169b65bde1c255c527e25d9d9f1b56a51f9dced4903f5cc358b4d878743cc8fb85421a301ffcdec520b03c7984b8a03130a10f4e352e5642bddd0ea9caf579087f2fa8449c015ba987c9c049c25587bc382ae8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4bffa8895d09f4cd34dac7f8935fab7d8607f7f70a1ff2dca647a3cd9633c1b4244ce42c922b5f2c1d6355b7c7255b9145f58d850f8b69c819ccb5c7e910b283a1720ea6441386cc2fc5a9a7476153a21802bc77a69321d31e4ddffbacb5efaeb2c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h502893c17f5b698fc5fb9b64629e675d9dff9f4a4d99f56530c227264e2922a96fedcb7daec281cc96fc102c5f6bbfe8c72ee1b05324c0a0279ef0b50b45c6393bcc04948ff900fd0fb6fbe18161da7eb8e153307d796ca667db0e97a565ba84cce7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5edcb9967f34c1234d3569ad279222761e5346f56474604a06f2b016baf6dda0338657aaec4e53712e37c19e1295419066cb3f07b7d056bc1b84e9a7e5910b82c5f6c34e13e86c67b8860524060baf3da50f0945bf7c80923b51b5f78a5d1c036e4c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e1b26913b573104e59ece8b8e5c8513a4104e483fed5d86847f5104e53faf2f70813cb39138c133bee200a53f1be163d807a7e3725bc428819faf8aecb21024b44d0d97506ecb4b76fb2d6d09a62ad402897bc653d5279a16b1949391b42437766;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb837739129e33c563510b2b05597e84fb198d3899971281f7dd30b4aa1291e51195f0a82dc8e4f3abc6a5613e522b19a9e86f52a8b1399e52f3781271159505f76bf2aedd6d67804128fc85c437ce8b836bc501a3b40138f8b3ae4c8240fa9e369e9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f451faae216c50b2ffb46821e7c42687d5f658fe58fbd0f14bb66f7dc5fa4a0cd370cfe7c42914c5b293022dbd21777ab5eeb8a9560ed1754ee62c94397912cabc72cd98bc92c3f71c41eabb800aa7d83946635f2fb5befc989c36fa2b49b775efc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa68c673d588dae0e75d345af2786c0fe2537fd8d7801cf49cbd88fc007f542ffb3aef88b8d465cde4e43154ccbe2265ede29262a783a29bf7b667a085f7833b74ed6716412806cdc313c482f9cb488d0adb61f2dbade1c90d30fb542c38bddf29d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3973efc0098e2bcfd71c50b267a0ab2747e617b1ada28f232ece6d6214a1b1585e92081e023323bcbede4bd8b6184ddc85e726487d1463337e4650688827fab309c2c908dfd8afda3c5e1869254eefbe725d5c54af56d5e36f2828551f7aa145e36;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1ff606818a3d35bbcc9d08a577d5a16a6569435aeab38897d6bdd1fabadfcc95808fbf07191443365155c3216ba9d8697b0782e71ace7905750fa036854e691a6e1a484156c1771e76b942a46658ba733a3e13754cec58d1e518b25c534163080ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he36f6e97075969b6e80a332c8e7048a933d2a5beb47d47b7669f0cb6405b43ce816c886460009015445357373becdc0e1e7f7607be9b7b4c67f666d50bce5f4fbac33db4d9fc60c392ab402bdb5d98ccad7f96285100e306c3d7608256eefb745db;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec6d3cbb5ef1bb6e8d91ccc8847862a88caa29d873228c7e4a19b80eceb18ea8e14188057836cc94208e47bffe92fe71fea37b08fdab597eb964b862fd3790be8b7eb1f3c0bd83ca589158b21a0d71ac4b493ca1be3f4ba80f1e3a1a08ccc44e03ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h563479281a0e3cddba5ad9a0f5a8e11e19ecf5863b342553b9cdd612396e3fecdff52812666d29d178499e9d658f995286c7feec1666922a1b1931ad0e50f0f8425822964533d1626effd883c7247676b022512575b22313e1db492b6ae143100824;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53e097245757e119b245ff9a69901933c04dbe8a5e224ef67e657d7b56dfeb889bfdce7eb4af6ceac8c53230a21876ca81703bd8e41c06fe7fec7c3927906c0d1df18a27929492ecce90afea96e0126a8374e61e3382d646487ffe587cc8f14b366e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2af35d14f970b44c1cf3cb6e05e65e6a5a9e5d4fd409e65429c2fe91c7bf2ae05728cc46a5cb8ef652da41ea63d21307a6d31cf13772f8c8389ee625090b604e2b2b5ca0c262492320dce11ca0e18d4822a74eb1387aa0dc8a9ecb1fdfa9fee62608;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h248d2e54eae45245980ee04d501841890dff5d08290cc49af1eb4f9f7bcef7b5eb0994ec9743b4008058e7e474cd1117639b55d7b76577aaec6bc6a05d14490f2bd779f99a56756d32ec3ec28e6244e716161dbdd6546be1646123eb46eb1a705ec2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2acbfedc265a0ff67d8bee318699f9c93e416c95db7cdff7566e2d557685422f6eb049317de09f55e0b208b33203469c46b02485e84cf76fce926321482ad2f66fb9b0afa416c003fa24f8716e84e44a58ab4f1d5e08c6daa2601e7fe838ca4557;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8241ca0f83da62f7111da03c954006d7730a951bee3000c60a9f1a1ecaac02818fbc26195a11b6f105b9f7c6c0ed8d4852f9c39afa7a2d232c93e086681331fbdded15c8ec5790fb96f3d86100cf6296b8ce35570da4e6bbcbc31475895b6d450dbb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a9626cf385af6240d7a7ff25e602cddc6cdea446207599c340bc0598739e2ef062a36680e13a1f564acbb9669ff84678b94add462c515bf82105f8bbc38f26b9e723b1e8682c840a3419dd1f2ea552b292c741c021daa41bde3b6ff6686e14804f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4337ecd972824a7d544fd97a362b92593279ce767600481281949774c0b1a621423ccbb22696f3c57d86170368c1c0c59ae259d45bae007cf85ed217ac4a093b9d3014ceb36e504427871c002ac4776e0f87e929429452f46c5842355e125076b0cb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89c2fc1f6e33e79fdec6e99437e3bca8b2566ee8b930be732bfb19d1a70741139c97d161b281c129e5a208da134b32c8643b36f409ffbb6b0ad277be014eae052006e6fd08d4992ecc8a222d92051088f02801b17f09e4951d210939da660814cb3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5fe4752832a27ee14e831b09a5ced7b689dac152b4beba191100819225ef697634568ae38ee9ab15111ff2db6fcf24793a3c356aff0a73b74a271d9dc31fd4094e90f2219fc401711ddd7ff014c82559e940ffc424e613ecbc88568e0fa687514a9a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd19aab34ba8fdaa953fba2b4d8a58742ee1ce14c209fdbabec5411b10b77dd10bea0208c438538a2961ea9fac7d6c7d72a61be33b19f235da14e3e642601ff754835c6fc3977a309908b265c3a09e14d6bce32b69b0d01b921f997e0217b3d62e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafc0e957e40a791ae7841e00062c86f9df8f47eca187d06955f74aa4e9f0f18e187a781a1f0aca5d555730c85238b0e8f42fbe2e4860770fc9adc8a40a3fa1b02c912ca82957b82fc3acf2d3ca7da12374c9ba8f8e721db09b29cffa8c0e8c27e84b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27ed5b6f2ed84b7d804137952b4f8a542e0bb7b6eca8c104e8d5ce0bbcbf3aa807e581ce9a63fbd4a9d2794fc4b31341a0aa864ad0f131b1b6d4938a57b132f64687dd705c141a6fc7f2e3f6bd800937720a6298ab7f6249bea1ce41274a4509ad29;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5111487a680dfe71ce029fefec650512dbfa5402e1e1340587552f116632dab992659294820cac7e8be97df476ca3eac255f0727e4c6adb94426b81a6fd0da515a019525633eb28854698db2f4b72652dae8c0676b9afc42dec697c56ea180914577;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h836ddbcbc8d28eb0173f7692a6fa807fb1fda2ff81f2cd28ad389b7190204923611af39d57493b733260aca8c2577e538e666edf33875d40b0d89925614f7be65a8319b833be9da902a86e3adcfe195b11799f9955cf93edb2278f38da28d3169718;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e4911be18c09214d132b2a1b24b6b506aec98d880d4cd583d3c79a0e21e85f9f5c8b23ae091dae8bc8154b9f63334962439439e2b4a1f39245c153b2dc905cf14f4e2bb305a7962f5870b3158fafc9d2dfde32daac5b94768cd252d1982531843a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7813b340849461809204a18b4038769080cc2be4b9ddce41ca62cd04316412c709c927427000797eef9c811233ee86cb9d2038741d9be91268f22a3e442114058d5cc03ac786c529e5e36ded6f76e4aac5f86638635ddbdf7dc7c1465b75ec55e0f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha491144c3358e9617324b2cebbed0a71a00e83290f3839fe605158b3adc2e9ef33a28cf4ed5f735366d327eab41cd48b1c2f663b5006ba1e3e50f785b841428d3fb6d9267fe2143a95c4878d8358bd90165d6e0fcff4e087535ea9505089b822eaf6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1745c6c566451897c8c0ad6d678cbdd8ff9d9bc0f74fc1cf85d64bb908857a9b99e990346109ff83a9f237f427a8684bfa27a0dd1acff8b84e50e515cb7da5034bcf3dd01b5d80ad264e5abf84f3a77f0f6acb7527fc422ac9d2195345ac3731e4dd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab8cccf7b5007a5caa07032bd55090e97081a137870c8973f4cca052de20bdd15d946462c12ca0bfa432b869de814507421595ba721a46b7c0ad2cbd13c1aa3a629fe441ce8feaab1ace860b4c04fc0691e898ad8bbd057faceb51d8770ea661f2ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ae8a1fd204d953c35b1203d36234827a7e90be49c8d976809ec4b248a95a6751ad31cf432197ca88015178ba1c82805b812d341fd889b2d8e528512b6a39a3a7753e44a3e8b099829ef64fc9e012b82d7ecf8b4a3f9b574e0b0b909ed90d6a91510;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29b21c80646d135d244ec81659b54baffdc166a8ce4e9e55fa96c97738fc5ec307fb096d29489821a71f3583101b27e1dd3f9ffe27100dc57ee22c01f24870bc36037a2ba722b6545f7a3b38daa23cb5b166bb191aff4453ee1574ca2e24b6abfa8c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc014af9f1a7be2dda7387a74e618de3ac2f2d561d4eb50a3a9ba78878111bbe0b94f0b00877fb938c6b2667703cb5112d053d6af7410d54102dec374e25a9595da782a2cd7ed7403517b73f65f205b1d9be46f58b0262399a90bdf6bc349b2362243;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbe9660903955dc770914e378d4ce1e977ccb32e5032a231b24fbc49e51066fbad4cd55f147ba476d4d47502afc7ae4ccb3a04493526faaa8beb16c26f7677996cef7e805bde2bb5ee3b2981c66da05a623fd81a9d558bbd89693a1e7c31193f4d50;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b94006054c157262b7259aca1b917174631ab1fa6a3b45704dff8525395873a52084b62b003a0b7eb809596241c5ea21d4a43b48dff55d9781704efe5262a563abe3db10b97e960249417437b93fa66d5c251d37d05b19d4288493fa68cba40daaf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h568b1ede4908a5d58ac9fb4d0d2016ccfc229268d9ad8d45814e5570cbbc0517f41ab19196477d2e39eb18f2e59af31cc771a2816f9d9f06050047d66c173a9ec4c3eff8c3d939891553abc2c335df1d776db19ac5325c92ece14d50a637b08c7a04;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba2cd69d36c3329a23ba72cdd7fb0a81f807eca1f297343a8b895250a7b10f8431bf3927945a1c7daf9861308637b15bdaef6163c8542acc89906e7e457099b01cb5b67ab299e6eb3904ed0f83b5b2fb4c4f7813b39f3d18bbe64fc80600635cdffd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec6c3b8d27659d38122d14866afc4ba95868f086c2f9adad0027c718a342202b67864f2c2fcafad6feb5c1928d1b856649c64743a793cdec40de5e3f1335d222c61484e85a529d691f58629d3f86ada48d2eec1e424f2aa2d9db433fc27b0b19bf87;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcea7d944924033eb9009b9c666397e896c3816705f5f6eb34ce4e02e9bf786dc4d30f10af0be0617591e526ae09f03f8c56bb889029baf768fe4359e676e0da7c603b5020a5e8ce5a3df657b0699b09b8b83a42cc95e38e4d0597d8a7482fb76face;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc403c619055c8a3bcca19a881cd1ebd95d227c2adb74d9d07d72ea5dc2c83c4e0d8be20509755085c1d0c84ff882c6ab0659c1a2ce4fa5c14089b57b7c220d3e36afab1145d720760cdb70035e88c9d574d45b05aa5302fab9e365b332f9ec855393;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf53fb1d8ac9be1979c564c6067c987e6dee9c4e2781e8057cc6269c77e8f4a8fc9a1995a1124cdebbe1a75f1779c2532239c9cb4aeae1e8e0d65cdd65fa3207d134692857bd9849079dc10eeba10cad0176efea2538446832a015b90a5e0031a9b56;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd803a5a236008791bd86a75138058112b88e22bc7472bf31d2f5837fa8faead8d82935c4e397520d51d9f968ec6441910b1d3966c0b606e3411641430798b96a7779c9eb401cf7f05641bfa98ad1a5e3acf5cba00913cc8c5dd5ab11257bbeb00d79;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h460f7d2ad284112465e1f63e4bce85d1ea8e6292c97fcb3f2afa94f94b056a25c11213b035f45e8a62538eaf133393c7750b9c1af92935c3d76c077eca1bf766009e9cd512274b0cc92a0500eacdead3690afdbb368cd6f472331d537e97f73c011d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c4160e9aef77292d224c272fd780be89b9065d9bbf6f53a612d60bc3a8504c565dd0abaade4975a26c706d7042951c2bfc6c998eb20dcd9d2120cd4734a106e774687398f75e680554f3a1c86701f73909079fae060e8bdeba768ee26ec4b24c68f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60a67fce64e9cba0c8aaa0de3ad0742705a1bd580375c67673697bb369b7bffe7ca8b660465e79c5a20fd3e7182136932cd9655dbde4716e90a97567f458784bdc5ce8e7f7247bf21f9d0e60e970067d8d985b0564a588f53c83482c2e9fa6d494d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe1b93aef877308cf119e7799b9dceb5190e4cd28dea1236d63c7ee122b1cca58f65346a117a38d1b9ce045e18702844a8419116e12654d6339d69a69a51f1e97f3b9a344fe8c72b24c53d1efdd68697f12b2964e3f5a3506760b5e318aac43b2082;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65f2ab3c46a1ce9088bd7013df08f034d1eb2aee2a4dbc7a6d4e27e48a747be404158da53da99ca27f421b755ce97d3d42044544af250c9dedb44b8f2015d0dab58509b5407ad52423ae2f28878d968f52612ad32405d33c939c04b2a90731e83cc6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2453f534e8391f8c6a99bc6906eddd49c00729707e7e23d7e603c7ca1239f886b66070e8c9a46b5127aa2a5a2b4e017fc58bd3361c291b69387ad2f291f80a34e6a16e7afd20f0789ea6d23597b4a7269a032b3c1a511fd46d846d4f962eedd0d1ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e7bf9866a54f8921ba9c9136478fc87d5d7107c1f04d179cbdc2fe7a72dcfc70292dd483f0214aef504169378ae5f70e6858788683278badcb59a4fdc6d29b54eeaa74d57abfbafacf66d0a4a55c43a5c9c341200ba2784f2a66382c1a3ee50547d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c13c7c73d528c21d5b64e9555c9d96b632ce8bdb2823a29931c58fa7608b405d87855473ce42bc3a40f4d733ff690a3d7039340d7154e47728553ab41c0273d359155d2d15260fe14d4fd3d2de913d8e69d97bbf1c7716574a4683bbf6a6cafee72;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfdd1d1269792777d53dafe29095f5ecb765908c14582269d501b39d462afd142d506ab463c9147e5e7e5a09cd30e31b54a93a4902efe252f4c6434e007c6277fc7e4aecff1fd1d2c7026cf9b252f8813c91b87c1f7a802d042ac67f51329fc6916c9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h735c8bc37a8ba0bbe7b370e893bd61a0d670a32acb3290ceb67d2cb167cabaff7ae42ad40f4632b3264a5affdc72ebc788fab498254c0f0f7e20c6304ce68ed5bf9a4437e93829229dd52cfacc655ac80b11dbc6f17fd54d817ede6b27403b64ccdb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb8eb96f4989f5472827d84c11d64489dfd7e4b183812380e14d36486bf38a244a54ca1f7ac67891f76d33d02b02eaca0cec4f427a3f3dba4d175b443eeb55d10773c25dfe9a9033db1cc69cf7edfbb3541e814a2236afd0132d0394a9f20d7a1fd3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35c1a8b528bb0f262c56329ce7f38d266306e03f6eba4e5760ac9b60e52a003165e5d0e1eaa543fc0a5c8529426872d55010217086efa4fe0816a3718044a8aa3bb5979601b92498dae5609d27e4bfc3df7cbf3abc5e6f3188de320156953ad76a53;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37d85cc5161d6945da1194b0bcca2144f42b6afcbf8a159c48e1f1beca5835186fb57d085a53cdd663ea35b6df072de03fce99116d6c6363ada3602518c62b3711076213b27785d2ddfea8a9526e644b9acbadbd9938a3b711cba827e3c27030ff31;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heaf467757558ee1a946ed311d8071be46e140cf67df22bc9476568aa6fcf02b9bb5d81899bb83f614b9d41c4e069963aaf3e3a2b13e2f639ddef99c1e44a06d687ee2f28f5bbbe284137e4388be749fe93d7a945ac525c244d50613ed77fd4f7ef2a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca136698ee7bbd20c548f50f2ed3697f3facaf98b14ad1d80acccc1a22a06a14c8a06d0a5853805b10660ee6fe8a61cb33c3b914683cf7c41bc1d1b218e862631229eca7e796f9a007a092a30ecd082c16113203d55fc400e9f3a92e3a131cdc49d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf623239325f999250cf9c194515c9aab660cb51ce5d920b254ed320d8e5b4068b8367fe65bd940ec132ce5365c7aa512b88c4d95163b8d1ad869d911ab345aea4e8d5e58e2d81154fe42d04cacc74471e58673c0a3818431566b1f4a3461ce04454a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ced0874996e4118651561cf865b31124ad3fa5e7724899018e3d6d37c4a3f40e68a87a3b9add711a1b3fe687cfa66d010c802c0558ac0dade66da8a89f3c23d261b189d2fe31babf8a98f82acffab44cf1231eea721d7b269ac3bd1b23605be7693;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ab858682779deef382e7851afa527b0e0c492c4d8f9a822e43b1da37ca00891888349102a4bcab6bca3e8295f78f757833f8d0a95e287e07e76c146006a21f3a6ce70d10bdb1036b976eef3579e5ba034e354a1ba09e0aec2c0343c534be073b8f5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bcedb0fd838d8adebdaea6f276015f891133eac2db847963cd484c0500b097b7de57ed4571aa93b7c8420cf90b05fca91a6251201e6113385b25a62fdfc004be885d0ea47e5ed371a21c023ee6a93e289e4a31a0fdb05ca791a30e98256e377c09c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77773e1e352a5ade5c8edbad9a69b45403b23d9bc46b778c402a651649b54778ec5ffcf84f6f4d73c6bd2716d8fd001d4b46c8beb2d70b65ae5251cc9a479f1e26685e262bfefda4cc93b195b5a2785778c82399f3106ff3aa48e9a8d668d8fa844a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd06b56d406458d32fe6949db9e4a59ea4583b4e3b09b9bab48954841854e720667b542308f3d1deeaa14defaacca313d7c33cbed0ce0f19e29ea9f60a3c784f3f0c447a272d0cc2a2f7271de31ee72bd3acae85f365d7835542d9a9b2592d17313d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf593fe8b511a10bb9a7c373e9765788475cff08a82d4a8e9153e077bbb026b75df24f61da988bed83024cc8f0d53ae023fa2540ce0815ef750b9c3b627de766877db0414a28ee32eabe2c7a78e80ae17c30133b337c45a37b4b2a4aec8c7c67178c3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66c375dc8cbab6a4a1e4b9a5161f8f7b2e7135b9e352e31a3e0a3c4e8f9d1149ec81e378991c12b6172e8dff4d6792a4132547a51d6f6ece44fee666777f05eb2963383c3d21f509d4a2542a8460dbdb6bbd0bdae0513219ed5ada92fcd0b586d87a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he02430c578940b82cb6600c125fafb1485f39a204ed24bc3b110294213354e6be4e40b61a0d679b29c27d4bbe93e66480717156cc332c2f4ac0ea1230e89b9424e2eb60ba7573560429f9354c72d39eb4fa2ee02b11e90278d3087e1d6fff87fe3dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc9520b6240972359e23d6b45c3fa3eb78ac59eaa9d5b66481fac6716154dc9e7172b437dc8848b66d08a0b1f8d3113bac7aadb620fe3e1dfaa16921586d806a1036ea0070129d752fc6f8d972f7b7612281814bbc33b8e7c101c03aad3ff5d5f1f5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fe4b3cc2c0335035be56180d949130003e5466031ca01a39f1273c950438ae76c36156f348b7e573b05af6eb82c274cab0ed16a40bb00a98c52516a9d5e616473db4868d35150c27025a96b9f8bc293811135934cb55b87fbe801778db5a59edcf6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h975632443973d34e9165d39dfec7b7b32e39e858af9cea835c566e8e783d5f247c5c6ef3ecca3aef3b8cc51ca3033ee0775669c8f3f2ead65ca88cd339434514b107373b67649e532b072184920e2c142b0f37b0a7f30f0a8788b2aa02d03b78d54a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0bbe108486860a1acd74261c8c1b61a050421f2fff6825e498c00d2ea1105443b2c6c38fb7dbae0765581e8ac9dd1e6a019dfbc47e01a44c285e5c83de318896e83b96bab4f0e1a6b16365a6e9b58ca7090045982af7231286ab14366ba22b142d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h214f2d080b45606a916eee55db936cf4c5263c4e216d58dae6f14022acd73af06bb9cb9c1f8f1107c07650e4ea7f549a758f22f940ad15b9d1551735f418661ab27ca778a30f9b2dfdfc1de09d9b5fb8cbc8bc7be90c50711fce4b1a1031621bd278;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b24bbb10d845e94f55ff72c2488a5557fefd4d09411c7e7cc1aae4ed6665d49128e520b0121411b7434a9d35726ad4e1d72b810066354e59f25954f44940e1a27b55b54217b9ba95b6116ba109c95ffef0a3ab0fe5f9ab9601c7b3e4c1c79471d9f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9efe8e4e298931c9026f64f2c39cf1f47a955f7407c14fe3e1bd14e395b41c68ef6633f7cccb6c1c2f51fd4175feeefd1b4c542676814b512b66b3aef16dae4ee87841744cfc14e2a3cf20ee4a90dd1dbfef4ff72c318db33d0b217b2892a282eca6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb52726099a7fda3177dbd55fd5047f956367f53450d681e9bc3a3ef4b13f361f0b2dc0d6b34af0fd79bd6bb31bf8ecc33fa11a43dfced61c7a72e946c1e44934a3c8a34d0e3aff444ef56b37bec513d2eb29d84256ad5d81aa80a90f6ebcb0f2614c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30adafa1ec9f544d510780a5c681c4fe701880900f365201f4c08600758b287223941e0a3f69be7be848531ddfd0a2d4e9259b1bab06a79f27723a6c9567033dd76742dc2f35179c5802413e6fb032a64a6089f083c4c3b42ccf431b1ba51998b757;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b45c7b8cc978b5bc218b5ef7c26789e7e4346434e32699c31d3337c3e8e56799ece75b8ad05701e8dcba2884bac96dc49fe6ed615ebdc01bc51cdc6f325f3bc265d3ff3073f3f809d41cb4f9242df6c756714a73e56d8678b63aea133be497a53a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd41672ed37b9afc53b6d82ec84314cb8eab23e147308adb51322800d078453147726be8f73bd2cdcb4b6105ae186bef147ca9fc899e7bf9f61f49306a581f9a3a2383a02f36de5a08a736024a3b3564a9e551ce3def0c7dd318282c2a94bcf8a2b0b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca4e845689f4d5c5f12fb8a843e055869fe4ce4c9a943a1fc44cac7711e991b8a733b52531dcf4b4eba52bf402fb2a56c9889a2ef44003e68b45e8f5aa507fd2e9d081f5fef5b50b8232ccef93df8537eb0ffac37c5642ff185d77044ed3ab9e7a47;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e6e429670d0e2518f6ced705fce5f49ba850495f2ea3173d4fb4133da8cd7e0ae13fd27fc0eecdaf8303e584e5d5e8d3b942e1507bf9e11d9287498fad7e81b374151b5c4b92edc946bdb5fc0b47a40e53facad3f1a1c278367eb34dacec3e9f6c2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h935eea5488934c730d0708d7121688d05c4ec9a768279e663624b00176be0ba4f18c8ac324b37831917703208208f2ddac3187a3a8a3e4cadc9636569fcc052bed7a3db886e5c406d829f59d2ee7c6e891ee31eb597921ddc0c8ee0cbf71ceec7516;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h580767db3c4b00206b8b818a3802e921fd829cb5fb0afc6a8fbdeb1cdb40c7218fea1eb5ab28b30e5ebb058345c5676280cc72fc5024dd1a060c9948a34864df2d2b5f4031652eeca32c6bf60c3a0164868ce64415cd620dae6652f2d30936f2876e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21bf076de20629819925a4dfcc7e83ddfd294734158f09cd4319d83c18f349ac6e05ab0579b2eb893851ae911fe67f4f4794e1695619ba98f55d1876addff7ebd30c193024a8d785b7777b9ebe968a60be37a445945286a9b63efb13e05657c43d90;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd13922d3b56d228e8323c387be10cad5afcb913896a6e18856892934a8c47307710202defecbc04d95c2a1dd81c69ab03522a439b4e9b91fce69b47061c10bf322cf121b470c956530bb07d0b326c2b9c59635a42a9a46ea24286d238d0c7ffab98e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcf6bfb7b5ef23053b042072899a1a16e92ffbd7e4ae214bf694bbad14f321ba59b5a72464d31dae8f75e53502bf139233d0508498b264e019104f3fba6580ab457dbb606ae2be4f9ddaf1a104464da534dbd6a2a37ea8ca5343e12fa1c89f3397d2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1e8365a7881ed632200282bd0ec429329ada66097f0fba9071d4826283f161401de9d92d7620c89e1ed4d1aadec23e882b58db580d8e51fa6c3f6bd70df5f71b1ca9a4a91cdcdc0b2a7f0245266fdc5c165f71d0d7243732de85e0409c11b7877ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfd5b08d390dcc0c21b92d76fb954257484518f80c084027f2e326e5507529aab433a4d08390ce3638081f3af2709969e7337677d8fc101ed2e533957b81b2a2bdaa1511089fcbbb873c7efff3d4fb50291bf8a1b50b11fc9ec43bcc5fbc3cf9d844;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd57fc8228b7c38a8ef42fe070a4b011da5bbaf0f054b7c9c7ec968fe20d536c173bc265ba92d929d22a3fd45003cb467c46c14796a502cc13d0cd405d292c30dee0c019b6bef5ff23d7f47768b99dd339aac6b2e1f1c5359a0ecfd391cff2c285fd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h681361c2fa751dbe1224cd36569813671bf2c4e02d005edf36350a848c1155b7f6924626dc7faf21e96dde656f484e4ab082de30d455d54fe9f45491cc99fed373ca7a6d2bc02f23b4f65ff03f8a8c6daff0a8cba0397b4e601e55ff5e8f8d88e34d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25e4841a6381cbc0358a8282e4fee84f96cedfb33364f22c3029edd74441481ee2ee461ec3f37fc59361588d904edeacc1fa0a1e00ff928762d88d62c9dcd2b43e51fbc5d3875b0f7063e4a2e0a34d7c5e95fbf473f2507d86df8f58e2155fe9465c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab78db9707cc53f1d9e1b74ad8882a05413538eb3a1115a248608c0b5544b5b12f83e3cd59d521fc23bd2acd78fa86ef2854eb5cf7ecf9179c9b6c551aaa703fca9b7a9a957e24cca1ba04969b98181999c925f3a04a8a9b60f2ffe1099863180607;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0c673c8b1fda5c019c8b77cce4a43081877b12d996bd6caec9b8e8bc31ddd0515fb9bedf56d3bd98c145dbf780b3a9cd4a48ea3445ff106534b814d23fe6ff17b35c25b1e5497450e10d7e06d8fc222602a26c4f354dfabff71ffae66cf676c08e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a4818e05b2c7140f9fdbc4e9c653f85b5a6dcb307be5f99ee9ca7e72741bb7a08f64553ea8179badbe80789bb9ee7af2fc43347161ec8d039a3b55ac0d44b227375ad4ea7e70b004827ba46735b4c75f8e74807d32b817ed5c8eead9accdc95d37;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6ede90862e1f580b91b777ecd794ab6e7a155b5cfe519b8882bbb52905f6c73df0110eeed296dc9a621c682e20e1b0544498cc2a6f23b0e885aa7a0c04dff97d7e34cb540a2a7cd586a326ff1a4be3697c275cd6174fd7b83cc0c3c5bede67b3204;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc94338d4a266b32c6e1ede8be06c4c2b07278c4f2f51d62990dfc2b9ddd78e37b5bcd0e2ba914a18cc01f8e62dcefa389a9d67477689f3fb9878417be8c48b17fdf6a2129327225a84764f741fc979fb0399ae2864e7505eeec3bc31de6a12383662;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h893b72a39721f36ee6f5396c000465d1b59e980f984e2f51bd115c2702aef1ae34214252a7fa4ec1e73923d808c59f9c44a20d1a42d054aa165c97c5ea0ad0421a95e3fd32301b09014fe6eebfe74b4cd1980bdd0cdeaec1f9753cb217646ee76888;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h533df3defac414a9c9d45524b68ec6e48d222d04b51b52560c451cf5ea0e6f5c84d87a63dc284e8108b51f7f2f9d64006c84c8ca0591fde0d06facf3727ab7c0389d8340b493a13ee97de91abd7452e4b936efbf59506f6b31e44fecd0e19a50cddd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2938d784a3d025e736f3c537aeccd5262e44fe970ef2f360963eef7c7a3ba5e6959098358e0a6c9fa0f4f169ab9ac59a95d372beb3b1724f49b18913544daac25980076d18e927a04e9694ccc5c46f7f20f2bdf0652ad3f4e1f76b995516d3f209f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51778db445527616a1f6a3e2a676455f35bf13f1c9f0dfe1e7ca82a596da667b0db4cce1a50ed8d5a902ac4e8019deedb0c1f711a8136d15c381008fcba11db04497f1c40a8370249e159312ad82cc562945c0113c1cf9ca660c285ae52478373931;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h421d1cb3c69f386fa79dbcef4077b5b569574b2800096935b6a1cccba1dd44e6eab50136cdfaef3efab3e385b00ed6741974d88290c42ffa578bf5ac64f6c76e4ec254d28e55d198135da2f6148d28f500874b3de3b8e8cbe091a660e2485a7dde20;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f6ec4928c47c03dab9382cb17073962b205492c29a874cf56accad7621957b1f2412dc3ced44cdc571c5eb935ab54eb1acfeb3421ab0eddd7be827bd0fb37e40b3ced168dfa3322771f357c856acbfd108998eb81a5ff30f8c876b474fdfe66b837;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha7b25c6bdda334d5c1957ed4eafdd0e5c9a4feff75c32c19820103b48bf731206a4b835774550edaba519b0b45f8d73992aa625e0245bcf42415a4b55f0fc3a98e1af3f0151c75b8daa4adf6a4157af95ceabcbe5fe5b46bf230b72f4072ffa19b6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ba3dbef9a85c3fdffbb3847735aac94be5efbcdb94d31f1704a5b23f3e1ecf23c5599e1e981dad0f2f00ba41258fb29ffa62904ee372d2b31be1c323d2ce2d50637eec256e91eefcf49e2d3f18e5713f7172e412b2e4067f6610112a154048b8034;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83831da0bf0c3e49b9cb8864edcb6968449dc79de4cff50ddb1138d2f569c787ea10b736a8769ed92f915a8b2a90735215641714868ddcd84671ee9b0188418ccd0beaea931f70b72b4f70b99c925304a9ac94501636304a08a12f46dae8577656ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32034f129d482d51a0d33f6c5cdc666ab920e82839952c01677fa4d0e6dd615bd56b4ec22b7ff743b5b78cdea58e0107ef39f342fec033c5089e3b0ac7f0f47f72a00e3b76fce4c23a4c399f01333d660d92becfda62b8eceb40625c8e67ca4a6938;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6bef10d16705bd64e22cacd01392abb872aaa813b4fae51065549eaae6e05c11354ec9234f442b0cfb1e2039ffa6467622bdd625f03abb16b0e5e914d33bd929a89f8182709a08886710196df7e43cbe8c6ea2a9d6f27988880af5ec75ad228ad4a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb450aecb2b67e5c7a011423f6ee30bdd48f379b314fcf414727d7bf93b820a0269f11b946a04b5df9ed00375509e4b5d92e2fe38108d4e4ffb5cbb51bc6ead0d912e462dcd988f28f67ad210d74c8390019cfcd50930401fe7605fa890633b22183;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc276f33f72ff0b8846b4aa827ecbbeae7ef0127ca04d7b90e0106edcdbd09de03f7346c47dc650d685e9ff66f47a44c229c9f982ce9cbd4f381ff610859bf07f7724427f8774acc94d339916ccbe3fce9363454e8bb28a5fe9a090c57dd3eb318700;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59cdf705fcd378cace7a18aebbc3efa2a1c980c1d498fbe01d64a5654f8705985c99b921aabb4aed8eb0a5781941388ee5c7617c6ae8057ad7d5870fa0f63fd6cf0117121c47f02bdfa2e8aa21ed3d7ed885d0932ad51de951573d8164288ec2bcf8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb46dab363984912080384b0dad1eb385cf4021aaf1aa384b86e874955f41260729d79bca12c649c0f665a6409bdeb073bd8f2e05e2d52abb5fd3332288018c330eb77ea5d69f61ff91dc31325b3ffea139971927ce737558a41eab9f43c759ee3d76;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3558f207705256224e495db127adc8a5e7b12e7509018c968039b016d087196516adbe706080f1449bb5b13f86246b4d0bc985b5725d6155044e85fa38ed32319f28a9c9cb6a415552f40c1a3761a21bac14dfc108a741ea344ce84dab91e34ab2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f77daab0a0920a841ce4820da01d1f43afb0b657ebe474c769ae709a68ba05091a3306fb8121b6dbe7f7dc0ceb2d34747acd6c7e9865ff2123789fec826584bc80cdf12bdd15ac269460559d37e02db81c378a948b070ef5eb95d588d372d9282bf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1aeff4ace73e5db9027ce853825831a091facc7beb408867ea003bc861c1c7c7352b394410cfd0de76f14c37c1e66a0c5618399f6dba72dd0cf2f9a5a7b81a4452de7dad6b53ca326fdf842ece31c50fd0211491680a2627c593cb86f890a5fd8fae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h131f0dc1dac112bed283991eb6f7073a15336a535a65ea26baa3e845617e68dc1e7bd704653b43da397a713068ee5dcee0411fab263fc2c8dd20e42563f32c1f606fce5fa96cbe979337e289bb7b790e4b218a0fb8e3d82167f3c9330e6012bacb0c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84d174ca3cfc8f42751615cf87d0ec916d1ebd83ecd4eb719cf0aaafd6a41b4677020eac495e8003a26f19e27d565b690b4369cac76635ad9ceae1392edfef8f97a61a8a2d2b138a5f19e900f63ecca6457ca6d3cc452715edfb7a858c9b8545b3de;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h129eb02594ff3b1f230034ce39db9f751a34590164f5ea11c9989ab6449cbedb3b28dcb0b9148e5ee8c8b1326650aabfef2055348de48855f193fa1cb2412a1ad14983ba9178331380528df245aa7d265747bc7df73bdea75a362a9d2e4bed1601df;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fe8ac50389f2a513b91128f5d06090094da0e5f91858d5be9ecca4b3e7c0a3ac9c1538b1c262c4f7005d98c1640df33df76b28dd6601e3051e04323e7f85a211b8e4f7d568f189421e0d9502551b31ff2e7b0aed6aae9092e24a2f0918dcb123c94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha027e337bc8e2a32f18f33ea1e673e437de222557d80abdfefcfed0cfc95977c3c5d3b05348f72bbe46e27cfc55d5e75c354139c9dd1e24d639739eb0808631173169684c4e139378cfb8184dd827c3a66de805d5bcec49b8ba2e2d90ed87d9c00ac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19713c65d766780dee50879b29ed24b419a36fd9fcd51def959c951fc1ed97a4141d754c29e0568873cf992c40e32a6b3d7077c70f78af2a3e395f7d53ed54a8eeabd00c38244d290f97cdab413ecc3bda802b1230e3ec104c2217da685e93d1c730;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3a869f18a3e131bc1ff0be382675f0b48771c771d21d48e931383c2e2109d3af2390e54c539ca6541983494c3f9a33fd8181ccb81694d74d6941a1b74054957fd304b4b5a70c3fd07d337bfc0a4d4098b415dcf8316b63dc25391c585fa66d3a857;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heefdf6f566f40bce4978a1a9a445e9b463ec9bc06f828b6fc2abed33b68dbf014628566d965cf5b7d4a39e202d5c6846e683210d60392658f8d56e10fd8fa586e405677f99b80ce4c8157adc23b9bc3e50f5341eee7b62ae931294cf54f169f25787;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14964f5f7ee1806ec000b538b87a68e048fca7a679d8a8c0f84f61f4d7a7820abc109a07df319586e0e34ee22903c207c0829b55dd6815dc0bd1f656c5de90840d0cb7aeca8ebf47f6ef29c9b08adc3426b747c06296a2bbfe450f4dd461160ed56d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4dac28955e70a5cc4573945fa0536b05315b4bc698276d3aa26d2f278776e00eb6975f602eaf7ae8bc6530fe3a744f56febb9574330d18b4791cef7c6acdb2faaf949bcfc3a7adf2a88436f0c635c728a8de82f84d9e3d6f249c000e3f15922e0af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h994ff4b87ba32d7c670e38ba986ee663a5a870b04ffd4ea6cc13605bf8b374035b853bee4f797b741f0eb31de15ad43e5629b44ff7ddc2c6adbdb62df4e49a26f25c54a36ba51d76b4beb2a3c8aa5158ad617b3854e373813ecb54bcb50a22182594;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6a1f977b4d7da8d78dfea8d16f6feb5cf936551587fb3b59712468d3c52ab79244714f319e0d3a277630c6240d382ef7d0cd235a16b235e86ddcd91c1df18c0e727ee194aff56ceb0a89850415b91ebf2d418acb4bcf41f122d13cea487963e2b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ecee7a069b8bf18beeb4ec9cf6cbb98267dc8e9a511d1e1eae0c0dd60ef0a0094b380053be43738beecfc4988e8b1424c2c4f698f2dc2359fe88e8fb6c6e07d80461f0ad8ff8fdcf6ad3f84c5375466c1da1e4e8ebba4f15c79fbf41746db54f56e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66731420e33deb7f36c5f8943950cfacd98be6c0313ffc163c664e905e89f600c84908b94aaefb925129bdd0b8552cb158c4ce5fdee714015dccdaafce6c0251b3c738a986b7f6a84ab40411df9c47cf4c7d3b0be96ea2f263a14fe47616a0c0c4c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a4bc5357ba684a6dfcfbaf59c979b5deb073c84cdf01a9b8697d953c3cc7349a18f595513d988a6eec0e0a67cb2d6916d8e46bc3d87a9a05dba91a4cbb9ea1d012751f6879c161955df3eafad847dd7de9580a886e4b3cff12f66abf870afcdf3ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4efe7ebc9607f5591eb466de4bbd4a7a6a1f39aa51a4cdb1be91f91ae5a4400d15d693a3687008a72758b4ec60c8dd8311e3c60cf33dea13b75e707f53ec44e7d21d0e898c1763ab56c0c1e5b12f0a9d8c89458c5880240b362a4f97e82bf5a2b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52e2ea38122afafb29b5ed8b73bdbdd21d4b100abd8194c88f16693444e74fcbd457365ccae3dd2a0dff9b6efdeb76105d704b2f0e2b77d2039ccfd1de79692ed95f238d1ca8bdc98a43de2fc195b14c4f06b7af2c715e8433a3858d826fb281faa5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17d8902f3b319e53db8d48683bfb2091dc8ca4b9494ed9d78a8958051d4987189e66d723fe5fcfd4a592a48484c2a07f6c4e8088b8ba16736dfa64c6053e9adae0986a350517612344dd1bfc7d0186d891df833ed169838d9cbe6de78dd0215ae74d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee58856b51319728fb6bb9a9f49c7b6f7e91227eab3c781db5655d5f439836bef29c15cd0824113e6211d6161f1a94784f77fc7156624c8110406851f77cde47654d2ace59b657c4c97d06035d62710d50568d8f0e833748da711053b2964b3f7141;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf642f6f2f5ab02a5abdde883f5191e2ddc2fa5f8cc20c3e4ba7744e194aaa945b9a0ffc7221a9a7ebc87939f42996392b6f6c4e18c86785fc81c466775953624ba3d3b5a157801409a0b4e78ecc8d2afeea8c696461a40bb27927a7a927f873c69aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he23fcf37442139d3e43771d6b94796d0d83cc55ee01b4c3f8ec37625f37ccc94b171ad3092e87177618f1d26762126fa90140a575a303a365dcea441da2be02f9ee4143e56027ded63ce670b4e38656d1ef2ee6af9e65004ff33159ff62c797b8860;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30d13da21adbb5f5151ea97200663e6438439631d11cc4b016cca6d888301fd4362738fd006a1271935f5fcc51ff88ed817ef59251f3207b875bc569a5474345502e13bb2b45f777d4d56c6726bea819540ecff49968e0c94b406ec1bd74ac81d75;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9544cabdd02999d1e98b3a8eedfdfecfbd2546c5b412577fa1770bb8a69b9034d484b8a697b747484ce7131ad81952c3b48a594600d2356896c35212df5d03ba6aed2afe020296f847e4db8b1867280a5e1c17e0666edb9d5425eb2ab42140df4de1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c2e748dfa730e8ede03e5d7eb46a8145c15518bbb8075e8c3b30bcf80cdc64fcca7260daa093e5e7599e641f272ded9df8e92635a498a73ab07d53683a7e2505ba4c349a149fc256a6d7d84728b2cd99dfb66ee388113510468ded9918e8cfeffaa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9bc4307f227a2e68a92dfa4403f5ca6f5f13cee713f6655f12752c6456068283f2131e17ad2403a23ddcd23af017c284f1cac50628f3b817b62c76c65d713ad519123f139306191501da765774ec7acb66d73958b85209b56cb29a1acf11464da664;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeb58ae6d8430e0386a114b75c49a57eedb860cd6afcb4f901679c3f27b6eb313511d5a5223a19c7e45366ec2eca4414e5fae0071e3d2d19f6fd94db54076296be7953f5bef608c00ef13e671fcd189b37c8befbc1f487cab22550014d203d697065;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9815bc9f46f26061862c2f4f7a3b778b5e4744a9bf00d70b9c93753db768b3061d3f76c68f5abd5bc6adaf0abab7f253d2fe791a983e3dd2a1b57824f26f60ef2c797584bd4a7ed4ae65d02f28339c647e8b7e8a65c0d9547007183fcda28b680f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfeec1575c6355af76d23880646043d40bf7dac2e72daf884b6983c85cb11a751ff17cf89df9542491c995bd95d1503ac1eb08de9a5f7a12624f691cbba3a172e414d369109dbaad5445a324ef2cc72b3ccf7a6945cfc597326c45910352eddc8a87d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf31a8981db7b8b972df42350f9762277667ae06581eac71ccfebe3430f611e22a42dd67839177fa5f9a9b9c119bba9a37e91144532d165753e4669291f03db25fc077a8fb549a5e27e727c5704cb6dea91f9537a4e3633843aef1bb2849d5fa3486;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd48a50a8661227f85bd34baf8679a2944e624372e397928f756cfb1a58af87c6da6e266ddd1afdd9abb9a7e322c6ba4a1d5278fa7887a2048df38747d4fde70bcbe052f9431d9a75eefafd7c01396308f540fc45992a85e7b2a9b4a835f0934262b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5932cfad0b81f59c89411d105bc0ba52e119e721d351036f762db270062e359c59c2c34dbeabe4956266a514aabc874b2bc6eac4bc9059116ce5ddfea6ac0ed0b1ceec26d3fb808a15ca5b592e70589a63228b222560c04cd60aa3c280b86cb536a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd7cd133e0841489079b72430ef09292c3c233bc5191a225ef443e72a8d431eb2b6b1edc3ce9fa145c9271985a34f94c65b34c98e75ff2be752b65e0116c9b228e10cc37b081635eb2ddf2210630ebd4d234f5c0f7e15103535b62ecf579ed99e20b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd31da6206173ffd9ccd3a06055aaa93c8f1fe9bde8bad693f4a48f566bc9df286b6cbecf5e69b081d14f7fa7da3394121542d394ca8ac31429433660c2abcabae9f7802d0a56a79c68fa9964c8ab04d7b28513f737828d1adf4339ba346bb34db873;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2739347bd01db46935aeb85d4a26645e3b50a3367ead0337f7eb009d94b7deaf6351c83829ea54725d17ba89e3bdefce65b88c9b8b99d93ed3345a62228ea0e5af1fb1c40a2608d06d30c27b70b228b4547771e19b0bcab8e0f3e794ceb237f8dbb0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1319a354ec8eb017cfb268535725e2aa488c4377ffb6b88a458f9e52069d027b24f98c89b90dc8d38bbab905cc6c8fe565dfeb03e32bef82718670a15ff2e37d8d3a9b8da8f97f31c219f7556339c34f25787a6af8a78d4f01b4ed88e250a9972818;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1f0ec8ed8b506ec77a848fdbad4a7b8b70b4e27375f907c02348e8ae58f20c5acc4121c42bbc15b26f4b40fd8157b4a757e108895a1df53b2788bf8ee3dfd259dfca5eefcb9ec18809334ba82fdaadbd786842fbcc702a440d590258fcf815c23b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3e90864add7c154f77b635ee31a82544c4d86f94a67b069e459deae8f99f4dbfc1e48a6edda4ec335ea5e7621914ae8cac4d242dd96bfe10f6e4631520515bd221c289f9a91f5e23ff996b2ee1eeb1f16de438dec9c92539e07784dd53852398a36;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8abde9476bb7b730d6752850a0911d67a2e694f69aced7541966044fb814709ae177b4c88bd6083e014e04673942a3fd70998cad7741ebd085a1a8fba61d7ccf4f85945c216fbe72b457fa87f185f8f89a9c5d3c8b2fe5a56240346708bb47effbe8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6b85eaa5fcdc37d6331b0ca9698abd212fdba1badd45da77aa6c12e4447582e99f84649b589ca3c4eb4bb04bdc6ffd6b1c7a8d980f6e109a31ea6369d4be638a29b5fbc22978be73326f006d030ba16f509fad58dd3d70592a4f298d23a06b81e39;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ab5f7b830ad305295e67a4cc3f194c9ccd4614abdf57cdcd4802c728c96faa45b2f98759f45a0db8e5e6a10ef73a9d923abba3bb387fcfdd2255e88c698e7908a66df63e76eadb3bd290bcc8c6f6c872c558bb6eddca2fe9ce7a054cc6f19699df9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c4bbec9ace50b911be6f2c35de9e0694c1c03360f1d6abba558dad76f51be787c12f0e057c6b5a464c6f99f35d1499188757a3a2bdabd24897a26ca46b0864870f07c66fc96730b134c526155d1e1bc917d8154ba3cd3c7b8ee2b7a303a9ae724ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cb1520bc71f0d64d0624b5b3b2cc1e8224635d8c0963bc8c111990fee7c7e25d632acb5ce49e33b15bfe1392fd2ee35459e31f3b16d973e73db8171f08a6fbb682efc740a656b9fe58c832d7eb551f344c43cb925c06dc1b380a3b3b8d25fb5330e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb4f5988e49463070b3ad6e20f836619e584e72648c43dcddf22d0873b10a5909a387e57549e795d5d93498e6334862b500bcc4d8afed4a9d4b6b997763a692f61181f93cafc307ca0b60162c250322e64a20447777acdee2505e92168fc39162145;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94d7468620ed70ee640c3ce92cb646c48cd386fd89071cf5817fdb4bc41b6d1c31a6585a1eef9748effae130a48524be7c6b74872e966427d16ad181c478834e86fe90fd6fa5672c2e9c9c485492ae821d92901c28c3a08f446fccee4690a5404bad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a4f306451dfedd13771a0d1bd8e2444a3355a5a009ef282ee5ec754fb269fe7977f41f2fdcbb2766513d053969582c9e194b0a9510b20133bb7649fbaea8a57d24ffdee13db6ca18faefce40fc9b46182dcfe086e2277b533a6efcb76ea7260b496;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4b90c32c0e0fb85cb9336c702628fcce30bf0a3dd7996c91464392b6734a7442e0a97e49c448ac32f86cd4b2d975ed8e571d675ee382f592f0839a4ee063878014bdd591b4b3caa6812d318bd6f76c3e067e83dfbd038ecc8fbd24eca12dbcda5c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf00b34b8d744694b87567063a953032a56fff3636e8d98f0e5d02db396bca6f7d1fb593eb1808cf098084edfd6cd587fcca111e5096b6c4bf6a6791c65f403187a76221dc5adfea92152dbce7c8bb70649ebe84315e31bc868c98f3be8052ba487a4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88519061b3bb0bf16d15f0c0e5956f6db5120f71c4ef46683a6ee288627c28b1056882523db31be6c038a1379f960d48be59f98910f26eca434db34d2c9f3e51c7d4426cbc8f8a28c85ab513d2f6fb9eb31e7a1185cce2fdc7ac184d77aabc6f45f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4043f7c273585798963161035e6e7d4f375a5f22f537b64daf6d51097d47e43fb40045f53a14423fca44f955fc6afd1cfac10d166c8e41b6c268f0744091c85d8db4b517674b8d8377917b6437075c65abb2662744306a8ff7f59c5af9830928c4e9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc6f8de9802d5e2ce26b14c6593134277a69026eed6efdb71df79a07eef122f858c5778eeced4b61f18e4c988e1bd30f2a4b166eb31735449b8bc2f7acb0e69e5a7236c24d06c6cffd5827e7bcb9a83efe7946d64f0daca2fa91e2242cf23161c14e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3170ba000046ee3856e04133cf9024d517255324130ab795fb272c0b54d0a8a0f00e1db3a643cd0518e60b648c5101dc0889b3462dbbb80fd733c7ba434571f2b2c950dce500d779f5b6ddba8dc287c33385595ae01b9444e8369154d1e0cad1d774;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6d4e0d8815621f7a6419294eefa56b771c972e978fc5edcbbfa953b03f69f2366ad2928c777c32d09d8e0e6d6e07ed8c439862853961b0121049db5b89b9f0f84e3c087b4d5d485c76deeec1fdb75681e3d60784ef7d357d806911126e183a9ed3f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9a94072c660e54f127c7df1a118b5dc7b2222f222e46227cbd851cf50cff8a5b5bd2e755fd56032f3625ff2c14ab8a097a7a825238aa8540a1313bb8b33208d058514979e17a1be4a94c2d17efaf7908a1ac1188b7afb049c11c0490b734a4b42a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe88dae09934935b0c3c39f3f0a7fc2ef9ba947f85fba9990377044f6d65e84ebe1655bf19ca3caca8c1748ebb83fe4038dc8422613c2c4cea6afdcd9dd8e2ab08580333975f5aec6e389aea9abc9de5ce37ed6d976694f92c2f1863eb5a512f8c03;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcae8665359bd77cd0aeb4f54ffcddae4de950324f0ef3b2e2d162aca710ace3883ff7a2a793127fa9c68049804a9f034fdedce3d36985495877004fa8be66ccf88356c43115d20f42bc8b24af534bdf7e869544ca04f1b1b3a09b661917fc72ce4a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92d24c6e01e72c0230ca4d28c71cb4d4ec926b899f2ceeab71f4516b38343e124ef4a83012d0981fce7607c7ff7a4dc28cbac541681c9a01631d133b94f3f8e97191bffc5bcfcdc35e82e4d1e57b39047463410ac1e18dfa676d15d88a96e8e3429;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h241d9e50f95dfad574cf7cd3a8f915421415ece170a3cdd4f992a2e665df02bad4e5226e1005b77e25595869debfd9e41c2a2b8ff99a8ef3c8064e07357f3875ebec42418a5009f8fba23fdd8f50015b0de4c66fe06b31130a993f8ef4886e7c0531;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1041383928a5f61f35c60132963dbcfa2cc1a733928a3849fffc6a3e372f98c7d1fe47b174bcf63139dc173014aa3b8827306e27f1005a5f40a2d1f140fdaab7aa429cbe046c0592da785eba96264578826daec26a488e4cda0758dc6c79894c42f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b929e7d148652ea5c7cf3231128d0fb5ce1647ecf618023775c1bdfe6dfaea814516644cb25e6e33a4e64a37308909f6ef7c9b826f53cc9c7b0852971a57c7c31a2df10efa82876732ca7f76b10b90379b1e31563a01e2cddc70a8542dc874b7d7b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec6958a2fdcb555172feadf78c30691776558da37aeaeb7af40e25094ecd368ccfde7a0acd17b9aaaac447a0b572f5cf3fbdc33d7489bb1737f0207393ac6f0f9aa899b53039f47aeb3be20b0301b3254e0f2f5c3702f90141b3cc401ad4e54e2a8d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8361bba34fb9d48392d0e603b0d6ff45d598857e879e98fc0d73d57aeaea727623dcf265f2f311f49c584b27e9f2946dc073aa024deb7a8141b85412b37bbeb67991f10bcb7c70c8875fe394e3f45925e7e35de66591b34c11cde7631c1e4fa640ec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h299951ff2c528de76068f03c1a0ca93476434cee1df36778801e09e02c1dc7d4fc346d4621f61c8c39326396af322176cb26b7e23b4179be5efb5555c1997893e55b4f96666b1045e35c9b5528daa10cff684f50503d80335c3f98dd4ccde3b082a3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc39ebdd38ee35e7eacb3d9a0a3d226b15fc14861009e00ba5ed385edad9a648777e98613809e6d39f01871e506b090c9c99e0e739dff8462fd3892fea58fa21ad3afcfdfa2533705f4420323485d5c11d0ee3cd75b54d98a1aa11d027901da95c654;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h70320bb7fc61275b5de7df44380b9cb00648ec725901023005d51dde5bbb073e38d23c83b35536030ca54950e40891e39b24002414942b4e60b47c4fba0f5fe8f0601b337920253f9fa9924d4b4c391330dff90784dc9d98fb4d507c0e007bfa63e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e73887d6340217954fca200623ecf526138b557c4565163d6c6508d67e7092ac849ac3060aa0534ed7ac37efd50d022d0c7ca5423da4bb0cb4bd32b01c745f5acc02718c6fa4b3fdf63e4429b5ad08f72e23e3e37c1f5c0ee70eac3ad93c4f4c757;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf20ff33b4dff72f8f4bcf6e4e78140a089b5b6457d96986dba6091e7fa80bb3c3d83cb10236e4bb7380c8f2af0c655aa138f6ef7c7a27a1ba195273c90842cb6e89d19eafc739e223f464d29a92485e6afe7707edd9872a8c59e59122fc3980bba7d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h796a838d3c0f21780fc90cfcebabc7d282ced7a0c713f3358bb7d68dee949d0cf4bb2ecd5d744045359832f50ca326ae55db2cb66e5d124ac5a0ba1c958779b1a2d43afd3a8388e3f1d3b1bd140f4451a495604fe6a90a2185ef91bc9b3dabcf9e46;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae8de668797a24bade26c49d190c5ea03416c5f685f605b847a77db476ebf6990d1f5e757b235aca64136c5d61b05bc85f3caf624d194d9504acd662cd6a0a638004b77012465072992d8a537426d8286744ac9335883ec401846a71104650113b0b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef7a8602bd57b306fa201d72b6adb1515bb7ee3e715c756c6df9c1ec904ddf1194338fa7b67e1a844bc7edceca7d781f3b59abc2ed1bfa960dc2553895a200f93d7788e62d4b7c2c37b22ae50a884fa91294f439f5e8a89729e2d442ff6a34c1c208;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99cbbaf2b4cb21aec8ff2fe2a23af6efa8efdb5793a628117e1c044a38a87ccd4888971e98c02208b3d8f6c65c71ab82eff7fcec8b4723f5b8b05b1cdd6041a35a3df1cf1096e670211c9da1d120f71c677a49794cd66e8556b9f6d17b8e382e9a1d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a69a5d0fa249b36f649b13591704014e9debaf9af892e77d5cac4d942e1d8e2ea4cc8b8d852517edc603a3daca9e8ea91c6acfb2598017e7bc7ba98913bce12a61aa1428d37f928c591612618c81bd793ca2b82e3abb57ac109065df78e57aab4d5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbdbbb83e07a909abaef91274a1d2565bb24ea4472a2678fb6f3154069c75c3954adfaa014f3c97f9f98cf199ae9be5093e84675917b50bf0d77fadeb3217adc02f8e621de26416087d6aad8612000abc049a85e6f52fe0963dad133129503bd7ff3b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heddc012f3402edb16186d202fe0845287194f661a0c541e9aecc56d2b02fee5b9c4ecb9b571b71545f6ce36c5222461bdf4c8ad5bd4534fc575820e6cf2d1ec29164e4d31f1d514afca25e597f4e10641310519fb8cf0f6e9d89eece5bea9502c1ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4235392b8dd91b16c1dec378fd84c183ab46e4691702775a72ba38c048767525f7aef10b1ea55af27d780d78dd9c28da387e738fac9fc69f8cad6220509d51665eb157cac2c5596efcc95cb09eb0115c39a01e35270614231e0bc6bd8421458699f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75538296f17f378b7967b63b337348f412c53e8cb272b183d1b568f14bff8db88c996fcb4b6910c660617674ea3d068d7e857c1ba589cfbab683bdaaa788a89083f6c221bade4c3f2c8b0faedb832f7473609cd2faf48205ff17b06b901377d84897;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43895238188d8eee451769bc7947998492a65ddf788b3ec38f443d5b88c7b3c0192b18ed6ffdfef10eda19191cb68ba0cc23e9e52d3f15971ce644d7398395e58d92d925d44e0412874e365357ccc89db549715f424567ae3e391f33082bba076f08;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88256cc472d6579555b4f307369ca79b3b87dd732f67bc00ce7c1e03f40d06492bd58f96488842f7707812bbf6e2948f41eb6a81c819d071a2fc049be04a16b4b792a0b26148526f8ed233b4218669983f66c121d7e7b20cba4a4de74c389b0a2004;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56fcdb6b401bf3d6864343b59b18ad0a861b718bdaa2856195b103b9ac5a6d90cab37052424d0f60055dd95e0b9b9ba5b17e00b682deb6286c7ea25833d55039fae77fcf6ca6d982d04648554c904996717b2ac156037fec81a89bae9fab2e45ddb4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h263ec3b734bae649a5216df6c7ebdcb275c294dfdac5e079baeba18f2f2457701a101981272e210dfc740ed5c3a733e8bdcfe92b3dfc7b665d1477e2665681ba959689fb367546bb47760f000704a1749575cbd0603fcd8476770dd830cfcb53b59e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16ec7e4076e41ffdf598830d0f91ae52df16f50d97eabdabfd7da10fac113b78aaf1d0de2132212a056813145ae2aa915fd08ba11bfa74f47de1536423903f76befaf1c54fd6270075445548cb7179c0197322e31f18fa7ba6bc55f1533236d01f35;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4b4f260d4220cb7b8d3a47123bb3fcd61640c1fd6c72b22656bc74f04f54f30f0a16d5d6cac9a9899350c9bd643fd2fbdeb4c0acb2699c668d2a1e6cc979971e088441d01a6cdb2b98da336b75ac13b8ba45028f97a016f1af3816fd6c70664c29a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha741997609372c526fdbf6c34a3c1d2eac3b524f2fd71b729a11ca41d49a771d1f858fa86c596dc061a7e52760999cd5daefa88ab6077cf537f8e4b32d42dcf06ad2f43bf2e64a3171acfc0ecf1580bef86cccfebb016b4a227cfc5b1570f7741314;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heeeb984fe26d37c74f6e91d26c561172c385551b68033bdfe958f12c86f26abe0cfbd852830a80603bb436a00050ffa6d46706d9f6bb88f30bfa2b6997f3bf877cfd4547e3eb0767596a167c0215e44b6a141bc813ea26d402aff34d13c3416ea99f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e54f4a67e4728e9b4dc648a3b2389f005e112b03370effd7bf9de531bcf60ec2dc8816f4b00495bc034c57fc4bed2f265746a99ca6d594aceb37b4eb91560003cd6000eb8c985af0741e0be6aab9338b569b9f74637c038bd385cfdbc5e882bab85;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f1624ada90f43af9886bb1e94f7bd621062a273490204c5de2a6f3b4931bc601ad980cb96821d1f83be14de5060253efe0ad93b1fe0cb84bd742f1176165d237f94ca2e52eb825317de89c93979cd4ffc908828f6f5298e026e0551b62bb02da2c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc484e9b1f21ae6edbdfe3b243ee2aa1eb72e4a383204b4c19fd4f44c8f98a6ae3b6e7164a6b1718ce71e22b41a3d21e0b05d78be7de435076b8bfb4644958962d65eeddac1ccef351065efc8edaca6c5f6ca845225c8ff32bf547ee7d35dc424eff0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h705c671e17de43eda7f40f57d0fa546f11f0045ef2572f4cab543e300e1b1bff3da898225808c00bd2bff93ce5f4ef12bcc09056a4c92212efc5d3588bfeff724078388e23b02d152290d5238c5325ad68fb5759598a03f7cb5779db6cea7ed7f0e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he30ca55c631dba829f494876332e380d32f85380706bd9284b13f22005bcf30b411d89fa5cbc0571c06917f75236714f7856c871cdd50ecbdb06418fe82dc85b52ebd2450071a27f83db7acf01a0d95e6d571fb8061b02a90a21aad4522fe03d19b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58508227956d12a8adce1d9a917fc1668b8579ca727234d7ab08aa571559f717432f855f7260d1e7d917c3ce70832f32302c714e8cda902a4d6b5a21d864543bb8a6fd315478b1515b750e9a0b34a2a093311b39302fd657bbb6af79ded25d7c9f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h208308fda0f36dcb4a3f01b2fec497c7c7b802faff97a82f14f7ee4d83370e9e7b0a33c2a5fd6e3738b5dd9da179226bb76bdaee2d562504da1ad4cd2d1925701ae603b440cf3d304b6360225ba4936a6fc6708662c77854bf6b84f7a10c81e00a17;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h200792c7f3307219780760761e56af1f8375b882e53ff925672f16b3a0f3a6702f9ba20a68d3e7fb1abf3c3c7ceec0a14298eafcf183327f4a751cfef2efa98b18823fcbb53eab7d39118b36239bb0d3ff0929507f9c8c0b67ccd6239fa850930031;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57ba2aa86df5e7f248a553733a1f82329fe48fbab2bb8c39fc1646032daacd45474f85f381767b9366ca0575f0426debab5dcc36ef79ff94d64d4aecfbf8ef438eac084214d545f04aa3a7db90203f5372c32e150de51daf388b7decf09af1fbd3be;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefa50956fe9bf62a347d85a7e350b6adc817583b318bd14608e223fd3ed4be88e28cd9f3027c50f2597d8dd0474384c3980647fdcbe2e801d56fb283f27c827ce5dbe488c4aac4cb18e9fe4e597b830fcd8802273f89e41acf1393f51514671e153c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c5b7b22e744f87afc075d1b65fbd9aba8e93b163af2c907f867e6d2df106acb93d23f649f9d8c4d415de2a31131a999377d92b67a3c34e82299cc95c35c27216276a21020df85d7bc0301a0fe9e7b9037e31b3c59bc53af9bf1dc0a6b93d760ad05;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8a2eed70d08ec13014883f3a4d6c46a9e92167b7a07f4d6e7c33fae8318a0c15457eef36e91706fff0a74c9685e91e84a3bc6cb1c8aec3056c8a835f793552c83a774ae8fca5c5f46147fcff5cf1303b99ef7d1ea5f8c266bfd61d9bb1c0d34411f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1575590b68e522e973868e64f67db9e5dfea002cc9c0cfcd6293a1e6bf1f590fdfa37ef0ec9fb9682265fd27d1a177d4783277a3909023ade4603aad210f6d0aa4ce5f76768ea8d3c2d00fd2e261c3189c41177e82cc146298eb5070e13f7d784f2e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86429f3a5943a590bd298c829106bada71b1d739201ca1e7018d4d91743bb417f4b16f77da21b9f57d86ee170108171ce9106b3e9407cebe6fd967029ea36777ab5c8ca75627a0bb8f96978775561fe1a3b925d7b51bd515eb0a153465b9b518a6ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a0d44f76a65c91faa4675488fcb0707af2db6eb60012a892c791574a8dc8266b28e583e92f3a2a038a5f5111516f6341706becec95447e4e44f0cccbd11838bd775bcc3b1f6d37cf1c093f4e50241bf6f68dc1185c80b07912d7efd348b8964f1f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeba2c2334b40f4daff78d07343a5480654101906697f28bfa3e626474342a3dec0b8fde4f65e82e1a323baaba321b70d5616bca1edf7009753ea4a6541c9ee96c655626fcebc7159b598102f8734d95889c1e65e34516059cdd32dba6e829f048e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7b29e2b679ef94057e3eb4c3e1eeeff22e71b6f4c455844cb6b57ffcf300ae9122585b8ce2d7216d284ad9746aa3d7690f724ebf72efcf967dd22c9ba5ece7c12caa82b2b2eb4357db606a95211e3868873e43290d30b2dff9045a854c2877e47ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4438cb739ab7687d38b56c088e10ccc53e71418d6223a3ed25b947f6aaa4896e740b2205076d17d49ce651d3ab663d652c8fa5141b97079362ffb6a99416326335082b49d3f818c41bb8f6a307c157d42d70057e692a178b77a0b5e733e62cc41cc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h487633a51e0dbb069ef1d7ccfa878eb212c220b8fef25a4f7907ad2929f73499fcd263162f6b51e55fd1c948ebb3ed91f1a76ba6c33ac20438b0440724006eba0142c4cf5d0291adc29ff383af69f75ff5a24a0ab5cc2e775dc7940bbb7f6774421a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc773e25434e9fb730327683902afff4836b19c05b199a6de7894f06bc5cb7c5c4c02087a3381a9406683e2c5a9fdd3cfb249696b52734a7a6b326c1f6496f46a3cd05e20886ffdc87f9dd774c664130480092c923d28111abe0db649c7779e72a7bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4413ab702df5c0597863142f265862387debaad3b69ae7bf2492f77ea3b4f663598b16a4e8654dd55a0a7153463c5d37c2a276f20c1269fce6efa90afc35a7e0207a46f9d1f20481118870b4748d7d21dc7c4c9666da8bfcd4f0cda7b9283a7674c4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e772303e05a9a3860587484b0fc31e5f3445927ec9ccd25603a4d76553c2308bab176b315e5c45ffbc3a1032e285c733f36206778b4733868e13e17c5f5070d0cf8eed07ede307b16444e9389f9b8416362d7da835d6046ab3e74e639302da0145e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h743242b4ae9f1718fb111436a958623c8b330dc67d102f6695976528d12b5aff83c6827f2b59b35f68f434b073a56069a209e575d3c9ec541acddde768f149fded3fba50e97abfaa74e0d4b5a02244dfa4bcf6d49ef0957bbb2be8efbdf77842017;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he247ccca6ace6c3a4df0ff47c5ee0f82eec019b4543490f1a42dfe9630f0e5d72a0bb7362ba1c6ad7fd8e7ae4d5871307cf5a695f516e4afa604405efbf56cbe41b42637e9f303a4d5cdd6874adf666ffbb7aa4d7cd137d718b9768fdd72964a99a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83313e2038ec7d8306ef05e9d8c24e398218fba4638755c5d713924f23737ca3afecbccb0121ad1ede2b016dfb83a77411e0cc161ca6e278e818ea189dd124f545523b2a8c591d1de522d42553bdd1a2b11c4f052a4b0f8f6b90868a4d5a31a5b22d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc395043e53aabd3b30a05de820e7b985f8b2c24f8f280b56beafc0a431007f84f179202ca26bcd2ca7b9b721d979cbc5956a074c3c9a5019d92b1835da3176885f48b1cb72689fe1313cecd74b191d95b6c6d11093fd4bdbad351778da5be871250f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haeeb33907699758a28bf5e92860bf43c8643ba8106c0bbf09914d9c2aea0e39ee7edd2ea701ad1ee1c6775d313dd07d2b403e71740f0388090e5bb14a75302ad01b520d447f1cc57d6c57fe25a19c631d7d36e65627af7f47548552a9b5bdc06d95a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a46694a8226bbbc42ad8e3dc49c30bc1a106e46e9eee08890999e7acd4548b8e1208ce37f0214b4b1b7da63ca5e0dd802b7cb7ffd6ab197cb13d9aa8d41836d6590c062bb7083b6b5c00c848567dc4a170677717b2e3933643913d19fa59dd67618;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74615d14e53969c40060ad70662d06343296da7ba8b89fc35d01f3bb7d0120a5a923f2a3bbb12e3bd4a2439d32abf9d16547be1ffd2a2ab9a08c8ad1e83aba65c44ad0a4a5df5b03c38ff87f3176d985da97a706b2bc517ddf6f312c551a0ea65652;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2256d5a3dbca3dd7ec0445d2094e9924aeb00ad1c8c7ae6648726edeebbb0cc47b9f42b8ec3f135c0047585d08350db758f3d4f2bc55cb2fbdd0bdfad7ce3b7ce0533e28d54e871e6f6a63a3ba5ceaa3edd756c3d49921a1a7f5c6bfbdc89fcfb21;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4adf499c5fc740d1874c1405b5656cc85bd08e242b2829877c814816815ea2a58f8a8d0504393faeb8e9e6381ee7ce3225f54a7570aea94c01ac1c56852671c4ac8a88dcf2587a00973248600843086fad47bd2fa3de756a07c01d55cc5c7a8bea4c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ba4ea3d9b164ffa5220fcfd2f24636bbba12ff9d26af73ea3c80702e28debdd94191fe89b45db218712aad95769c0e4af82ed5127a9f723942a5497ff80a5eb848ba8e0622ea931b3bb64b327277eae7eca7a46013f3faab6ff8ac9ca3ecaa09a54;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha624e669720063940e8490af1a2f65b7719567ee727f635869caf998253473644102c20aad19adf46c4c48dc2b327bea4b0cf664afc4bbed43db5442d9602ac868a5f1a9210f999cfe689ffec3d3afffd3f8e594d045d368fa84d666ced7a70ed6e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57eceea49c98f6d1bb5363584c4a508abc959fc069fc6461e29d26f8ca20aa2c09c7fe5c0a35b72053c8c25fc4f41fc9b159520f9ee0e15591d39d3b5caf01e8ca096273eaad79d7b0af56fdfded9e94cfecad9003bf19e6194cfc55f3c1d85cc59d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2087908567ba7b0677544a5fb994a92bfe1a2e77eba026e108cf00eb2b5e65c44826706655ccc56e552db206c99b3da4b9b37ee60f440698beeef61a9b7a6c8a0132288743698e92f9457ed655d6b03476db22f560e30a07712b4777925a7275d98;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74c613c2908007b9c4ea132b769b25b4a604190a5cced1889c09c889cb6798f59313c8431760f314b693bc2e04e48680a17af64ae1f267a31dce674e9e5b166409c517135b3a63fafe35e5ba3bd6f33fb2ae9380c68c45a606aa62e7e09220cbaf82;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8fada3af435bb62d54a2d981ec15d98acab4a7314c77c87e3936d2af7f3a47f3d7cb45d5faaa366379f4c092702d5eadd47c72ce3823149d53cff46b3cd0600208df57ee6b52dbee393ed762127e379c591c589926b836ba4d8a30cbb1f9d497159;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e90e764055515a8f951724690947fb8a38cf8f4199aa6da9ab3272972177529bbfe34814c00dee6aa6190edfd003344db41abab7662f31f61bd76e7755c4c4d521d098f573d14e94c176e85ef87ca32de3a491e6f58be44e64c7132c8aa60f112f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4694ae8d431b21c3b2b3d23d28335cc62450be445ff08ac85df7e85fc0e3003ba36578c6d8720e54457d9050579583db11f9e570dbd7bfbd83f2b2a5367d573789b0dcb3fe62d21c465db2e1ac1f3d1a7284ccf141e72781bd526ce8f2faebea774e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h721f2392c8a886b2d3486703f90ef6536ee5216ef1d9c77a6138d017140c4aa7269e2bb64896b6280856ae340b848f5c239cbe5e376aaf18e374bd396763dc4e9f859787012ff7d83e37739579a836757a9eacbe693fa20a26fc463c263583307360;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa450e8988b9126fe3988eb9905bd4ceda919f8a4516887d0dd6a07afe0af5faf5eb78e9c2b851e67c559fa7efe56bf9c702ff20961d7e5efaa10346fb1d7021814203cd9c41aba291b8b8084e4d0946b84bbebdfa2dfb5f96d5b220b038c499a215;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h373b07120651b3ee9af03083a70213071c90c8c8862215f32c353714ff3617572712d26375b65805737211142ecf1aad1e9b2aaf4cd8fc9483a099f542638c34566e98f00de6cbf91f04ef9688cad16d09eb71ab552ffc38ad6dff120dc046de4223;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b9a7870469f9aeefc5b5692b45c366f3fba803a9cc5e0ed6d5b94e38608489f97cdb979bc607bdb54ef6daa68b971d3f69c2f8f50f6b5d7fd88f2a23e720cbdc9b3deeaeb3313a3ef146ce72be8a98e6fd3766396364b13034a533213efc926ece8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50b998a4fcfa36df75b4e37f95e77b408eccc761bd7e4611a7c14673841ddb7f70db67677d2d30fe4d901e9786e83e05920dbbac8bf29fbcfea0714fdb0b065c6d7da18e25af3b8c58abdda68dad0ca53ef29c5bcc4d54e6fe69485926eb21579008;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed07e194fc63cd7c92634bece3252c0bada1be4bd6c34e550040f905f7fb24ca012500e44aebace2a5f07efde90546da83e749af432ea02aca6a192ca08b846c4769595483efc0134b9776d544eff49a0b4636ababc3689d7b54bc7704f95531ce94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0bcc7c9b7d8fcc2517f3eb44e767159a4c54c343eba7bdd545f7942a5665da7d9967514311a7f04de294a8ddc68dc51c7552a28b84481f1a3a4fa5a97ad42c732dbc5259821928b167aa1a4ac4dda41454daacec8bd32790213dc100b72f67f88e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c287e28679c0cbdaaec1aded0027a90d36618639c1cb6bde483293cb171d4df2ddd9a4338adf994bda57e5a3bb22ff72eed0bd021386ef96983db69f7afcb017503d889bc168ae8db494969f9e1d57ca9d781dcd7b2ee5b9842e1a7673137cd0da4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8bf434e4565eaee73a3f0e8cde1ca40086f3117b845c734082e77d09ee8ad57405e28fe8f7d3cb6f4994b5056b08b20b1bbc29244eaeb01cd20a77509024dde353c51857beba1cd7dc07a224ada318fe1d09aa040848409044410d04f706d7e34ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60545a81494a31685aa4c00b325a219e0cead11d2c270b2c7bd140690e57e36c20b0a06d190c308d550f7a5b6ebb73fb75b753e679457335a24909f62c855c091dbf080c51d2b15043a229e19dd3ffa64499440952804ca25d1e5189e5332a86b863;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ace898371a92522c1a686801d6e5db6786c994314bd33653842943dfe68453aae813715fbae9c722d9e11107d6464e5e35494db25e8a853fed80b99ae0c718e3d783fa2e2dffe5237051772cda219e41560097b56fa64152d879b514fe30f96080;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3c2541ce38c93fb8f063ed8042d4e9551fe4a09def774d58870c2d2434b53422706c93d3c16099c4270d0913d873b4f0550e67fdbb42965670071547801c8d5f5b1ecacc27b377c9250e1f45b0b1ed243b06a05ffb6773b30ec6e4972ccf8d07228;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd59837014b17034848792204f213caaa8f065e560826e9360913f9df657f0925dfae1f86f8b7f73bb2adba99b8a5dc7fcf766556ad8fde4e77fa57188ab1979d702c913e8806b4bfb457a96a6c58acb5ea97d85d4eb38eaf1fe9760f18869c034148;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e04f68d8a0bcf44cd810731f18719884561cb315ed88ac307538b855f6601ef7c09d9a7a465e82191191efcfc2c7f18adab29893161ee1ffc2d457772e1f82c4028065bed6e6ba3f43f7465f81e0404c8c61b82c967bdd83af02dbc140218509ad3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9c4aa1513b2854bff483c871d59c3f0e657d1d78f4c4c5848e5cadbda2ff61630268b400b2b8efcb71aeaa86bd8fb7d2691d35a37ea9e68d30d54d0d3b80cc1051f4426ea9f0c5b4308e839cf7782bc3691323da81fbf5b244d583de7cfa515cc0d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89417c4f6b86411e8697e03166e6ce2b315509555440e279989da0b2927a3071649da2853d3543262c6a2799580450e4b18d5c0e0c3e2bce551f380017616b86ff5cd5d9c01bb66bc1d2d090c382b1b75d6f742c094414919077b10ddab52fed3022;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b88dfe30013b766dd9aa2d6071a7e54f8e589010e43c4f40b91fd31ffc6c8360d5ce95b4d15a44e09897a0baf594d715a151098d3c193e4eed526bacfb7050c3dbdcd45eb72e2cfb1ccfb78e5904f17e07334f55ecff905c96ee6b5841147c139e5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd84da800b64aec23429cb1e51463d89416cbda2139334feef51f7db8eabb80508c7dabe95c37d570bd8cff0f8b1936d785f82f98de05c4ceaa4d57e4a41821ec6d323c8dffd52ea82b0b879a7bbf18a7d1689af3a73ec302861a120201b360553481;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8856715ab03300e545332bb2a51a16d9582491615ac8598ffe240b215130f90477b58d5da2a98262df9942fc3634cd19fc321266b710f10c86af0b65f722b7d9db4980edf5642127b6bde4f3fa5604530076fc75ae6e84156e29f86474ddf4962346;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf616d7f61eff3fab7885c416ba25cee2dac4ea21cc86f13f8ba39eed4b3af0a443ba32d7bd581f3e184931fc2f3498bd78beb94d9e0afc92a9b8e669cdd7ba7295ec2de5d6ac20f326c59118ad71dee5f004138ded05cfa2458c7ce0ce6c8b0b524f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0719a519afcf404cec6a1c3d01c1fe101ef679270cbea7e25d6ddae486f1311268a0e326bce67e090770184025bd6079f2ca61c4f55186931a7569e03da623ce29170a2f3c1d45440bc8042f9a0d4a160e4131be1e665fcfcc3984882a692f45934;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5623bb83b9c795fb863491ae6435caa413ae6d53bc77ff2dddad491c1b906491c935b0da34ca80b5592af4182dbc2163455aa250c7a887739c32dcc85a8dad8f71d9985f364b4b9347f13f46df00b60baf0ed0c2efdcbe266a2084db40dd173b0d73;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha69e6a13fb07cd6214b6f30e5bbce3d0968defde443a0d54283842a782bdad80ed0344bed8597067ad0775545f40b3e90bcde2aecb51b2e78045103f8c2ec8182eeb36d749a191f91416ddd0d3fa78b55bec8b7924e1fedbeb65152dac79d105fab1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1dd03627e2970be083c41bc187755029c80774bb5559b0bad5c49d153c8543178690ad6e529d8abfe65a6f601c5398d714f492e0461f1c54b597fb680f748f8988694980d4f58ce6fb3aab5028340a67ec7c4432587708400c15f0c7964a7f97ef31;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h943c40c4b79a37aa83f2f6b2564fa54c596fa6e39fac261312248a79afe4443641c82b1ecc07deaf5d2f26ac0964914f0be68b0eee21123c3481e8f7e576c42e34ea982f20e3cef217d7cdf08b91198e970e1e0b654fd803c904ec3e2dfeb3455e67;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc04f1947b0abab416616484a80b901d34f174cdfbe75ac75f644c4d85ea92ca69361045e748a374395906f77f5c36737d9f6842da9a7ae9fcbf3c65c2ca61cd1afee5a0857bd12e7a5ed7a1227e2f999772d0561e515397a094eeea8cb15d9062086;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc32f32365e5c9852ae9e49aac56421a162d7ed4a54bde35aeb6db9bad9efc4a6447cc723803025fda021f0cb1f7e3ccb18db54927dc4afb4f3d8a58e16e8fa304a821e23c2717165a07412ec7924a40c4cf21b350afad907656b48b199a7f8f7945;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha49084343d3e07e0d54f34b9ac4f7f3965277dfbf737deb5dd970bbfab9eee6509e79806eb4ffe04c6bccac6157ab3d484099e04d4d3ab12d1bafa3472b2df95dcb22d7ea477c765b6bfe346605acee48351f0ff8963cea57b03471cc7b7dd536346;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e09ca2ac422893b660b08c6c510a880c4b4b11cdc335e35c511c0d41e505ff9c5cbaafd00a7b80f0c6ea9d9e5294a8fcb3f8fe8048e0bbbdad8bbd222dff004e465a8abac9d953cb8a2ed9f25939e74ecac1bbd43d8cf329cebc803496c1195a6dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a68395bb5b07da7b6e5a7b859a9e7ce9af869c08c55d217fd61e6b0d4639ae5e5278c82358535b612153ed2e1562afc1f99cb8ee8c8617341f947960c3b0a62508ce4b570decc4aca6044a4dde4581ec8fd1754196f19b216b241316232e73bc82a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf52dc5bc8c213cf073a8ea2453abb4a49ca2da930ed3b3a93916325eb1f500918e9b5b0556e24d5636d11d712b5aa3513bb1dc816c2d3bf646c3c5dceb57c64b92e7f8f7b6973808f700540e9a2ce26ee25a7affe8949535b44a83ced6ef6057409a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5613c67573f61b982ec39b81bd76b0793d4a76f4ce3d4c5369a7e707bd0316ac55cd2cee560cc84f595726ca8a24df5e8588f9427c079d8396e5f3c3dc5c7195ef959690a2cdb652d9ddc866cafbdf4fb9fba05fc3e8ab8f819533c674f87d108f59;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15d5531ce9f1f0bcf622a3f6e166ca2de8926ff16baab2747f64a5d40922f6d3285f10962124a4be03fec45c2b17609008cf441006515f5443d005199163e6a9a80376334fabc450c0c421ac6bde241c711e49a6e51c497ee0c52685d836edb51d0d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26a8a84a364b1db6e5d272b39bc25dbf919fd0d62fffad655d66a6a4b8e0d6e8ff648faf68d69674e50025a5ca2ab1aa291f2a3df730c1670e3c55bca94608c1ede3b98c4b88495d58bbb38021b064e9ac9e74abcf27239e9f51b83db761799f68c0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd5be36150bccc7f9ddb70193a22135fa744576d632201a47dc2cad64ab67e98b9619a2c046358c38dae6db92d379f3a362dbe39361aadcb873d0bb19b2b6e31dcc98809029fd8ae2aaef13d52b6f8d17b9736902c1d72511fd0b5ed7cbcd50ce80b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h806cf46afde3e93c643a8472b0d6b8cccb275071b823ffa6c04ed915ac06dbe9f834e4ca03803ca5609c66e25fba74a9a9e37d553716c00c4885fd606ca54a55d98ec2650817e85b27706a65bfa97012403b1064d01f5b7aea59dfe35951d2ff7c52;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae96ecebc6c3ece6c701f91e1f8c6f23c2319007317fe00329f0d8ef5d33026a13d54500ac1e72f83d81f64a1c3c074b69df9332a57aa5cc3cbc3da23ab233cf36bab053e62d42a7d2ab2732c29744df714c3e53896402941327492fcec5dfe7a33d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b607349cf0ad32d44e3172e85942066ba9332de5fd6270d666d091b356257b1dd270c9f3c5f0880b5e9cae80d5d61ad22ff82a01156845444b050861917dd4434c8bc365c91baaaedeadb99442df79ef9d719446df50d96326a2eb6a6ef461e515;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha55d9b76870598616dd3dbb51dc6d22578a2c68bd7e3f91b705d7230dd179dd667265479411de98df7a143ceb61c25628eb47d55b1f556d52325c4af259e9a96d152fd7fa1c920d8fd7c5b985a3d12c6bd6fe89b6327549d4356493eaff135d39e5f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13846523f6c27f8129f0fabfcf0d67bb511f431a7ae1077b2dbc284d707e958e6c5e76fea3e01c9b2ebb11729cb9751194ec31504511c613557ec5e3f050069c5d9d94208018ab86f8ad8d56c593635218d1c8e96b92bf9caac5a55ab863309900e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97241797f8f3da22a58fe61963f5d026324d61245eb6ed120dca08e5529b8d4f5e5d9867b8d8688988820bf69a56772f464a7543e7827d1e90f4fd610f33b4e1476e347f550294f2f048f56f6ebaef2337156e1277a68e993ba73ea6a3ff9c0027e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d9b1bacfdb2dc8128cad3f368a166b3d8d7d128e510b0fdf3fd6293c9e5364b84eaad818b749da2c2313c18c3e57784f7bd3b6f55a5b65ea633ad7910a9ef7e32e45454b28866350253bab0334f585093ebef92ce4e3d92eb1bfea0910eb2680a8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h867f61bc2176b41c6e07b369e7354d4a6f7a1062fed3624a7c633209f258bc3b34a6fbc731f70dfab521b745f0a02c60449c3e14f93a9bbec6e171b5767d42434dd241eca488c2dc689f1a81438e329d34cdc0ba5e7f5303acb9902b2b2295a662bf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b5599cc72ae27f72ee45c2f7afdeafa297a25c1ba875258ba82e571b5ecf51174ef8eab7063d524e1ec1074ba2a3c174adccb029b27603b23f686443b3cc23828769638dbdc14971430d0bba971bbf39f90a31b66ab4ceae9b26b714c060795594;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b59f86db8b76c59b035adcc7d8246db35fdaa5d0815b06df0e32ee350b4fcb36986e4c65ea4d68e327f2f3d9dfab3bc73e23cf9f9ebb46e086e0aceae78021f0cf49bea14e6b1904b44a680d33bb94d4086f7cf25a8c4a4c417e696261e147ee390;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9aa75788886e52d2f3658856fd1fa9cd21af3472f5f5d1e14195501d83069556066c5b3aa9cd672073fa7d6c739b7ba275f90ed1179449b314d5421b5c70a0ba64d853079e764a7a4ef2b4fdafa0161857e334c030de2605c67787f82981c591cf6e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e79f50666a889d531d590ffba322f16ae0f5e5a9d4f15ad61b139f7f5346a65f88f1031b6670ec41d4fab09cc61802af2b323332b43bd5ecee945486f7dbbc05d4fcd07c2fe6a1162399718042ef2a5654a27806af854f667ef71b2325d558bdd81;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ebc926303a452be74d6d7ca5d20533feac81eeac26ea6890e638168e42594add07be274c94f86d25d65de6d2e8500de4710bdc6489bb310c350340c9d0ff8b1a4a2cdab2b736e79b8953b30120f4890bf9a86dd227d76cfaf4a90b2286e7309c7b6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51e5f1ea3713ed5782025e573df838358a8a8c1d8fb2acedeadf24b62056cb05767ae963c9dbb551c7950d6e3a8136a404d93257c5842036f0147c83d8ae01cf2df8968a56d0d84ee801979a89c00b5eb2693196507e747be1d672ffb5e32f67bc94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ec6d43a9303407d1193bcd2eb06b532827844bccacc52e8f836db34854082c316b96c827e4789b39213e1264e30dfedd67ffd868916cd111bc3845491382d0c323fc8fcb1f72b8801c1d1fb0550c99632eec95e9e126b1b3d5026c7aa73c2c7da05;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hccd1b7c2e5b9af3f41a8f72a6f42543002f6fbbbf40ec8c91c5d75ac639356962b70a36e5a96b81b9dd5587756a8cb52f59fb1ae57602919db1a3e18640b0417dd67603469a481cbaf2b8ef99bf918b0e9fc09793648ed1a0d6b3831c1b24d8a282f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41e25f8c71aceadcb41545b17fb9a6700a1fc72f8432722bf75adc2423c95bc2323ae24beac42e63c2b77e2638136914ba0344276ff17c39ab94638782b90fc7a7d10544d289900258f2adc51b69caa97ac4b6fa310bf2e10b17601950b3f4950481;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd729e1fa46f437280fbb7751127c5835f8bc09e17f59cdf71e6d372cc657c5fb9ae5e9c2cc4299b445ba7c43b9955df500d364cdddce274ff473467c3c8d1307b7fb1885628856e80d0c06df7a36223d7f557976ea68c4e5ebe12bc8ea42a7d0947e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0c5758aea71e8aa91da93d5f08cc1fb901a4559841ae33a4a61378093c6e8572ba55624e7bede0bdb267f7710cff13eaab9f398bcd9d84b881207dd041a0b60ad4d0fc1cb9785a56ff62abbc545d60fed5fcce671724ff4f54caad15a67a5e50e00;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd6bc01be738d8fb7c55fe0797afdf14aff138089f8b642bcc9f8fab8f0a1985e4cc9412919465f9a50df00dd4b1cfbb391b7764324ae05065fef20100ce5040bc845150a21d7593712a47e9a167ce418947489a5a0409982813408a0020e16cf65c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1178f640c543929f0f1ed336df406b99191de1c5e1bfa38f4b789f1f302458551ed1ef3e2c3f35f172f213dd7b10a3825d24250ca8b6633a2b4359f54ceaa01bc33ad9efb263487c8e8561711552afa0011d23daa5e6185c6d2624bd517f2acd856a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc73bfaed765a36789e6b839c00513900483704e19db1e22ba4ba7930ddc083bc9409ad9587564e7c8248c6e7e971c47c43e412245c17e8c2a89492c26e7a6c61fbbb0c5cfdf5936171f12196f5344fc25e4d19b06516051b98217d0319b6cc3ab9dd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bd0439454fc9c3443eb4370241cbc4e03397b7de2c16bae57c75bfb3af5882b5770a7a8d74a9d754bfd1ba9f73b8d388191902fe8c09a36e7dd5255a33839d164e18522981c994fbdff6c708cd52a3fb6a6fe71a00030cad12af12a5efffc6cc218;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd813a231f347f5236c624e17dca27d0235485b7600eb529a16188f67fe8af10c25bf320f128fefb0a9d6eb81615db4545e40fb7b652efd1b79652192b69cde786dd4c8687621377f87d1ead4573ca50e093854d9ca5f8f2c74d8614cbb38e4f1654;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3fec4649defb55a3e0ded256070a687ada86c5750d7f10ace62119e111cc6d2bb7735f0203e57eb96093cc8e5e454c9e681b98d04e58d7d46075406fcb36d8e4519acc7bf6a62437acfcfa09e3534ec6851d07fb227470b690bc515aad4c76f6d24;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5630eca60b6ee276c0ef65a42508d27deea692e6667f5e000d79d97a0bbd96b7b747b47cf1aa86ab3c3e33b93c916ae595773118f682974eeb6c8da3adbd3008a67a18fa881fd4cebd238dd8f4067a8887516a450972af2af745dfb9907b4d211b16;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47251d62b33fd083d21f73a87ba7235cdad23774094026d8dde512b29c81a4661cd7d5af8c9e7516fe658df9b17f882383adf8a6f9fa4f036b65d80041e07e8f587b443e6d8b576644a51800c93a8b4b2f9d322a99c60cb10e04a2f0071efec7cde8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60b22bf10bb5ec30970faaad02f645c4ba3f4edaa20c9112ec22cd8488e664afbd434153daac45691620ca4ea48b42ee4da50b303cdb9170f80ae16edf3d04588e50c4e9d040c04521a4faf5678592470c43109adf696bc57e60cec618c078ca25f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc83b0e128f65764e0bc2fffe39c13af3d8f99aa68bbb5b3d66c5d6c92cd97e69f5ef13cdbfafe88fc2b68076ea9c9e47488bee3f09c4dfb8ed9e573c7ed85c7a5e81f000d9859d51d9f648e921c4279cdd9d200c00746a79f833132da25888dfca38;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb76ff16ce6f293fd9e776952964d2eb89758be77687086bcd644323916bbf3bdc97611cfa667c17073c5126edfd1ed11af2a0b0986ac9ccae553dc5750ab4a99d12e318fc2832d314113321cbab73be5b695ca169a0c7eb0a929c6f1982b93097bbf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8817d62f6f44c76f97f3cead0af7dcca7a38f207e92905eb27e87843163e1f23039510468e41b40a14b12bb2f261fe084a1e2042bea6ced53e310762ee7b3f5578eb0f9db725b386626c628d6f312b980c940c94bf21f8b77f35e9c8a6eca9a5daa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb960327b105b82ce137fc513196686f5f9fd3efbfa614a3954a3566cf1e44d75ace8e2277b14f53b2e881fa538bb422e5ae3cbc1077952cad27f3ff1fe74aa213fac7314ea04a4e0c337c4ee7daabfaa5186b85012825ba7981e467037d4489d845b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h254a4cf80ee36af872af786dfb2225c4ac48027b1909afc40a5b1a2b5d00522c5ed054eee3bd8342c352e1ac0224a59b77ea151eb05284bf7cd30c335966710374c648b4d908b4ba8482b8782267a51dcef93eed5d8cbb567a723d46f60b937a68a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8df7a9e68592f16a00ac2c5883d09dcb1473deb4dc325c74998c5166860378cf3330138da746bd72444afbf045aaf5c02c9d04d64ce92bd5033fdcdc0180e5496e42dc80eeaf9437ae749c513c4d5018bf4fdca9fac3e9a9eb5a1d42d0ce889fd544;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4a90fc8f7130e723624e6849b2338f092d358c586c27754bc48bca39e59a19e64cd5fb66b9c4af84b0d14a469fb56165a90ae4884ab786214b311ea2bf765bbcb2e5ddc82a3d2eb9df689badc465c3c68c930962bc0dca00dda2410ec142f7513e0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h440fbe6549ce291eaa55a9be914056f1108124fa6e4a8ea1541452b69cbfd6d6a21f8c30460aea08252240fbc532713230f518334251dba2531a9c5b9dc84302891f72ad0d2cd093818b3cd9e028b4bef1f481fb7b7fbe44036cfd9ff8f81d51883;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h277ee76b04f222b5c56feaeb4c257ed371e6c0463bdb81ceb31e4337d20e09430d046634c30a04678d0354d80c865f9615f010040fceaf7f41070c66f3b8ffe17a7b991424af149b0c6d19835bdcd0db720efacbc0112afe97823a81c0d00bc9af95;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc933de9f9cac5240c83fd74803a107f301251cd744f8b55eb1a1d2418a7080aecef17e3838e56bafba31f61d5942da704239da3c2e0a55515e4a9727bf0a8e0cb24186d284209d4119b18f2e8056768f7cf0ffae1053a3dcef69e5f77571885ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d8454096a011ec67a04772689213550240515b13539b458c61aa70e70587fa3e6ae5bdeae31dcd8456557d7c6cbb6c5a4c9339fc7f19940a17788d5cf395f9669120da0f287fc32376a17bf7185af1becdca1564f2f49acbb4201add6ff74c1bb5d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5142dae4e9848f274cfc136779b323f7683ee27f26f72b593d5c4ea0daf5a01c55eea64dbc0f26a8bf04fd77bca2373e985b66f5b74f05f274024b9aeba62b6bb754a80873d62e96f1e2fea6b5056ecbc33980cb6e1d924eb325f7848987bad1ae69;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1addd36e8626314a5a96bf98131dc0fd35cfd7811a3557bbbba4459c2d94f2038dc233ebf2140379fa8b790b5e137e2c98ca5f150c2941b7bc8d8eeb83e9193fb5fe4e2d04eaaeb5a5e6d9a8671fda404c7d677e6f898c64ea6692507bfda8a9f372;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7a6a2eb22fee8a1562dce8fe8ab1c1bd99e917230ff1a8ac3b85409bb9f23948d26073c01333288f909564c46bfee78c0056779b03da3eeab31e19e76f7bcbd7ae7fda1374fdb722e474f8d71a2c607e3a860af8f90abde95578acb0f716db0d300;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e370b8e0d83a9fd37804a4ce242e40e5f26039e9d66967b7f7079c747d3612262e7fec925f83069d5ccd3c7d995bd7f994d4249214bb9c0c603199bc985293cb8879a6259ad23c40a7779d2df827ec6034bb8e8ba73ec5e887e9da56f3a3fe38c88;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a5e986d8a54896a3346da4e1035000e85d810437981203bac915941d63f4e6a3d94f0ffca48fab70af3db42d5b0b255f0001b082f8be117a24c795b624d00f9913d8754c9a2a4c1f55f549173dc2d68adcdf94cdfedb3684a1fb08a8cca06f7aa4c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31ed052f38c73367b3e7a0de54460ac1d53b9c986a62506fd7415f1458c3c157607fef9f3c54467b5f375a0f65f1a99c87b06682de8d6e31cbcc51c3d162cb740940315b4a558a0c38542321dba9cf415429af4d9a23bd113d81f4e5f9dcedc484e4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebccdcaf63f18bd05156031c5ab48c51e6af5e6a1a03392c7b1d3f28550bdf4a32aab28f1c7be43d3e6a529a7bd359c8dbc3e3da0324126aa45ec489e9d5e24943f242387293713da0f9b8f80a75db2a3d0822c00a34282e281b8f39f1647934e800;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2fea2a68fc1ad40d453806d35ade3516b31c4997f81bab5e94dccc6d0173b0cee361bf4f6efcd77577f5c3a5f794ae7b22dcf0500e9db9356cff93aeeff78f2d98859ba19f35c8aa494b09369f27599b8b2c6dd069d79035e57602f8a4941c78d65;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7badf63d0f557782d4ea99bff2829d68baca4bb52e05dc10d185add6d97e3b07f684b0aa7d17b84de3567801d54813a59cbd98f373030fac8a3e97b44d3ca3323d70049c7cc12da7b90a755c3158b94ed05df5618079fecbaf6a1220dabdbd63758e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heaf6afee71efb6dca5618d24f19108f004f022b4f551486ba2c3c6dd794c142a36e99874f42c2f7dbe04b471ae647a42b3bdf30895634005f3dd519f03380fe4951cd1a1a7a50c89ff12c54112e3a763c332123e74909b4577910fb5398e6229d006;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8bd31d94a4ffb054021466934e9d118bbc314aba65d568dc49148b79595b02a1228124c29d589dfef7f207182fbdc62521c92f90583d7bb05123b79fb15ed462578b0e41e08c473a13bc63fb131c4d9172a81bfd5931cca67964bdf3d91b4555f94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfaadfca6849e940e48a0ee6735df15b77b2bc900fa9807ccef9b853d8afa319d16addbc0244f6e5b954561698b9e723a1af426329da42a0ff435eb0223c29e9e7880bda84ce18942741f4c33329f5a5784f347db95f61d0dde577b439ce193b8f2c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b5723ba18bfa63841ed2aace869bbc771d43cc1ac576cfd1c3cf2c00d183b8757683db0468f73cd86b982fa14f139fb522f0d6cc7baf5d8604287c9da07911385774cd359c31323a02d94976a31fd67a13671a356f191daf7ec72ee08a0566756dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd704321364b9e3abc4a775fba62df05bd5b6fd77f39b8f1fd2571957d2569fbd6f29bcee2b5480e8c856c6b935b7b5984587a8af6088c7009f5d84c13373bd2ce81279d87d1947638e393a5f9f4a8ed9337616ce152d4f34b9d295c42785501c25f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5241d7c1fda243fa5681c687b74d72db724e74cabefd77368c17874cfdd98ab3493b30d7c8ad6aef13b1bb31cd692aadc0ef5ceedfad495ea0718fde77940b03e595e3cbb0971298fbceaf278a663aa71abdeb74cc5911febff8fcf68af6f36b474c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9d1055ac293dc0d599c70b4e39e39b957ea563f13c8cda66f18964f6f233f56af3c3134681221335fea124d1a7186cd71a09479f57345081bb0f060a59a75c91a289598282bcb1d97e06c62ea38e8dbf7975584c97513d983037df92474021e750d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e86bfc3facb6af32820993b86ea22e46dead8190a5eed8174a833ebfc7316259faa7fe5efc8f8fd07a93bb6b98d86d8bb605f5acd0fa0d740f27405c7459301547f9cacf21f727f6844cbd010ec5ab7ab44eba26d5906ede58d96ad37a78a519047;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8474c975804c9195be9f3e68bd72fd43dc508dc9b3b3eb2ca7982b018981c52da5804ed83578a84d79feb073ee346a22f94260a0fb67b6319785879cf6e2a717e728c706d7719c871bab600c2de5e3f376795336a899e0fa60b13fc59ad19e25b94d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a5beac98a9be37a6d56c8fbf12040604d6bc920286ce397f15d3b5bbd6c85b0b566d7253a1a37a3a54bd79af2ae7e0184a063abd2e0eb6cb9dc5319616bd6876c4debd16e4a476adcc9cd44af5bf315afb6e87e2de67f03ef2e15f5857f75a322c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde9f9f799c0fcc0541b61ee67f721cc8a8109c8cf2b174d1f3f49b70e099e20df020f8b6c1727e41797c087d3cd4a084c3ed9ae7e1511f19552f687ed07352494b531d90600fa426c8c8a80eaede783253346e7e7a6204de4a4b92e4fc23bec82814;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c875522baff1a76a0930e24f36d8ab7db699a11f7eccfee187de7d3264a6276b7afbc9970f08ebf6cafce138f4592415ec2b3a10f9647f280b4ccbad48ee5ed2b623e4b3592107d3fe0762931de6644243c8b8d87b17a80cee5bdeb7a9d34c888a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f7cc137c08164f1474b7b562dce3e3b13b2c080a0306b9d908f415f4c43cf8575ca612fcb97ebb1949197a389ef5691d610de517bbfa6cbd465f42012430cfe774329cd109e26bfee52d01f2fe2ad76e6a459d04f20cc56b4a697c21ce157889873;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h970849362655c393f28a07b322f6fded3491297a7569e25e3d34f76ee01b1dbef1d13cf9e4c633a715cf8ffc43523c45a7923c5341d33b3cca6d8fa33bca765ad1f9e8dc43f9e6bed935156078e683057b334ec076372b8f44afe09404ebf59b99d0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99a20a49116ef75a12c7372bd2bc7ff57d1d14ab2033a72fc62bf9a361d77577daca959caffc3bb52828f3b12730118f54cd8bbcefa024564f44796008f25aaa096221980d248e91f6849dd24188f46bd713c900664b3ff635ae0de038f4cf5bfd04;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h270748275c055c6b84fde45193833e78e1c470c052185af3b582d8831cbb71bf6553b533ca2041cd01d997b39931d4a36aff5fdb88a5293edae01663e2ed2115deceacd2372a73203a68a78edc6448fbbd0ce72313587e113e5b8c4c3e56e8ba36ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h290309541b73cb8cce9b062b7471b67bc03069cca03736728675bb7e9aa9d7ec89fe34b5fd3bb12572806e19850ba82cc0c64de35e8b88d4da80e8d8f1ad5f45c9d575eaff97d041fb8d7d0731f3be3ec626b3dcf03f127f279e2342cdcec386e179;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d8f73dee846e243d08c54b637f9443729b5f76686ce4d1d54886aacc00eeea18c18e6b9690ad1177ed39ee847531394f342ffed095248a33ce70e50513c01b699bbb3bfc8abbb32bec5bb597be16c8b2f609d081ea3dbc399cdafb35ff3992355a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b6c1564b29c16af6650e3919ef3f90947e91ea938cc3c8f03bf4fc14319739dd537b08629e24679e392f886b04d14fc8f0d17c6ada0c432a718b68fa743dbcfb042abfa0e0312a1841ec804480d5c417e171ac831b25992f8293246866ea23d33d4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde34aeeda3a806c7f191806baff35e539eebb9f45d0007b8b3f32b9b9b598635b1fcfe47cf8f59982443bb1c65952de3cb2c54e055ee8dabe57006210e4a69f5e502210f67b82fc44c0e935a90ced680eb2af406a8c90f3eb89121f39eea769c778d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd03bec758977a5a2153144a421e25e6736d6352cdd6bf62f71480cedd4ceacd5e132d3ef16b56f225d4e9f655699c54fa5fc9c6c5b7b50b276a4e4c2450056b3383317ffd661cb1c5faa74c7f0a07c69c35dea2448ce7c44e6b79ae663abff7c1f1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0e350c33a7b2e7cde1fdd1d3e81d9c46d97ec1d10c3f4b6a053fa08c6e03e16ff1d7741020229559afd5440122adfd907d6957934d8005d8df73d6e11cab719e3b2c6c6eb268b1abff55620c6cead940badcfc988c68b9e178796eae342118be1f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h241764d513f1f90eaea27e67ced1d3caaa328ad3782ed5fe48e6eee5b87bb1e3f6ce0b891f169da942786435554882a76e2a23ee5a306b75ca47e8018f355680b028db2ebc777b225bc325479b64b7a6aff0baf56562a9a7de7d56f5aa8491790f3f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c2ad80bda6cb9e0b0eccadbcfd6786f1b4d22e4fd7bf33932dc81b202848f7f452df08186231704766b7a70c1e328bd89c8d420e247ab93fe0639ed196502246c1eb6c3590671a3a86ca1eed388245b8cd0ecd30af88a33f021684bddd176647149;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he32cfd1eb3c27ab1829bc22c13c2ff2774e70ab62f099690ba23d0e27df3440aeb731abe23c9dfe1e356f343dd2675d5611fb4a5500a6e1dc4a53c077060721b371b524e09fa2034937dc10d937568585ae5da7dbd9b8d1802a15ef33a79243fb85c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd00d10be45830f51ffd819d8078926a23597bc5e75f3768b6fc12e58c28ad4537f6d561f76532fba6a8ba6422dbbd96143af7a68825e14ad5ba8c4b14a5e5a3e7c02825a609e493af94e8184a4f212fc88f3520ea7e404ebce1172982cfd75b68fb5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h809c20e544c8f6f4291db9a27175a7ecbffa6148fedf6980515a37cffbc261392a9c743f1a9081de74227f3aea06adf860536be8369c0d44e785c3518112b3c4da2dc645ac7a76e81a63a4f74186c23281c569c91abc03830d7563de2ecb0f75885b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cc3d104029830b81d9dbda3ad7669ee64df1ecbe5414f498cd108222b06d73870ef1bd6523247c043f79843587b29b26170bfd8ea3dfcb40a6b5153cfb76fe5bfbbc84036b89ad258944e7edb1da46dc9e4adbe4e60cf17d21206ce9b472dbb9986;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacf617b2b541d9be6e49196ae1b994b06c6f7adb9899ce652eb8bb6543201d99b6834bdfbfcf3dffbbae2c93bca215f1ae49860605a46d1ef133a0978bb851fc13a55d9c1bd5b2362f3ce1ddcbd539c6082fedd15ffed7226bc3b6aff04e16dfe6a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe90ada690e6671629f1ef8a56cf56d8706446e10bc5e4132f0983ffc6deb56b541843b281ce90c106e518aecefaa15cdbf1b1940e4a006703f56270ee88d9ccea3e04d539b78a2585172bd4728277093bc084a07810e3114e07d595cfb9d5426e74;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdcec5f317163d9ecca2857a0783fc7b2f96565df01027cd1312752b48a8c578bdcc0bb86316038b284a26a3132c105ac0a897b8d665942ba94f4e0ed48745aba1c77c1737c1494cea3cf6eaca24358a57e5e9930f1b25e9fb109688d3373766ca11;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9de7316faf8a0d33e0f3101a270138c030911460a0e08b1f7330d73fb8d983356fd21b47d4464ffca19d93c121cbed48dfd4e201186e880777356a2a53fe72dfe9ddec07a88a19e4849c232cca31e92382d9dfc620b423858adb687b70a7c60fa917;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92040c5f4f04a3cb27430fe0094fabf903ab7821872c5e012b8da3eb454817bd4835a46128a5dc6ff10bee909e15e91fa5311e83d873b7bd5a233d6b1971075fba4076460c82703fd4b344ceba8541c036e6a04e4cbd44c78a4ed19275e7296e7ae4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd33b4ab7f0c4b7530e63c41a97db503f379972afa019f660320f0c5204f8dfe2fd3616a1d456c197a4fea912ff158feca26396a21b1336afdd5a080ffd4f23618f0467817f274948071c107491e2370d812d4a61028ea9700e83885085e268cb402;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95bc538294c44fec0474126ef27e21e6052a2a363215ff43e8706e57eed5b867a288ce08193b26330655ebd84c40f4f51411787cb5a6bfa50b312c9bf612d054b2e38cc5cf9eafcf3041a0bcc2fc3c9accf7fc9de5149ad354f8356ab76f06974bbd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92a082adf7a35a34955dc6e84e74c1e05b7ad6d47ab58f5a49772bba449e06781fa11f03e3cd4e4fec44dc25fdcac5fe66572bd7760a4ccaf5c0a529a34b462d26345af3c068a998f0d78c92f5ad353f8847748e9f7f0dc3492c8f78a085a3739a4e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1cc04b41890ba237a10e3b8349075f1ccf11299e76b76072d3bfe7db4e78369238048607d9291e1ed7f47daebbc46c01ea7e5376c2ce84484679c40eeb7c9e2624acbb6cbd4c7bf295e855a057d804cc281b6ad470d2b110a44f8824680aa8c6d5e6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97f56491176c1efaa68bc5bad90ee8b0ea3a25250a86b3542dac7dd6c1faba3122a349d17da72bb2284240fd6369a63189e2cdd05271881c7d5ad642523b1c2172233b5fcf24d9d1334934c92ad39ff96fe0c13c49431567911596f04eb2ad0e9b70;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22886358e170fb069ba97f315dd839ad007d715e186d1ea46a389286b304bc7654bae437ddf6c3df334da318acbf06d2494096ec8736050bc59cb9ef2c43dc1296c0630c2e73ce9c8bc43d64ea1c2bb63e68bcd33bd91b4e34224ef066da28a30212;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61dba374b856a8614485e3bf67a3d54c3548afc965ea23f770c866fb0a5f4b1dd6c596690c664dcf6dfad16ee034517a7e04e8c5b1bdcc92f44ca686ba9c10b07a6a439d932f4434e25f0c62d99d6f005af0e9659a10e9144460d195673d08ae0c7c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ac3f6be568023abb02487e104d92c6b30b81859c1e28aed425156c16e5f03f43f04c8b3436e1cdf9321a959c98441930b7f06907bfb512b50808051f7c5886bf0b2d267816b5f36a5f60681e4ac7c434d67c2c10f8a0cbe5dd2d2820516ba3c3893;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74bf9c0276f0f91b44e0e2d1f5c0a6aa512199c8ee01e37e051127c7883d8cd05f816b4745f8fdbd9bba93d5866975d988cbc7b196b573f5ad6a0b08d9eca01e68923efe41b9b0e492930e5c7ef21a965752e7ca9826196f9de085234f025369b133;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h152853f70262409d4e048e74b7caefe8b9171840203e1660710ab765e9d843647fe07434d97859f01f347fbff68cc9074a8ab2bb8baa42aac4e2a0f7f39f4f26a504abfac9bae734b0b0ee66feb1aa476b88b27ac5c223ebd4642d625ab07ef08290;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab32056287893eb5f1cedf90fbd2bfa63d50782492d1c5cffe0bcae70b580f1b6a3535181b304342d35e9195251bc066eca4480437a3359c43e2f64f7e4eccfef59e50942b734475e77d80afcd94d589d398d1729b4a2246e755a08b495e181f6f26;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d23064908c8d8bdcf353bf0d7795b496c060640363d169c4fbb1cd5554a8d4ebfac1e2eb0777caa5c5e54faa08198ef34aa9caa7d7724725a51b9deb4f455cfdaa010f7913c660e8a3a392e4e4d68c82d863baa6a4623320105af0b49329935eb3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8b7ea109594d936fcc2144c6cf6b423ea08c57c032052b7a2ba24d4a893d1dd967b399d8a17754d9b67c7f0f50842590ecb20d33107c60f545b0937a8bea80266566ce12e3e58afb104c06f35d3183941cb98cc0a0fa8ea0d7c1f497be2c2d126f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb5e0341b79206e5d45aa8ae49dccbe7ef960a4f1871817229e8603f20a6a3a2b12de301742d1c2565226f0eba956205033d97d7de335ae6e0f17ceaf283804dd1401bf29ed9c1e5b791d63e4a31b6220262c0fa35706b563db8c7dd0c82c2f60c61;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65ebc940b2db0be2866a3a03c6232d36255adc811977668cfcd46fef548e832587b9c925afd2dd807cf15e09ce9b6d6012cf9e15e1c71f57df281031927f0368deb351e722de6358125466b00105d99a9d23919c00fde660ae6aa9ea1e169b61bb4f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc303df935a9ecd2a105bedcafd7f1b3ba4b1b5d91873f1e26e42aff633ddf62f263dbc0a1d2cfcf8f0464d2cddc5636da8a7923ddb6c2cd82d24da8a60e6e3b29c539df23636e391b8c81a049d7f1f0da951709b197500aa93cc934e22408bbbd90c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b8b2097cd33382f9a27f5c228851a819890bddfeca52ad23aac237914c0c4a9dfb59f99fcdfd9004d64468de05599e0e94d50590c5c498b71fcfcc34fafe31985d3bf4f9293839c7b8611167211ac18c44870e8a55727733c6953e371dff7e676a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45c96ad693a98872d69d0839d4adad3ef02407ccbb3e7b76e18173ae73cb39b15958d0ea1771079d9638dabec570d370ed2edd1942a5331d7c6183de45d164319b8b29e74896b449fe8be1468fdf595f5465d40d731041dcb10785c7a311a342da97;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fb45a76725926fcac2f130bfc380873e543e9fdda5668b5052ac4ebf203f74582ae1a3fc97b0a97128b33bb2f255b0666a6b3ad06869c8f6ce4394e353bbc4c55fedc61b9eac595f2d628c508b802a8b64c3755f244aed99f0454e79f745163d2f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22086ed1004f6a8fe5cd7de2e9009eab1e00c59affffda3b150deb3b9d151fccc960e4b076f8421135902fa441efa820655e47de6dc8a32ef6e1e7c73be353a4e10d9bbb84bc4e32bda58ee42eaa3bbad294b2ef2c2c5777c71082520526b4086949;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35b226ee6d35daeb58e059fe2d034c187889abf9fe64dc8989da2dffa584e94e17a221cc4a4aca27d861f3af5b9518c6b1bd8029b162c147e001d39c04ad5a698d416c265dd908e56501cda953fa6e6b1876de7d274401fc8703419ad4611b680257;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8248a7860dcbca5e0ec623449a36ec77f2a461cfb5d8ebc2dfe7d35faa82a9d2b9223eb8e392628ed6039989def9146f0b951d7e08d0c1d719c26bc540362c038c2dfa9fdcabcff86608f93915d2b8f4d514b4e63a683e1657f34cc7fac1ae743e8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he76ffc89f53c35691a69c1d9edbd2f47166d555c21616bf5e267369ef8b751c5c6816cfe00c34d52c62c6c3f2105847de9cd01fa1c37ef5d4fbacf3bdf3c7ccafdb6426ed64c9f2d220389efb105afed134556fd4a07fd2a303e948c22dc8141973f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h323a4f2004a61f2dbf6fe30b34d96a7e3e2fec4f4f013a3c4c81f4515e50217e7436cbd28ee74850eb295cedc09917e543ed2eed6d9072a7dda3fb939bdd22a35256a31971329a0812c57a6941867a6ad987ea9ce40afe909795a5d7270daa9767b6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5c8683cc0d118dfadf7fc26f60a1c75aa37e924ae8421a26b711499a5ca606cb6ca4a09e0fe70f99dce9fc331cc694ea11092cfff1381c57d76b9a411881d1759013280e1e649a8501e857784af29c9c6f475ca2cd7ec357b001491d1231ed88c78;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec08b8d1d6edc0091781f6e2ae85b54b16de5c4d60f0a13ceceecbd5bc60ff2023f5abcc9b7610e1eb2cfa10a3118051f5a277a7a129ef8206f7720046f2289a0ee810e4ff81755e9e23fdf8ee6646ee4b3f49923bb11ba142e935f4b5ec24052ff8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bda3c9d6448326ec86ba347d27ac5a59d14ba45719cb89e78c507501a574c500cc3eb9ff0a94f51a982288f432ed2f419096a8856e2ffd06f791365b8ba652ee9c25114247ac21890bb140ccb2c52535be121d9189364fbe72c0e83f2c700bf799d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d8bfd6770f1a2084cbc5114e874da8acdf62ed7dc1760148235c7f98e4dafdb47ecb646907d345ed04324b3e8f43fce783c344363dfffa2028e6eeb87d1c4d544546fffc30962985e9cc6da562adcfd60b3e362ff49f2fb2ed0a1632129dba3ee94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4bd619d747524cd2265530009c4eba44ef74d91c047d69b6cff58b2d38604761afb37c79908e3d48b3bd17ae4960e701f97606010b4de1472d4c79f69ad7030d740106e7d094aa12db0cc9befa85249c2c758152d76b1e2d31541e71ea805dd94ea7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51d5e80e804eb38400f28543878e591fa1984c0f2fe38a87cac977001a00031c3ed23a49142adbe980c56ad0f49e608ff2becb16997db94a8dfec45b0c3849a423c16740980870aa901500abec56f60a06d7fa4f31025bb997e3ef6b8c1a821b1bab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd30b3ad1fb1e135f42e23f839cf221a0c2d9d447859a26b47b702587bad7c772722ea471e5ef9d2d32d662f39cf66c5b49ac20ef5dc194826f3b83f4410fcfb31d13b78f9615ee457248f885c83fa982357643468286d791766b7900f0f17d2b9b15;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc150966fda9e3a65c91eaff1469439e2d0d08426db494e017b4f3dd813540bd3700e7051ee5338dc6a161a646843ebb0f4fac6e0026df5f5b1aa91087efa2ed9a78199c8d9eb62e6c753c6df24047fe246650e7d09784ef6c91051a8af15ee7e0adf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf881b74a34d16a5fe87c1537b211511801332e1c69bcfeba015fb3e2d4e93e94b71cc6c94fce09783e4aa422e425bae94019ea4a0128d9e008a3d6fe663acf8b0afca274201c2668cd9279df7d5ccd8180560017f36665f69f4e020427ed669cbc72;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77d008f4c80874a3e291f56656546c22e0d85737f191d79b9162a85777461e7b1fdb550d6c297e51d692b44fb6800631ce482139f16d9c945e562d33e194c4aab9bde1695ac9ee86ed29d7a3a6a14c930d9e9de65718de31f490eb8359a15a6a6f1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43e4eea9e4f3e5d861963bacb2c2dc933e962e0a454ed960426b55d72ef40c111042d04000292dccc354f5a4496bffa039ee86b49a47e7480681d07aa0bfa264214621fa99671b40542ca727c789754f0ede69efb85801454c780c33d2c7a18ad651;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd1dcabbd5873b13b127b021ac31e70fea420a02c8cfc96a7d68525f090424bafa94b318b98cc6d7a1bba66e12f903408cb8391df7fec4e960a380ecf93df2fbfcecf33b39ad1e7d81636378a68f3a991ee2cbdb696e831e9adc88315add3af1ed3e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5784de55642836aea0ab7f77bd725a6b0efcf72125abba83c24f1ec2aed1691efee37fae4d0e1b888bdcf6d9ea5da79519ca73f31513501b401918baa92ebad8eb56d0b0b366156d37ad18d1feb9f03fda9872c709b7174e261922a60f670213dcbf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf947d3190ca680c4d30c230b7158fa7c75993709e6ec98778f0d4cb72b98baee39ad04035ada97731a29b519dc61abd80e2e431c85da05d049f3f8ac164165164ec6f7b2297fad5384c628e3025254211acf43cd279048576a0a0b5b1f74bce7911a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1aa66b395f45ce4106487de1a86a6f8f4147d38fc7691d2776d3ab484d4526f135a5d7e08c0c9c796ab0c674381c3b866652fbecdc1ae96494fe15143647f6f2dd647e1d32a5cc30a8b15c0d030b2d39545afe6fa2817b983fee615781889619d0e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bf6e765f1cca0eddc4fd3b75ebe2b6b1c6419c0e0db0e8d2eee0de3da27d2b1b494779606744ee7731b19a553364f00e9fe8f4d4d07df321697a051c6e09495dca49d2fb9ff897278506b37eebd953e40816c8be7924d5863e566f7598a0ce58ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fd2c895bf69b3c54c25ff864d260dbf513c5649741173d687529b063a92e19e254166348eb5a149adf3be619aec49cc50cbdad7ba86613f523715826355435207fc989587f19b1faf7ba01672608c4b3cbf114e60e136c0766b73ad337c1bffcfd7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14cf266b6865d48416b593fd1192fef28d7e17ed2efa9c29fba5b81cbbc4518212bfb944fba13117f71237ce8188caaefba60c4d30cf43b107889daee77314deeea4bcd363b0d003645f3553f649e24f29dfbdcc7c0ec89f14c7e52a502123634437;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc51fb841e5c3b29717b1bd39e51cf2a1f381e5f57c66d481bcfc7d1476e62fab7b086ac882abea1941701c1a8828252720c685e43722aa638013bd7905460cdf3a3b48dba128604085b451ea1172f6c39e7fe26566e3e062a6fa73d8c0eaec78835d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27dbca212b5fa5b7f5d496eb1b7439f70d533c80ac6047920b5aaf8b8170292d4e0a864da1726a340ad9f5642d6a8e87112f13ae1aa2b4d910f9fac613374d8a9dad10e32c5b5f687072144cdbc376d43efbc769a2e55d76d4cfe239ecbf74216a84;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h855b051bd60a53b5394c34e70f00805fd45c6cb53904f42030897f9d4e51c583fb0c224dcd1ef85d2cddc330051e9d7a20a17b143f0bee495085c978caf314a3e6edc09ae96bc0ddb27620765d65697bf2f3f88e57cab936b401a23309e10b812773;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbebdb012b58fb6c51968f780c7aebfd48f174d3beafbb42a2bf710cf83a870e54a1ebb39c113cb385ac45193f84e400527031f506cb529097722a96ef64446a050c3a17f294f510f02e2cb22df658812c091e7733329ca5b02e3a18af80800ab51ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c0d73dbb3793579930875fa25d2d0c3efb7fd67e39fb29280bc9fe3b17fc8c834bf712dd1f822cee21ea09a0033d8cb93675b4c01d4f21bb0cae2eb35aca50df0cbc46678904c8161412028b7f90ff3d4109f87c1b9d4b85f6d8b80287f8176b093;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76104f42212a94a207147df6e7cf61024ccd6a108d00eeb553ed47f054f6e8f2e92439e1540284918e7189793a5fc62e8ddf1df9f230d68de963b9d5175bcf95677d80a39df77e0d1f810476353a2250bfa5cada1177e086ab05865f2ecb29eef89b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff4b71e820268495a938439fd758f889a6a248271dbebb5f57e8dae5201b7f440dca534685a9953b39614bb90977e23ff05ca7e833d2d78ede5e009bd760f76e70cf1fe8fa600c54464c5fe4eaefd726012f5c6557e64ce6ee4891af69e58270b324;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h715f3f3f03b3308787bbd75075f59d290d55b78990305d6a5f28d967f5ad8d8da2ae22c7117456a3fd3abc32898c046ccf91e3018f636aee719414115b25ade61e8dff5f661c9f227bc2f6b44818c3839c4e7f30fc39496ab83a56a29314f3d57c5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6e2a02f6911e98e96c0304fa3e18555e896fc1f99fb95539fad769a67557241811b283f082f750ab7b9fa57dd23bae17a13875bb74c1961570660b0491df7dcef479e1d77ac90e1a200fb874f2b2bddd1750ec6416a1edff9b812def31ea22eaaab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc280205bca63ed26c0b88a7dfc3a94ac445e1a6c33e563f70dce742eae0ba6b4f1976954141120a168e46633177c3c195a23ec89deaab8b6688a0acfa80fd640ba9080c49441f107b218bd14ce448901e5fdf0ea47e07c913c0056cbf27883eb24d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcddc208a66b973a064446f531f01138212ed059dcb9efc634d7af5536f8926f515272fc7c2a5b5c359cca0ac9d498a2a1aaa513a7f51355222e8eeb2d86fccba0f54c60753771acf94cab16d76aecbb163b34f7be7cc0149e651c73baee2925d4a6b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b2a7e8eaa8d5288afa271d5f7af9dae61f5b7ec7f87797696087c38b27187412db9d4aad364f63a3e8c71a61dfd83cb46bce570c23c350173ae9d1bb5258989f573ccb3c15a25024e3487eff7afb11fe025002df9ca12870256d4a7743cb43bc732;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d1003fd946d80834ea17f50a6327aa348118cadea5b39b939c00d4f6a66414580b33fe9a8be320b515edb19b68561d366e92bc165ed46c70f57ca58f52287b192c343e3cf6ba44ab1f8b720ac84f3174ca53794820ac1c98daa8ab199a824ce0f1c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d7718eb50ebcd4a13829a2cd124a196c2df4e3e5d5d80eeb72704ab124266148f9c82161cb017b76c2d9c14327317972c8acb1203fcf0158faa5fa08f43333ce9025a1d4ca60c658b5583a304db7832db8d8cbafa9178215d65f4565557eed37e36;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha379fab0dbbd908ac38a52b34852f9b096a57f82ad223d47bfc83128cfb4d8b3c5d55703bf6857f0fa9335651916f9ae6dc1f368ee53546a8e8a5ef81f0b97f6b5ebb5d7b48bbc3df294dcfaa7a8c99e805ddcf67e61a825d603df63d7933b13b702;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc33490abd0c6a1d9ef1f96ebf7411e2ceb0f569f83e7b2e1e5e53e20adda3b8a6f0e9f49ae48829eca416774c3a629cc8e1653a05461b6e165e3c21519d9211302a712778a9701c4a1664fbd722ad55ac41251ef3ca750715f5fd00e3c60da84dfc4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc571832359d81917e4cc9c1843a59ba586fc5a911b0c5166503e757b0cbbbf99239922a72af1972eafd5e82222ebf36fa6025da4c70343d73849b5eac49cc888255549b0a36a4e3a4cfce7f9447b58bcf3449408c3e367c037ae9da882b96f12e99a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h895f2d6cc7ca78c69d2b34dea5b6251b8d0393925c36efd813fa4fbb7309e00cc026bfb4c2b9a86779e8a9911aeb72f0d538e465b8bce76755d73969acb67f3345851d35a054aa4e97c2cb1a0ceacfc5293b9344c4a41f8eda23cfb9e8e3a29aecf8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h882c1b4c6bcd7f0d2ce32500d8a97c4c7852497a05a7e76d7696d436480204699a40a8a148002741d4748ecbcc99367f6a21e5a19e344845174700b5d3e4915aaa25f79c736e3e64eb9255454be63eef3a0c6296a498f67147d35d712b1244b501b4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9dca30c7fb16c4e33feb7aec1d5da3284a5dc47a5a501cd99cc7fac24028ccbb6bc9f78ccbab72f74babdb91594ec0c74c2c40ca1556d8d6ef1a14243535600b4a7c064ea857cdafb0633535e35c249f87897813bd6555ad73ef523ed41df2003d54;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22643f1cd813c0a16b6fdeff50d1bc51bac866c89e857633d9c7eab45304d5f66507186644694bd664876d92e78f6c1bd1cf9b686475ffee475fcbf65dbcce56453cf03d1a0eb47af040361eaeb973746aaa24abe7dab61d7535dbb4562b4f2cc396;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c1d1e4628b1ea4c46c1c651fd76a6e3850f6d4a7ca7911de20d9b9cab0860be479837f2b3d10b1c50c6e7bd5b95047ad4989d473712b4d9c3fea23fc4013314b3c4f6ef0b8d402bd3246c9c3c7dfce4f88882d80ba7d9d2c1fa3e34137c79a3d39c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b0294eddfa03a24f4c766dbba1675daf8df56295b3f27cc1f47626ff16361afa284b93bcc37e6d556600828f75f0d9e94e49d39cd96853970400f943ff107eb8f0eb53f7b708fbbc11b36d1b70ac6bacc28bfa17faec0d7a167b8b1970ddf71839;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12ae12d1bc1c9ebc8302f68093a8ddb6b31d2abbe1de6ced6929f40a78051c4449b38271538bc3e1c9c3e9e8567a4d4c61160b07ac1c08de2a95abc5424700c8aaab9e1630e8dea92287e658483c68c305a73af05aa025ba9222cf365d30efb1e61;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cb05976b372ebe03f58246260e6c15f96554ad88b252b1bfda09e910825d6e464d5fb2dceb301e93a42cc2a264ecc4c9059929d6e4e2208c425f1451dd76175a6b9e53794a9e74a2abbf48c78da9075dd13ed0d4a23673769a0f333a280137ab10f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13b257149f316b48d699c4298fde0fb065739a18e4edf3079c2de97c4f58b3ad22b1ddfefd83f622744f5cbeec86edd7fa9642b2d7d95da1d0f547bbfc896352e35f0bf721b1d99ff947572be74b139a70b83b64e8e92974d9f2361f9bd70d02f7b5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b18780f2599277aa58617ae144e17e7728d29d6028076d8b6764ad27d124cc81be9d75de0111b941d8c31144d987034d4798962f5448b0c4b4a183811fc11196b0815ed27f44d97df19794aaf0653c8b136acc5336b7021fb3699551bcb0a90e21e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heaa99d94e2ee7da8cd280426f579269581a70512292c8fc5faa6218af2258cd84fd5eb85868a0731008c5ee4fe9a0a663b8cc9f950f33fb1cbafb98fb130317e82d808796899edd4f5ae33c2426673f1488134dcb0021436222342893a19daa20041;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7be28a1d92b6fe2a8254b2c11c898afb19d84f3128eb44654c0c3756718eafe90b2a0fed3b961af0d35890ab48aa9d77666e1a2c0935ae04494be19389ebdd0b47c636d7504907032d195faac7d1249847c9ed85629afebf8f42115d93e3754f681b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3c9d7fb97e4bc1caab77b508c7026778a3183d25023b39c038f5d6b498b7bc896a485c55bfd60af1b7aa7e4544ca70fbb0313605a327b90b10c66a7cc80d85fb133ad96605f9b9626b0df96c8f1cb809e28d5e2677175cfb6fdfee825061798092e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8359348d5872b22fc2abe73f26cc9a3e4460ce6fafd61f2b791024fbbb4a03c528a31f786d73185731bd40a78548e1c5100734be7ff768c9e114635fbd039035dd0a0796e2927d0b638579f0003382c1ede5cb67f60509da6e036df3f2bba3b9541;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf113cc6972bce409c4d38bb4033caada4d429c0cf2f76ff5e758a7f95232cfcc6eb02e94096b8465f81a42c4e5149a53f2d59fb0ceb0452ffeabb29b1ad58f2c91d7ead98c13ae8b362edbad28bcb696802c9b8744820574135799c49ae5fe5e3121;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd592a44c732980141a446f924bdc9a9015e1f97b332aaa441040dd18999dd140ec2f03ee35573ee6aea06d44b700fb98c239041933347429a8862d8ca6d46e80049ed73cd2507e4adf7320471e8aad03796bf2a379b08e963987b017a9ccb5b7f982;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93870417ef880d943028f342ba86fbfee1516424419068e86c6024d07fc72f55c1d512816cd06ab4904670641cb72ac267177b6bece2ccf58b1d877ca1bd2034a3ea8010a6840ff9d1211560bffcbdea672f29e6463a4f6f034dad3699acca5f4370;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3026397b326836eb0560125f0cddb7eb7a9c26773bcdcdca8098afc34894296c2edb45ce84ac3c790362114ef8af6acad91691f1834db0b662bd085940358c8faf060445a83219ca0d5a01417f70e75885fe4bfb2848bb8515d24872c3006f444ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65226c356e771dba0c27781d73ddc4e47b48b556a74d96984bfc284c3464bafa2eb5dbdd40ebbbbd7691a41c64a9a4cb003b7c74f089f9d4fdd63adb0df918680ea4b046754a5cd02fa7538dff250931b8a1ff042331c8c83f7724387bd2aebc306d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3109600303525d2e8d9eb99bedc5360355a400e824dfd374513c314963f394bb440872dbd930cd9f676de3e897233b8a83191f67810a81370f3cdf446181ff7cdcd20e466d17a0be8019d26cb21099063f999d9d4d9148b5c5f5c2c0e18d2e37baa9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c070ba49a9374e0848d22a53acfa0a4ab082fb2219ff287a448a45edc45d6296c35267f12f130af27a9cce07de80cab3ce073ad06c892b37a7e993af012530da550112eeb7d8ff805df56efa2e787470964b6e22e57b508a48de3f10f45aed4ca63;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc106a62ed375eec82b60407f4e3ee6f6195b06aa37122807af6b8088a458037b567c98104011eff30938e3396f1cbd7ecca5f1cd051e7da0f36451548f1c8debfaa2e905325c11419c995f9072c6e6719bfefd325c78a53177f8c2738f97c7cc0cd3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h946d1296f34749e18c5b090a2b3a4a43c5e40294970e22f9906b43eb38845bb47d6d425f3da78f1acfecbe9cfc4dd5d2ddf16c59c3c156d9341a2455c6bca0dbf45bcf6904c4070d10fcc70c8fe0c010f3463a4b025668d5926669cc335dd8441b24;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55f4251bd7bc9ac98bc06ea9340f641caf215a1c13ee825fd5f3f0ec760a6fe67fe6382a61fc859bcabd5bfeb49a59ef4022b9d27c60e6323797fde17c2650d657767d3209e8ef1d171b92443076282791e0a986122b2463215f74dd8957b2f681ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e17fc222284417485dada64915054ac329ccdfb91cb16ab8ccf6d9ada18be2d91ac51234e5f83ed3330c340602313b87f882a100c93f02ae62fabf512b4e8e39d8bee56339b63175e80dee445a20b35231f2953041115ec1659ea45d6877c224b38;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha726993602f2bf3e72db9e13c210043b1b32256e6d8e8928848153ff109cb71579298a4741bc50f733a93c81cb15b7cf49658626bb24e04be443c140edd12198fabf939bb9554e59cf0a845f7c746d21ce35050988f2600ed5c5c9bd9440b8e08230;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0a4a9aa3cff09544f1cac0e9ead4055f16116444bd7720366c838cbfa7f1e08a78afbbaa1e706c4c78518e93818bd41de5c5bda1047a7e85914ca3360ddfa2a281db53528071e648258a50c9104c161cba6d955c8f96eb9a1e5f8458be406f4a154;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3a1e61ed94407c0e7ca969a200b95d22b81cd5d19349a4cea5a13a193fc43c061d62efd12f2396409abde8c2cb881660ee3102c34cfe05e577d9677f185e4cf3a1bef2878b00b36c6fff40cb91d18a2ce4c99365dee872ceabf69f255b14177ef72;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8f9436431c56367a54d81d9445747a47e4c7ea5491dbb733799ec0cc5c4d4c495ca8bbab7bea35829061e2c3914da598f22a79535a8b03a3fdf13ae27e59dc9dc6f375fb366778128d1c6b6216814575d5e0b86e848dc97d103c261148b4f45611d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82b9595c0c516f22fb8166d860c7ec39c1b0dc0313e8e809bb72f115b1f5ef4a267fb5c4a59eb09728f5a0e8e2edd8fcafef7335fbb55b7e6201fe02daf2580e212c2adcd3f0d1574332a6efbcae790c7b8178100804af1c07cda136833f60c4bda1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a4746e7b6828074979862d1f2e5c94557568d9a9f8f0e4962f122dcaa237a07deefc173ef5e29e42a98926671e4566f97eec46a8b587311f850a91af1271ae67542b19d294787a7a5e033ff8792dee687b5cc5234603a9ba7a4740b2a180915465;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d9c16b81faa23e68b4b40698fd531ffb79d73bd77fbc4a3c90dbfebffae5dde85b831d0968444ca023c374417174d2862d336b95e82a2677347d24d3f095bdd0fab1baaad2ec46eaa922a835decabf1548a4f69eab7eabf6c531d5067f10402628c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0cc39b676a1b65b5e0d0f64015ecb672cd0e3dc9cc95601e34f47298f3aeff991e308c40455ea4fd153da8cd80bc621fde2fba59c028e3bc116e29de297759c26a622b9f4d46e0693901c717c16fc18fdf61b624071c0c20a93bf904673de755278;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42557f63ea6b4f84ffd1fee38f315f3c7b6e356431f304276dc302b7d4f146dde683e0c2f11d90fcbd4ebaf959b40e2474ae60cb746b8fa9f97a89f55b4f86a4e8c06402f9a2648bbdff44f476b0fb91c04b89ec820b61417be3406491cb07fe4397;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94ed7b34312c56e84d21e8209b14357e8db5a106254262b7f999e7c398e62ec90e1f2ba43b5e6d00b6c6dbc105bfbddbaee9f9cb1d216ea1c3e2d15048c255e0f9f635cfe648abc6d33a74e7e46bb0f03b664273e009abc0167ae64aef72aa32fafa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab1af2542045d986b05e001d14b3276a05df70cc7c828df51209f6c33db29fd24d6e90a148cadecfacde049773812c34e74f7b2b3b2b2099dae279dada8832bd8d1c71513eb19a3e652377d433b15bdcc8898f7e3901b4bcb8afce677e462795c8ea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0d6cb3e664cf0508ed96b76d125ab6d025eb484653cfac2cab6da2b39bd4ca94518d7bce67853442e6886fb0b9e993ac8bae7d60235b184a6da4b731d2405b8cd2d200e0a241e3a8f2efd8a7c4c5257691d18ae7271920c7046296b03fb9191aa38;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h761f510cbabc63b8eb3dc3230a2778c592e1cbc5697322b0ce9204d6aac0cb33659c4cfe7c3aefc9baa0a0c5729e3f5f9be54b9e070f96697eb44c0861cb57e8e23a7fb186c1a7eea406df91bc8479ae059f417a30f5ad045f6af781b3af8a0fe3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f0987506a480d7e9bed88c17fe6d594a53d9f54c32e8365fb0eb965d412159ac0ecae2ba9d062f5dd2cd86770573a1cbbe9155cb33f7129ed13f3d9b185492a7282bda15878b115a8489866209c404c929aafc19b49b0f33b0a1bd515dce8d84e70;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84e2d18339aa163e0bb7cb7ec4297dd0449533747da2864de455aaaa235bd1f252bbad503fb09cdcbbe8c698057abc32f56d1d8bb9bfe8dc66f75ea7c821a8891a23adfba2a5e5d718656fff42a78eebb346d40d6e026320f90085569aae70322ad6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d8a777f4f131aadb1299a1c03e4c5351b3fced7235cc39bc273262473f683e610f83c6981966bc806b3f7983f7a433f1588b542d4921fbd4d22907995ca487df5bc820662f31448de552029c892794d3be4ffa7ac95c334a6c5e143f86807eee7b8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1c24dc5b1f9ddd96f4bbb15f54c0c9ed52dd7e7b1c218ce218844cf060f239af3e79daf00cfcb1529a43ef6fa3f4d2e993d4d03b7a103ea14355e4eac507d5ffae632c3fd2d0fa4ad2f7465fbf11d3c16381c0fc824a2c00e291295f86976ca48d4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ee059f6ce24d1b0a350626593cc35e3a14b3fd79e28a34e97766da88ad4c7f36f3a37b4f3df04acdc76fb3e92b811c59611c2a52c2ae51f62178570dfe392bd307889a6c6e50d001a54c6e987d4ba30a04cac9f2c46bf33c3acabd7a686f07f06d4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb68f1e3d0150acd369493576227c6da6952e08ef9b38445b655fc7649e57743bf6fd553cb62040389ba103e66c73c55309b76a59c334c3e146aad5ef7e3d3aaf64c1c5154a694a846da0fb13e48fb5d37ebe1d1f936e785a80c66e7eab83c081759;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0f9376b046cefd5886bb12d5ff246f04c78ec4a4c201ed5dced513e795f6c3981aaee76c62f33fb6a6a1d17261895628a241ec298280cb163950c7a16499492372b0a8d3222853d180cfdf9219a24f4581b419f77900ce2c6a50bafab6cc3d58477;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa342a4eee705ad9a3d31c772716e771c4329b12eb63bcf9abf6b6c3b7584fe3a4a8e8c68745ac1bf748533600fda690fdae503bf201212d81a094ca0ecafe3dadf4afe266d2a108f57b565dd1465a30f47a3ed4fec9022d4bb5b6c717139a60334b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4dba7fccb0a09f2c8e4154e48bc4d8cba4e61e7022e07a3e87c3d35bc6f2ba7c47287be21841d6ce091a7280673470e9212b7f2eb5b594be53ca624bf6d40da0bb2dec985ec70acdb9193aa4642df6160168d28608c7a6bc8f2d565bddf65730c706;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha69650746add4662039a7c956eaec3225cc86c38bc86d5343fd68cb5a772b0891f851a54c7470990c272cbc558749c7f69f1540b07e43a88cbd852b70e8f4837bce0ab5f4b20caf907c0ffb3737b0fb918c9fb3fac5b5b85852798186d578fc4bf59;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b12474d08a689bc2519cf3a4b04a4c3189fdafe72f0474a346a08b9d0a697d47cacf7964e963ac90649d4ecde3f8a5eabad8f63502dd6b28bf5981a5f4d64ef1fa7854fe3824176d32b7bfb6a0601f75969555fe89baed3de8c0d2abe09547d32;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5c26b6cc9cd9f6b25a5c36a3b126d9dea6f766e66a8078a91e934f67fb1eb05bd5b24d6c47317b307093b2e7af0e167b954fdb539be938944715098ba574019ffb0fad3639d3dac94c1cbd4f5671a0bf146ba109e615bb6a77980ede6308e5433ba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83ba10d3cea496eba164543e2bb71762cb7ecf6296b0aed49b37591bc22fec0bcdc108b8e10bc3de54582206d312a23cd28101fd09ec3e50cad19ebb4f6d7618fca0e55437d94b33d41c647cf68c765bc38c1f855aabc5640307dfbe6beec4188660;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3d08540dd7ef08e7fb79c37b61b852c9057e0c11a61a4719d3eba922c42260e8a762e393a34d4ad9be770dd211f69588cd45af55508c4e256ab9d108d6eba8de2e3a111c6ce6e6e074bcd00798283e46c5add455555445e348632c8f46b209ba4a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4bc8ceab502fc86dbca24e3d9adbd70dbb279ef7813105f952b8aff5a3eab0840a88a2d0e3fb673542616c6e109b1a2d61f704ca2697cf07110cd2b0141c324840da68f36cbe97e799862b7be5aa79eda168b727995b0c71b1aba222d28f198cde4c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h752662a52ed3b2c6f0ce474f60dd3d88866ada1480dd1b524cdcd2b3ed97ccde8fca37003370a7d0506a854ff902b829262f69e596174ea9c3d1c1e50992da83d80976b163180c63913e25b24809dca003d1f15b8c405f56b045079ef7c83b30c116;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4122cf9681681e40b2d0405c86221d8225cea1b474a995d60aaadecc8b9047eec467eb1773e42d8eab194c4c7edd6c0664ca5634c04e8a93b68cdd90a13ddcde3dc0130b016643012c224c6ce0733872db62732380eacbab8516fd0ed1fba32d146e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h448f82452ecc39dccae6408685e57348d40c024edf4a76ade89d416a45cfd59047498993a46372a2c5705b6c21a3b4a0fbe33ed707add2120009121c51280c1c08e267e4aca029dfa5cd2e1eaa3efa092e9ed58499cb712b8f8ae5aabb72db2d6074;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3022bac236bc33331600d27e9b4704c4d91c24ffae22b0c271d8797faac23ee8630d8f722c8b61b34a64dca7aeca0d6faa5ce13affec2606c5b9f1a5604fe8c49a12380a4d8395066b6cc3a0db43f7c72f5ec9ba1a9d6e832f4aeade8dcb7f84bfb4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59fdde64e47a90f5d34d8ed4a59f082c94bea9ed563e3e1752cd886ea104acab571870a4d5d23522b4ac82e145862b1a395b5ce5a43de826a53a200caf17b066c366cad150b161c0ab70f449aeaca809ddccc3ae29d4faa90d3c974f4b9f38f7767;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5686423b30ba9cffee33b7313b9a5f3f911bc91b0d458e1821909319ab38aec013b8928f2d0fc25a6789cb974ed48dcdda1a8769575599094d226f86f1fd5af371828e539ea1347df06ce30ce9934246f26acc4243aa0b1e512aee21600a3c527a79;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecd59af820400c7b5e4235b2581ebb50fa6ddf75dffbb63977e9de1736cef0d0e12c0ec97f92e543dd8977380512686cd1bba5a6513abbe0d4c1bb270b2dda3104cd5f2f69b627d30b718335521da5f348853dd5b72bb31122491970a644c44b9748;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc745b75c39b2d8509d692817a5474bb83fab80f456b9d1f6a78ee67c09eb6c0f19d0adf973c3dab8a940ac568211f122e5117e915359bcc7e9da8fb56116175a6c43f87243829f6ba94c8e52fc43be482f18c25599b62d1d968c01f331f08c12dbda;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44e9792c3e4e0974d75731ad5559a1a509f36b5a664ad1254b5e0f5d4ebe5156b156c354857e646bd717756a357eaa38ec3e527a93e627878765e3dcf073f3b3928c58f16772045d49ae6db7f0b3be692b798b86901dc6cb08d7dc6f216d30c9f9b7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3926e31522c86b2008d9257854a818ef03463e687be4f50ff8465440c3c46fbb3d6eb0cdc442912acf58ba030484c18accf29a01c1b87652ae4fcb8b274d4ae11773b1c50c00e834aa131e8b1490675052336729441323b4b7d67fe8bf78edd975f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e5381f429a0b223505939be20ed12694880d36762f7c7a8dea7f7007a1f33bcd12e23dd026be458ef813d988f4b68e4906f6067c8ccfc34ecf4bc3068b31f824b62d331413e9ec03f8141f687c51def3c41fb62fba985413bf8a6ff15cf080f178e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc11147badfc5e35745e30a3439d99261a5e9ab35ce731607f3cc838deb2dd3e2e93dc9d6f3ed20269823feb11fb0e24eb714972de954db32e1f05236c0c1ae6510b2a216ab7b8fbfd2c4b1868b5be53ed93a60fbda756184adef1a488c91d588ecd0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had6107c0bb6019d051c764aee655c50168686af875644a52ef14715cdd13f49bc1efcb109c85774718a12981f21c79d0a96bfcb2f3316cfa3d718c66f1c7953b5dc5b6d169201c3880a7c2671a804f8b311d59e5022ecd3880be441c03b3dddb63b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he578886535cae552d4a4aeb348c84ac4a9c469d14a1f8fdd468efd89c9e5ee26e60a71cc70ae028182a6df49c33a098c310632f224061ad6328b15bb132c12d70019b2b5cbbb58457b803aa7f84a9abda0dfb726daa51634ab5624956b495975b767;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d0fcbf3453544c85f8ce569af807e9d7f1c2d44eebdea20f6328bf9d3632243171dd0e9d9024591f54116b0fb1eeb28d1f35f768e9a8b50da3b104659f31332fb736a8268b1b704163aa8ca57853a286141b92d9a3771a988afa55e356b0c2369b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h272a7cd1c8f40b86981b2ce25f796da23dacfe847f8e5b41df3b133f5923b518978acb57aebafd26c624be066298c497f5b0d5d46bc649334bbb74546da17e07b1f35f75bc51d83005c2292e4aa16153499218f667e43fa33060819a4ca646c1b0c5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe51f0e8005cb1541c881c4d3b78e1b3f8981a1c9b6ebc123bc7f9ecca3dfed332406ec1a54ba7f33475700bb36309bf727a7dd5509fde494b01f249ec8d609905ba3e8078ded6169a10bc43d7b9854229f1983f891e5e4665102ea6a13addf6325b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dab683d70ff71373a2bcab9881fd54fa3ec9671260b4367873cc5e85e4e85dfb40fdf14bc03e439d3859b14cc70055a7dcb8a47bda84d3717a75e00a41797f0427b425ee6de8973e93bf2dfa919198527f6e81bdbbed414743ca0ac0ff5f6c86720;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18bfb175a6bc45c12e2291f8bfdd693ec07b783363c35ca1fd337522b399beae7e625c4845ceadbb7cdb10405e9b31cbf031544ea9954f930a318134e77e20b77a92f86f0b47f0bb23903c1a0e292c6a8be83980439688ef64f134d1d2351ba581b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94883d8a43ec846108fb1ac79c00f5facf56a291ecf4fb5d967a1bca75e0d6f5612601857418d694b9b8942d2d0766c771315c42917993e2f47f34641ae1891b9d8b43724e91ba60cba76ccfd20d081160222cc725b77c1aee17525bed0e46e1f0f5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f6dd18f6dc2bddb07829b61c1441f326f6513f75e9951e6a0054e815661b0ec1cfb0f2fe2c314094bde79324629073e162a7d36b1c87a7fe3096e58272a8a230fad6fa51e4c1d693cb49da5fabfc10cd966f1b09bdd1f0312aa36e941199e892b7f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5629f374f015bbd1051b11441b03b84b9908b9f7db3e33ab3eb9918ab01eee052e91e648d86149d7d30d03ccaf0b46149380b51b1d957c6ad3b8fa42a462805f657bdb63c9d5fde24327d60cc58af782067837fc98f38efbeef2b53681630966707;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0997f6cb56bde7bfa3c11287de7ed9f516a216885a290834a0013a7f95d962eda88321570aa0eeddf6b59bdf9f5f0dd61e720e15bb894037335bb25225df71424311e5677c60419373ca6eba3c98f987dd38ccd2da5969261c29febdd49a10c687;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9bd158fab0d1d63ca3d5770b92dfc05b8727f1b68f7b93fb59f4775cb0995035724e0562493a721bc2c1512443b681cd025923e6591d5a2f85f0c3fd8dde9c2a7058a176486a4fc4204d3aecd187545d853cc476f3869cc09bf6c0274e35a38accf1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h721ae617aafc489ed79dcc7190650cdc7bbc470bca4e2511b4db5ba16f6fa42f85e0d80c5e8cd7cc9be3ec965753b329fc134d6ec85cd91cc7c0f98be8c9b85d7c04a6f73b73a214d3aed476036eec88a8862190c909374f19e64d5a2c2d44ba55e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd8ff162e716c8c2e338d87499c24e8a695825800c4beaeea790df164175ba3e9bd555dec14e3226f7cc75ea356c81261c564231293a84648705b56bdc1859e0b79918f5b28333b2ef386f2ee26378f6999cdebfe3c48d62fe67eec8c169b8bb948e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f06bb6a9eb7c8d2eac04410075cb8447c35ad430aa8a2bd194ada142c931e8e417758f5ab0cf5adc000b611ee8ac6a9cb44a31dd7613e5319bff2fb7e0bcbd0553408404c2defba94249e275210f68a55cf023576c6da0b7fad09b04abff999674d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d5cb8cf00e8022f1c4fe2a0ffa057434b6f7e02352317ff75bac1d3bdffd3ed0b2b53909769e1a24a4a732e7f0f566e9eb3ede27ce179f17d82c3166e9c3b2511c65082ecc8f0e5689830e7fb92d7a1765a5de294e3408c20a0673101df646da465;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc42b0271bf24f745dbddcf64a9d4cafee8811133b2917881a2b06775a2faadec5f7323ad1a2d3895e4ed3390bd07a52a5a77f8bf07aca665e28a7a381d8d59d3df0a2ca9afaa4dd7d83e39c7270f1ce9de8abb08686573360d52b8e7f874e6b1ae88;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ecdc093e32d79d535e5c37cfb01f878688e86f9ace570932431a2149b075542fc0b3181c02538cfe1702a503605b0c82cbda76d09aadd09774cc14b50664df936237b5a03ff12e5920106ecb9500bf46be2a9433e4c60fc0dd563d168b2f48a5ed3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1853cf5cb2b84a814901806e5ea138497a08719e5e5fafe4014d470ef7210564361d87bac6b368c7c7d1769515a84015c4b1e179253fd7f4a81dd1a09a581a4311140d9cb1fcfa9cf6d8767c8ca8a74b81dc32d9780728eb20717017c5d8e7969807;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b6874df7cb21a0aa29a3e58b805cc181a4c3f0dc464688db2c045e1c278367eca789ff8c17f69eba993bc9612c905c8d0f2917af419f9d38c36397b5282b1263fd32baa87ab5a4c9c13395282ca907982f948a0e3114feb5f867458923c1c0698f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8321c1ecb916688b9223771971684f03723cfbae3b48d679c707f7d28f1c88b8c4b71cbf9d5befbd15365ed2f9132db2c06708afa3653001e768954f97924a816214cb29c4b747672368940816fd1cc0ecc70237cd8b41412918016875cf643ca20c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ef1a8a068edbda05af886398f984a79dd188e1216a1fb4fc956590c64d84cbe026e56ffd9be76a430ed7c983a9f238b63844d2f04adcb8c89eb8f1f54f74043ea6106d66df118cef42a8472560b0ad0d5d71075f4550c024a55bfa7d9e32d082c93;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21648aa4a8f61e0d8b9ef0fb1785460c16a4e786818a2cbe5656bd507ed2e863df89a4288fc39c7680701c10d54568f5ecf17c7e81be3945790cf0e59686d52305af6f78ec1e1589023fa273f1d4900fe2c445e4ba63efad756ca509b9ad609c39f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60d6e6d7c879ec6e8d35d8851ad49f9c0c437bf97e114f88b1877d1ee0f46a864ca62864e0db046f47e049a81e92db06132516b6372637197bba2be65092bdb30b409d36210570c945f1d2ebc4bb91fe84a4d572bf180ae407716c4bed957d667b18;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hada7db25e75130a0242ecf544e17affd3fc1b5f62e2176a4a719a408c14d58e86b25eabda660fc53fa0ab6992a6790bb9aea655828e127588c651aa115bbc5c709e68bd06bbff25f7479a6a6eec8d9eb04a535785ce43975e115aa903366023a5523;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha194dbab38a39ba1a6c0873fe83b00523c858fb8c1c31f139e2d9ee8f621420dea29b9c3d1b45dfd419731991e31e5ba87cb53d7444a8eaf2f3989d20a7e7123cb7d3adc59d92665dcb1dc3d224e6193daaf9ba997eea92b115e2964d0eb92d4b067;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80cf26f8f98f5ea87475ba6ebfac96bb512abf6595ce1466d10314432948e058b3910830964a292b86bc1c34a112e13487ef4a9bb79e03c1482f2e7a31ed2fda762dc0801ff9fc6955ec49ef4a66fba38bde4b4bdac711192271ec1a2ddd8d10e538;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3033485ce4edce55e7f65c6693db1f448b03a5227c4c1e63af8ccaa10f2ac36f31685dd449e3daf5848a14a1fd352cfb8f16f535261dbf10d78ea40186037a299630b2c8e02dfdb1d626a27dbf506f400ea1b65ba3c7249749ca9549c784569cbf2d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ebd373b54af6e02b41f7cd545d334442b8503882be2daacc026d2ca77350c5f661f6ce90519bf6b84842f0df19c592bdccc584deec0f7c49a30846a78dfc67d02fdd4629330a1e85d661e863135c25c43c8ce09e349c9357ceeb8bdbb789e324896;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6cb2609d84f33408faf895f3bf1641e5b3770d8ee45faea4f07bfa654432565d44628b36ee6acac4dff8782f087a600fe8d8a5f17c5509a232a0b2594d7442dc962498c8c82c4931a9d9a2391221591fe1f3fc14486b98a8c979c9b4dad459beeef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5e581d01a41d543184daa2110a30c49897b07462f0a31071a9a40eea1e85d013f4dae41b2e91f9726caadb7c97d912ee24160f8ae6b18572c91bee1454a4f28b89df9c77741b67bf58329fa06495f54a162e4db05af8b74a2f7cbac7c0d9eefa6db;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc8a8f52d54da22aa921ec67eb46a5a48c93bb95d640c0d432aec6efb9cc122ce57b6e6566a49777c68ea386c2be42270928acad56bf07e5277a6c997824a94e2e558fdeb78853176052ef9bfe8e76e0ef27feff04eb9fe31d1fa58c07cb0b9249eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0127114f6281aadd8a772657bcab122aea4e951260b02fc36d99d634031e2d27f0cedd43c3f79590938bf57b59d48adbbaff40a1ba0efe12bf17a5b93b615f996f310536bc071b0c666c3e855a63e4a0feab34d7c70d950cc8d5b2001518961abbb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0e10620d36c5e0e6b6262eb60fdc96069dbdd504af5b877b5cd58433be7552ab60c6b79a23892eef1506423697d57cc63ede1635e05bb1e6d4b9da1e41036081e41d50e2f83d6c9a4f333517de5e31fdf65a7c99c0609fceb207b59403feb5ef5bc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28c148816fa354aa8985601cde6382f8d225b30102c425b239d66676caf515280c2093c6a7951c6eb61ddc978403c4384defce5327f5a91384569b71eecb62deb857184a164c8ea6d50deefd14115df4d70670cd16ea61d8b12d88128a8774a30041;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13fecbc6ee52e8b135618e21a413079efa262c3c4ca5cf64097b627e553cd02ed29dc3f9096a09f2922d45d82086355fd0c6fc690ea290a7982c842198675b914c3cd7e76b7ee81df57223001c7d3394017ca9e55d45e077e3449f0ce589c21982eb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb902f45d3ace98c3912aca65086c79b895a744f73caa6f8f6563867e2250b60beba3a8de1f0aac1062d986851efa0cd67730d532891b9ee43f3630849682f4db2eae81dc931dcc159a5a9fb39aa65b310c2f4c4eb1cd31a82bc22d9d4beb7e2e862c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72fb116dddc2e38e72e3abf7de51411bb8020a52d05436e0dc420d7aef7e1f3de54d6f319540a78373c807c536aba8ada1ed78f6de891a91c3e612684a212c93755494c5efaae26ce5270f4566172c67c5cf37645426b01837dc0d8d5ca487adfecc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18650cc7c0860397b10582b42ff05f82d94e53ac65f9a02614cabd949935bd0952ecbb24e5f2b19579376746b68d1ae8aa0a190cdfaedc02f4ffed8b94c83dac8d1823a11e5ace4990b4828d7698d9706cf0d97034f7ac73a24a609ad77aadcdd23b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd00041f2ff3cb84fe9ae0e255b446062871809a762274393a1576ac280757478eaab01de517a4828c410707f7e57d9d82e6afe291da6c5a8077869ba40cabf8d5f6d9d4bc9aa3fcb05accf1db5de4f9fa0821521256b3d706f8703b5987cec690747;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he668e940f73c258d39f0d7aa5d16c2986a715dd80606b798423a17dbd1a859e3a8ba86e1abf05ff4c3952d5ad6363a45590582e5379ce5dba4e3a3f0c269274c7affaa3cd34f7fd013ba2ab1206a79cdd9b387bee3024f65d3530db9cab95edba238;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bf92e5fa9b6e700ee0e04a3cb960b7e7b279fd47e6f419d2cddfac848e6af64a096fce3f880746df92e8d06f0049b742bd1747c1e7201b45306c0eb04789317610309bc449797c2c76e6600bcf487ee28fbb4b18f5e1d1eb7726a3eae6afa1d7564;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16956c8ec63f714a1cbd967c765342a7c7be28d286e0d323b84624013f3feb0f5d76cacd87603ece8b3fab4c5fbeb04bfdad383f619503d92962468b36f9731403e7807d4877554c94d9f54045985ddc9dfd8eb8548d25218d3defe3fe421c67688c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71a67a3f83265b87f0248bb96584cb1d61ee4a5da85437d5dc7531c4d5d5e17cc8074969a1b80dfeb115dc3575a67a0a50dd6a6ea14fe2bf3e4c317ce569c39b71520b11486d89b0e6701a0db8070df086dce5d802643da01bb9df1cf0afde055d2a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h740f995b184d889da51ecdab5f3b060016ffe703b90bff286da6d22434e01e9f608c7da259419f360640921945e81878b52fea37f097b41300f9f22199c0e2102f35fb071c76444e553751cae9c42d2c22f651a2a9aed486c700c26508a55f5a2888;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb657ed4ea83fb28f6127330ed79484f315eac3425b6fe510bfde1462ee786d0c9ed564519afa4a6567987baec191f4557b836baff5aed282a70a1fd8ca8e7e4cfa7dce99949ca081a446c26a45cecc0505dcaae75f51357f5dd16c837d4c690c7a13;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8437f5789f9e6b6a0ab286c8c003dff01c0be4d9f04739cc68e8e3ddd969f52f72b97eb979f2f866d52e802ae010746fd2829a62fbb35c2b1aaf83acbc00542f35afc95742998769a61990576858d5565432b2ea772231f76e584ec1ce9be85ca0f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h160a886e72f778a3e4ca2c1e5b728e22ad5e667e3178c79e6eecfd0c3897163222f11130905f72d19da56df9ec616dd1ea9ddfcd4f48ed26e30f55b92e78af6ca3cbcb80c01c9af343647ed619459d9b71ce8221fc69c494dda84cd98c6f64e24d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8e28396de0e370b646ef3736980be7b4d58335c6ea5fd815d67597a0d8ee94a3266ef032f1a690760c008b85ada8804de68b1db35e2a04af96fe54313a86c4ada060253dab2c14c2e4660f049fcc7108c41ad88dafb5dd3ae64a49b12bbd2f988c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc3bcc8eab5e42dab0933087729e6e5dcac426b5e47368149bf94fcf06e4cf5d3b36f359a38d2ea80e520896e80da6706685fec41247bd9185edd50e75d237898bf8a492df9b52b496336f600804f860606831bff486d6384991d02cacf9b3d4b9aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dbe6b9b0263951e190387096123b7973661ebcb21fa1e18b114626c4909ec8e9963c768cf8e2f6ec0c92f6045909d5e44f51b45da64d7b97575f57522ff53c49050fb50b4af671176007fa72444a0e799868fb0a14e46a91ca9fffaf45f27acdd33;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96f68db478c03502fc6a147cc6811a706181df502fd9cbb773318f4d1b1921a5ae7cbbe6b2cb2da61d2950d016a80613b6159483759070bcb2adc1b4371e2b79e07e204f0eef3b43b0a9be738e280dbbdaf6b168aad16a148436ea026b4d9588701e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe179af324287e459a4ada0206b222e5b83ebfa6be812269289ffbbe22d804fce13617ec078bc46382e7a3f97b9af101cd71f8389fb2dface7512d3677ada01e239212e515ff1341b08b2b783d64b261e7f29c1e6c51a6f495d020f9212deafe633c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22e3588175ab2f4992bc881fd12d15f0bbe37d5f6c0ca1caab5f0b0224ca979520d28b8ba550fc0a6a69183c0617a93d843ce0fb6d1e1d2553410afc2e4afc954fbffba310ed639ea7c287f3b8b3efee648b80defae4c4551df34a2dafc324fd8bc0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8f158ec9f0e070e9a9ff8a687378e79b6cb43c4717c1e0c8e1ebbf0d391fd66d5939e392da4cfae4ce653945a742370b41dc39ab211b729166d8306415fb4ddef8deeec829c687ef7a6887aea6feb7b94f57c914b55cc12ac37ef44e2b9d8bdc1e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41d69b2d39e6f88ac346c8fa75a1fb8d9bf637bc9b67197187392387cf7f2148954e1cd2553ad07ee0c07a736a940d375072d237373060d560082905566bc138a4c00d5934ff29a38f9d65111c203a599f3108714dbfcb85ea7b7e8ec2e297328a04;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39b0ba3cfc2d745b61e4757947679e2f69f48242c7cc570679e01074fd0f7790cd0e8400b004e963fa3ffa75cee0b0d1854759bc60bd4f5a455178ec1fe484258c20e3736a7d74d5bfafe5f548330f6b166da89e6f2409c45bd7d516d9af1118b76d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ad05930eeb1180f3b88d1c4a6bc9750ddaae7734cf82211e8dd5ef3a05249314ce6b01d8ee01fb696e0dac5d2053328480081bc9b19ff2199872a29100a5fb7d6a4ef00d29b74f0d3c97912641fc84f1394fa0e502f34c0624285645e477906dda8;
        #1
        $finish();
    end
endmodule
