module testbench();
    reg [21:0] src0;
    reg [21:0] src1;
    reg [21:0] src2;
    reg [21:0] src3;
    reg [21:0] src4;
    reg [21:0] src5;
    reg [21:0] src6;
    reg [21:0] src7;
    reg [21:0] src8;
    reg [21:0] src9;
    reg [21:0] src10;
    reg [21:0] src11;
    reg [21:0] src12;
    reg [21:0] src13;
    reg [21:0] src14;
    reg [21:0] src15;
    reg [21:0] src16;
    reg [21:0] src17;
    reg [21:0] src18;
    reg [21:0] src19;
    reg [21:0] src20;
    reg [21:0] src21;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [26:0] srcsum;
    wire [26:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2be0b191160b23c24518a7f67f97a97195399de244fb2468b0f5a83e22a5de046c192ab13a82e25254bd6c609bf61d6175285c39439e46e8ab8437d2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff2d7df0abca67a847ea2fd8033c00d5f3f9ce0e61d97399261bf23e19fbef14acfc5bbe71d1db5193bc7596d9afcc383286d975ff3be3f92cfaee7a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e9ff46e12f32996a12b2ef6aef677a4e1c8dc822dd39a13d7e51478ddb0ebd08183523cee553ac7198697994cb4b95eb65088d7340b6cf414e13b7ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e07a61fe4750d7527c0e539d8a60cd25333714cfdcf26ec746fc76d4afec57e61ba28f7f06911fcf47d60435b6c150831f952c3af240a42557eec942;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75e3bd5895f17dc4bbaee57fd174e343ce70d595ee340878976bfed2c709d9b1b9cf3ecd2ed5b4064e380cabfd4884af9e09edd5dac717f9adc818c56;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had7d2784bfc9e8cc09d95edee007f8bca695d1f68705807f76f2decd43b6abb5d177c4aed3f6736797152cb4752028b817702ae673383dfac80a8389f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf5590433ade48cbc6a369da4dc455f66c177462989a07e12a49af6c4078b4c272bc3d4bdd5a169405c8daada76e478935af0fdda3f9c510327a6cdcb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d84818aa5e380b25dd86cb974f5b45aef2a459c1fe7ee6a20632bc43d4be2b1021e5fe0e14e29614f61d1495dc91a49843102df385e9ba0353acadcb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h707e29ca2829dec9984635e12d2b103e07a9c487682ec6b9dada59ffd1288147e258aff0cf9c1d5f01fdfbc5c69c42728a8601b55c1a4759ab0c229b2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5e39ae877c4d6c94b99a365fd9aba5c820154235310f15c6b0f7700991770496a6533b14fbdc00a9a9be652b539a5caad2d629e4fb84977502521d85;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ce150473f544fdb088e3f94f40ba7bde5d0929050b7d909fb79c1a2262664a46e97452104a54820fd16b51f6d038ecadd9a41a61628973ad49c6c946;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c20ff3995917f41e7494a242195175a6738e82a32957b6fbdbe06a03f0155c5769886ea7057c44c7feebddd1da90a2643fdcc15e88613f6516f49fb8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h292548626c5f8018e90136e70f143d0ea3f3572c15ec466b07d1f311c3c5e2acbec0bb259742cf40b38c4a5d453c01f223d160c405a334c0f36c9f8fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h280f9a74be0af53e2e7fbc91ab5c83ebd7b61babf7cb51f9398127edbf65dcbcbd6199105943a26753f71d96a4fcf32f6138cd8e14ca2f89bed50ab69;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9b6e9be4674510d422f17ed7fd79d34c7f2c9b2c39192cff567f825070432b8d3e61a670860e0c8a02dfa3e2a3587748add91d0911b61417d9ac5ab2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37a53a9f237a1bc75c82b8543f5d2a06c5e16a95dc09749714746beb9eaba690673aebe9f88af4fd6e227736ca65490275db220c30864cb4f4125af85;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heaf3c4e8468db74cbe4d206badfefc9116cdc5066f907bfd22f53542e73e91c500bdb7420b1b537df14e652bd89e97518a6c328868723af0901110560;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96eb850636eeef15a4562a47c7080409cc884f43f2a7d29dccc4d12d83ac08503e315d9acaefe359c8eb26bcd2b9881d58d7c18f39a73373ea28ffbac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe1b03521505e490a4df10691ed24a05ed4911e6dbaeb242f29e63cb94652cfd645b3fa6aa494e2d2677f6beeac585aa0d33100d4b3393fdcd3139f29;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h788990f79dd1317d730790c83079efc0e13dd0c697a0dd7cd51d4b714b917605d23d03ffd6e72c8f360c693cd764d6a9da4ebd9408cc92207e750dbdd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ad38c8c864ac75e78b61869dc3b93df06e358d0a08cc47bb327d44e52fa1ff3ed0ddb17077841fdb60b020ed0f14dd4f0e4abbfc24580098efb04239;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h300b9406c6591481769599cda276ce9f93b39fb5d65ec000d300077dd1161ccceaf0ea0d68cafdbe54677f87ebb924ad64d98ef1b8e1d5b5f8298cd12;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34498d5499a17947894fa9557976607e47c2918365b885549948b631082c4071097b23223ff4c799c6b235c064bb00b9bc82090c73e82976aeb624b14;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c5b98546346528d7d5d38dbf49779ce7c11da54daf04fb5cec814a962b9dec9cecd2d0270ed6e9a046d97e875a1e3abe0d925ee413422ce2990e1c90;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71d4411af37a71fa54534192a6c383cc7ea9eb8618c60e719d61e960fddd584ab6a2d255ddf3781b405a13bb4d43417ab7f205976a7fcca88384157e9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64629ae7f881ce75b7d02c60981ea554116f4b98a0af9830cc4932e44a83a825103d0539dc0a6c2ca7676db50fec4911c6ce48fc5e06f008daab3a4f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2543f1fe843a618d8c82299c592113db95a1b946a85efa5c86ad576422855148339833992acca66e5942a1c061269305aec3bbe8197decbe59214d051;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h252e30313c0431bb4bdb8eaa4589c07004a2c8fabcf11abde2d42907d015dbdb2c03a097e976296a0f656f405c79090ecef8e1c6e326086e6c8228ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ba20acc703301cbaa9ca2a2f1d1aa6df49d8af7d9d254010fe259c440e7e8f94282cebf7ceeac00517e9e752d95379ee556149029be845a5925e1022;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd975fffac6aca4a2c651c10956a3947202ba50706e4f43841ab48f08275f1c622d0c4f4aa3d6dd804388f3037bc0d0b42802ac105e3ccb461e414737e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63f67269506d88e5a394069833b8a25a35c343f3889ac1f6b7b2600461472e03fb12a52d312db1614c039490d510b693c668c15aa853cd486f1e515c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdadfbbb51e78f638535c0f1b4115c76cd4ff50f96216e4f645b11ef8e863421eb3e448bce3d7fc43f7cc2c4e3359dd04a8c76530254fa04ced56b824;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec335fc3e4bca61ee162ae59cfcb9cd6dd85722e70a0db223497e6556fbb01eb3310d2bbd0e2727b4bbdf700169dc844e8cd521fc82e96907d9e3592f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd64d2a0283980b95dda3c52a5e5a57ea382704157dfe4592bb66781158f1d157d41ae897647dbc4f2343dab29685b5de00ad1b8168481a9e1f3e6ffac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc79df212a38ef7bc791991759374ffd50a5bbae6e078c9491125ae49973eba7dd002bf65998f40ae11fee5da7bccf25ec76838f1c9111c9a62251fce3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9867a79a4aabcb0db68a39084b18329b1f5dd893cea7d2511ac2e8e512376b1e1d24eb13bf193421b3a60b0e927c0f97e5bb46132566897fe9ee0a103;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h232325d8c2e3c58db8b1e9f1a252d4134a3b1b6146f6aa4d8dc4b93ce95d38e66d3a6204fa47ce991f0bb13af7d7f489f4860977b783ec1d93d926ebc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc2119cac183c006949666873553d5ca7aa09b06f79e05165aae08ff4a6910cc9412382a5a702a82c7d13a535d580899cd64966d24040f061ba32e83f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9440a6cd0de33d6f8e762285a19a358d28d2a87980f29ed39a8aa4ecaf30fc62908182509d5528bd8cd367c80a2d408791f668d8c4db81113b01b343;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46e9cfa02fe0223bb23e22b5558d40431d4408a5418c391a115eedc5419a09c92fd9b014969e552905a2bf6cdb53793a97ca21a0a9fd1a77d9d6d7599;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88ef54c318e0fe7f87523ac9c392e3c260c3647b872d43177926e0026606bbb69d5a69fdafcb3a3e7dc81ba1fb3dc6e2a83d5dc9b2c7d83cc2f116479;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3b1693c4c83c202f5321763cf4f734563a8e5eeeb9b6afcc7f055b7de48f03fedf8a99914d723d1761cd5c1e936532f03ec62d43d77822e81a1103a1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2b8d62c2e26bba3e2b81f0bb91e9d8b191d7e132f3a8d171ff398aa46fe7942fddd906c56429d86c5e598f2050853ac3aaf797c3305193fec4dadd1c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he17fc99bbbd2f17adbbe192b0d53b6e723451e6935e12f7fd582ff708e430604e8a5f2d73072ccdf7cb265deaff390818e946ca834fabc3a10a09c7ec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44788f70ea5fb728c5a1faee309c245ceeed786e133f5d2d8563297c666d38e881475487f1f7731ddc7b8e3a5e07780ac494d593a53bc0962a4740367;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb655731e4a96806a95f7c6d0e4347f2eb781ef5f7cd985b8815e16385d042df759ef8eb6ba5c63ff33534af8dbdeed55633e8049a3748e15d19a77cea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc43592be6b481c3e31638d188191c37649b9db7b41d05f4904429e0356f52ccf52ddc63bd7a3c5f3dc30e8b928317f05df8031dae3374faa3a1032f92;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83b6b0f3e3dbc623f62886c54fdcd2af9c25294fa7d75ab773e722a7b3c91ef714802b6505fb2d6cee88a3fa86b9046b779d4a44463a80321e48bbb78;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf936a7f67160a023c858d976cbf2e779389b64eedf41835e7aa52a886949963b2838f5725d626468f32f37a3b872c8381b2870fa2b29a34544e58bb6f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd90289fc48eadd5988d19a0ee8c832df698963358c524b6ea096257050e39d8fa44869efea11701c21334b5542b698e3198e0477717274472a2008035;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3dcd635b04cc8c02b14aef354cd7da07ef302ca81238a7118841a11cc2fa5cac4de6334896454d8d3ec3ec4f8af0373ee0b9398157d36e822d0b4873c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33bda5fe7b28a8e90178073e3b05caa37e5368d083d07082be1aa6567c80b6194fb5b9239a8f705a82f3b264c9880b63b3efd73feee51d0b2617ae973;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdce247be739977096db66e57d276533f4f088c96927c0167d49e3d18d59301d36b47c98a63e17ba1548cda623568562c37165c1639cce38750701b01a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f628136f01c2151fee1ad3aaa835fbe80169a380f0a28cb01f8f5b7e91952029d4d9dacf2bd1895bde6887dffb559b569e080663cc400673c2daa7bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h648cd5fe3002918f043bd08385b42a1f495daa6c6727cbaf11d7e23faccab61c7ca2d39b601c993ac738be0393288ff8c620330db2b8c6fff36a512ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b39dd55c09dc94ed941332347e21be01185dd7c804e98646fd627abe3a5fa949aacf3eb227fb6c47256936cebaef49b68c4b00ee5a61031229dd05de;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b834ffa9041016566c70f99efa236618416791e5b04287b9d9d1353f92e17d23b8f5432620f828f2175a3c73445f861255ecacbb2767dcdc1f1bf1e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5c84cb771017365dbfd9095e53ea28778760f3262c35e6f6183b58a7c3330bd68a92139ec9fd1470a54c41dd7cbd031bbd760745d3ecfea82b531b71;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae79693aac77844d07972f52a9f1c9f40f4b47d958d58e1fc1125a1ef9ecc733b6641d94eb5ef27b64b5974ef1d2775231b8a6e2e10beb1e4ad3c586c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf898118ce97110866dfe5b22526460d2f2d1ca0874fb11618bbd1d51d5f8d52053f0f10d308677cee6f58e216268880128c375b0c5215be2fdc0b6bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d052331f482263a5dd76e1a67636a370f58e625c8c77a96fd5a85705adaebf7f78f31b0425f542ebfdf8741b478c6f1a88bf9957420470bcac9360c8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24711fcfab0e1fae4c06ccc92e6d8e52a09c815f730fde5cb4e8ee96b9ecdde69051f48f7862491acd738405e20250d29b9dac51e36243105a5f8807d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8833509613de65962971d9be482cf401e8cd02d45e4a5bfda7f1488560b777d1c434ecd087d0f13ce49c06bba3e7e2d6417ff4502717d64d28edae9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h741f0b1fc1edb658bd513ea5e90afe973012d877bd501badfaf63eec058ccf6d1f3134e59566cfb42d34f2b0d5d1e1f303e322f47506c736745039e60;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d76a20d7fe5e90eb935c8e6e0ef359c4add75bd287ac80dfcba31ab4526a7728df28fda8b9dffc4eaf930c4d67f474a848d13d2ba902fe0268b21fe4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb568cc8eb5456fe2a1eae5eb2d8d2354135528924c69f88f45cdae1cababe1c250e1a5b3cfb85334b88e1be4e0f8383c5a3f18170881540c11176b9b8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd60ea691319885334a11173e7339b2c09358f89d02a4b802adf06ae014cd7e8712249a8a1be666a306c326db1da337352ade19cbaf42ad889d68b79b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h347888f645b31769c427ef5364596686d446645aa7c2c1fccae285cbdd64d3bc10d8d60c3ac0084ff4fa9b757c38078a83edd56a5976bedbfef05a6f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc39900985fb2021e046db949012e3e888cb04faf72d9a7003f0c3df1e7215782cac03facca85979f7417f5ce2f41e060ea8f833cd887d0906e0c2b1a1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c1fb483a5f84aaa1c62198f5c5d581692e8b5e80d5475c1a3c1590c9e93f16492f1b82419a948fc562ba493cb622f4d40ea828b7795b304b9c6b6eb3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b69830fa112359ffd46b6c2542907ef235c07a759e286e4b45e8a5cb0d9ab2d0611a1c2776ca2bd8855915e4f74b1392ab3b88ed8897dffc5f449539;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e12a292c50d5040c05cb1b503f8b0830e8fcb4e89359f8f42066135952c1a3d9d30a0a94d66805af39c8a23391ad4e69046b691405420a525828f4a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h903c5c1eb21076ac932d49e36ef8b050df9aded63cb7e5b9bf85692c0179e7ea4d6121a64640c738715e74f12241f598f4eab75936d4d3c301308d04;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cf1bf3b193374babc6036ff17adf608802234554ab2aa1ab96be0c4ef7b1ccb8a2bc3381924dcfa4b173625632a5abbfec8b13c1b92e8d1358ae2be3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7dcfb7d2eac6015953bcfc2a3522f68b99ae20c00fb1c3510119849964cd0a712a9fcf3c40d4ebc94543ae0777e6eceb57aafe72412330b6652b79b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha76ed60d68fed6ac63b2ac90179f5cc0c64ae7659c7ea3947ea7fe4da8ac9952bc983aaa9640da0f141ff18bd680e3634cb912abf74c4b9b78b0b3904;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc21afec0f7ec54cfe69406dea9550d2e080271ba5ebb112bcfca8a627376c025bdab0f5ad6a6d0060bf268e9734229e018ea83a8b73ad11bb4a2ccb9c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1dbbcccda73ed6fbde0ab92b142516dc4eafdad6695229dcd8df3e7be643a941b1fe3df042483c01f97cdb4b4e56ee3a2d23b466747e06f0782793e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ca5d03bc26bbaef351f96453575e964937a541dc669413b9c9d28363054b90db7339fce4380815628dec1436c581fe5373b90f6a5dc98f94e8573a1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24bedd43ce300c7619eeecd6d6dbdd25092905bda1a434b36247bcca2f2b96bfa7920332c84a10eb977416c83b821d68ad5f3dbe9d986cfda42cf5eaf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51ba772a543e86c8d3745f11d4c8011a6c8dfeda5a719d9e395879343faf628841cfa6320b1df243fee4eebbe95f216360137473156ee030a7f20ca33;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12e2e7764e697b8ba6252a998eaf7716b2a6b695f5f893eb23eb18380b83057f6c38eec888ece41164476c98ef1d5819c43314450c24e64aa5155f68;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h202eb2319b46c2d6354cc20d1a7293e2f6b7cfa78deab907e354e2c8fa51751a7a58a2f3a5e1048f24622127bb45215b5ce1dc5ca95a19209a4dd43bd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd831a9793a88592a4dce770d20538dc1e81b7eb8eff6faa420858417e5f990de856fafa84dbe2c8ae489531dba7b724f37dc74c9ec30c5d759c712ca;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29027447627b16142cb0a0969881ad15e4a8f7be93e266ea479716d40640a689f5396b5b3406ff9bb2e6e44a476ad3e19c1b3990aed9e6e12208a3e91;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfe7c82ffc2489b98e37a99205bd8e019f8246189c7da120997c2c7da987c949ed5e4dd5df707046656452bafcb2847dfbe3079fddde9e46e869e62662;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h225958145705fb0f50a8494b3d29cacd77dd20d58dda98bd47be54ec85333af6f95bc290abd263ef21ab6331813000f5a8787f75000fbb8de2430e69c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15a4a7b9f7d64e7b6e92e6dc2bb5d24d60caf82f74f66f8504ecc9c8f95d994a3cae394c36bd84844e381ccd53e0ead9390280239ae69040a19341f9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d165c98726e4348a2afb581c9131371a4d71310c7dac19a8438b5819d56f7b275a74185b1999c562caa65a9a97e6860cf2b085a0df62b961f57b1260;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda85f14ad35e61972bf0001748de660fe04a82bfed219b073a0cac6d5f641df9468069238ded78bba92f85bb71c9758d85e6db99bfb13e5807b70a3ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62b56233c3cd329c2557426e03782b206393061ee63325763996eff6bc0a22ea58261bd69f9ea0da9665ee12ab2e4e0c49ea614548d4e1c34efb448c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha687afd3b84a74e2b02ae7efc6d5e611f56ad4efb6519220bbe14be17bb8ea0c5f230a834266e8bca0c88ca73d1ea1175bdf64d1cadf1139632ff55d5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9eef2022661f9ce694dd4fe689fe97179697b1761857241bb8780659d739547f9c40fadb9760bb96a416acb5ad31d587c5c1fd879394388b564701d7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87fab0a6338130354b7bd4644a36c5f907476e58293951dd2c4b3cf909d11589249760f0c551cee60363df5a27e4289586aa56b7aad0c63523dea958;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h975c13bfeb297dff3928c88fb0073c94e5a9f97d39b65c182f0335a17f6bde1ede2bac3a7b96c8f413cf5fcf2bad98d4ac146557a9f227165457bdf6a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha15d099b30c0adb95959edca5b1ca79a38e6ac8fabb0ac4ef7a2f50a7bf1cc8cfcb2f9372b88ae066be9c88100e079a7bcdd25e7400ef892fbfe0774b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91b118f0a3c41903355da9c401c74b5125d01765d9c30bb4524f48397ea74c08283727ecd8687c25338775415c64ef377c67d3a630fef4e1eecce61dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62426560cc6fd6bd622a47da5dabcf7bdd4625e276cdaef3d09c02102a2a438469ca72ad9d15f8c7b1246ee5e5636a3f7ee548555dd863779bb48ef02;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56312f2e50e4102b9b8c566370d153a21f766b4abd1c57f3c85b6a478eeefbc5f629964c583b486d85f713ce73f8edda84805d06d906c9c3f9e574d9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfbbf7a2b391b002459aa49a2aa6d5fb04d70a1690d537b2108e37a92f4aac89c94c4084428db83420fd77b0c8fe44b30809abba85d34d464b4126da95;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4d3b088185b65356cf081162ce15aad3939eb5f06b3936a283ec46c88c5b82bdf47d522369533f36b0cd9feef0f52724d95400f809fb09dc861cb25;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3158df67bcdef6f5c2de4a3b51c3f2374504e0af4ab0d8c9e661141d17c7dff9e769e7a84f6873daf90021748f1472e77bda8a583a57c7b7465caff1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h594d3bc45f8438780eab90063a931af5e78308b6db20496f0c388c47e5e78c8a2acd83fd8b06419a3c56b4fbabf2b9173eb2eb006e69590e30a8cfec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9aaae20d1c5f15e01f0b027f8012c8565a3c62a5392ca3a8a37421a852e7c7032de434efeffc5ddfec41832a5f858468eee78ee2804371e4d5958155b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3cc651b17e1d6de1aab0e51f4de67f82fd53aaca4958caf9a3d46306e8b054bbb8fad81ca899ab9471f9587b89beb4255dd6fd01a4daac2a9b70c099;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c02cb5adfe99f0bbc81e81b7c9441d8fc55b338a06bd8a987e40e49da07deec8bc923bf9d99d98c65eeefbdc898f229681878261388e5d7ec6216385;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfcee52f3d9dd670b18b0244a75cbad6134b42297cdd4e67d1de4da8309fa6976a65cf4a3d869715748090125d9fa87d4bca43847ce95fadba4c76b29a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ecc3c86989be195c67dab9ad644d466030f91c32575cf81e9d3d632bbd31d1dadc7833e41b1b6f1daa58343e45ca07436390c518d6ef97c27bb03333;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1062c5a5d64afc77a3a1929ba33cf09ce646b8adcea0a140117650553d4fd0373d0435781291a0f1ad50415d77aa0699b2d679699561351053a876394;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h957dfe904d582488245bcc03372301212cbfda17f993ff05026f3d1b9905fbf61e7977141508462350ee7d94d9e18955e0efcb89cccaea4a4f63d5777;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff4a466557ecd189ec9264a0651076072600d66352973b07ef407adc2cc98850d1e224d3264dc61cbb72bff44d179113399ffb5238e7dd771d79cf75a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c1c1efe94930e22edc7afdcd33cd5791c37f82c1253b023a4afd446c2a940f263103ad00f6f0dc98fd1c1c9a332e1391575c5b0d251db876d7241e3a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb821896ecbc061ade9797eacd8f9400afd5a321fc054e4ba8a713144346dc1a6c8fd740fd8bb421a7645d2ff5bcbc18f6a7ab5226a4d297b9b72b902;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f6b102d1ee5bac00d249dcf0c66a2a4c9caae78eead3783819006b4f3d480d2a5c159d05cabbd2e2cc9948766c5d3bb6955ba3fe7eb93e5cb4ab50ee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15e40df20ea1ad749f4df2e61abd8142fbde59f503a7126c1596fc162c6810bb6ce8a131ac3a767bb72aafc65015fdd33081b2ba1dc3c7020c7da99e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd294dedf8cd8cc12aef3e352e683c4a718100a679dbde923d4fea1b6b0bc226f54efa4ae840289205ca2ee3764092ebab5e1a8dfcfb91791b77efe333;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf9b531010768a311ffea7e186fcac8f312f64a021a9a9fe674c5f387371a51ea9c791ac76e6fdba348aa71176d0c4bf24433aeb0808e66f2d7f6402f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e551ca8544f361cfb76953812f91e6e972741af24406704b7d0e7823d883f74b363e4dbbe26b15b249cb8e0a17e636e931fc6d04495f3f0110775bc6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43c6b36f596641232aa175cb94269e66d932345a9400987f9e6c0fd18919030ae756ef5f04c2fffa9831465bd909fbe6a58c5ece458ed80b5e53b4579;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haac74a5c1a0035e47c14b62bcd73557c7ac7c4bacdc0f6238c86223a306d17e55763f4bc6518610716e4440985a0faee8283e85f57fda7b924828c83b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24319f3af28380771d4d1a0e0de0cc2052200dcae58dbade822b46270808d43afff472da5b78cdcdf9a39839cfc4d57f09f611e62bcc8be3c627e3a68;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d9e3104bad5cc419950bc6e2d6ccc6e3768208d87656a4eccd8ed3e8e6ede8e529c8afda3552c57f13651efbba5529720c441c500ea869c1ca89a29c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h802847e67a3916653aa53a971505bc1b952db0c2cfb9f2066fc51b4eb33c5686a289b742e89d3d61138235851f1a7231d6e350eb5bdfb08a0c131139d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfbb9a2bcfa30889c5f74801d770d840be18a6e2e5dc46064eb9c8fb2fa7a83efad176ad61476c6e18d40e11395cb398457a4fa1c55a38390d1dd10dae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4f3143e30af42b5a7b3b635569f8577a1310180254dd0fe06737b66886dbafba559627679af284369e033f9d8ed304ebea594eb244da28b38016fc5e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf776c6c1a9c4cd8b873bbf2eb1a3a93dc33df6e4fdabea6018683c455a28217fe895711652ae2a821993a1afb3eb5710d99ed42f053fa958d64713f9d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bdd8c109395d72e048327d172415d2043ce8ccd5de04df0b614779dddd3b02c25b32c7d2f453c35f8264dc8d21f1498787eee1daed388d2e64c7316f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65d35fe6325a5088bfa05e97c180ff7887b475db17742f50bd4ab878e703c231afff162e726eb9c18305bc655c678769b12fa68d1d5b41a8c694395d1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h123513bf6d21dd62feb36a66fd7cee18d32e1934157589bdff957ae1e5ed1c99914ba70ea89552e27550a3645f6d445e0a94f7666fc2d5c5dd8061717;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94e8b2d6cc3773ec9059e1d2d2f11f673a1457a74231e627d4c9515f9b3f24d569c80052969b9da7e5a7fc17a3614f729e3e409593ac4e93e3904488d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h329de089363867a47794bf4b7a52975e914af5d64c7a737a0d36d9a663222dfd7bc475ebece46a537e55acd99ecb326240d15f8fd149122de3bf26fe2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86e9f5b79e20840d142fc5fa3eb05e9a512248990823c5125dcf4f0bb4af02317c151204cf77bd3072f1eb71076e244b0db2ce19b381f2bac7253873d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb898b51f28ceea33ad19de2b81e68dfc109ed1fea4db9899e4e07aa9ef77719630a7dec04688df3fa62a5a7d04312337695e71994b5c341e3fce07e58;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h801ee6508073a67d6117b0602121768ee14e37324cdf485b17908359867af3d5e7652faf3c811fbf8b0e64e6e400425d12792498fbba916cc49332e10;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88c96a9f9133e7263255ed815e8a4d7afc82dbf8fdf95a7738d8c578653614da5c465f1ae0c0b36db5d3a8d1cb42abf4da5686775e9d94a51e747e706;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81cd88312d555bab9549484d40ee265340877666b96af5e1f2deceadb2dff9653a1fc0a39d9ef3479a24329b423ab05d2993a1390df9493864046e11a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha41c470269aebed7533d6f7d1aa06571ba75984268b116ada8d7dc04d806a7530631aa06b10021ab10490a287f35a893dd6591931d608878e852cfc65;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha08ba5179489807ec1fb5d50a17870b53842f9c75ea1aecef07b1bb40bd0ef1a8fffdacb4b0ba0a4a48e5c6754c578c34c78e9891876b9fdf75f2b4a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8077007ce0880e7681a728383af3bb6a43f8d141bbfaf9e4fc4599c38650ed840c4a732adf61116997f39b06979be6e7ce54712d2c6cd36de1a2e3f0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hddd619a411416c05b6ee6ef9e2c50accb65e0c10bfa85bf5a7ff6fd7cad495841782b4ec08f733171c89eeaf4817e20e6e3d66a1489fa14ea23b799e7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2692b8c4bc40eedeffa2ce69813500469f4c1d15ff408d87c068a20f7bb4c6743f583965f9b2267c7fce36cd4eaa2f5cef33952db0aaaa3ab733b155;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h453bb97dc377689d3a610ef7b1eab74bfb0bdd9319ee7814feeb178860252df9ff4e310172a4f64154787741536bbdd0e9d2d279442ebbe3f7fba8802;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b0a0e4cf6b973046e7c2f6ccf2c8d8a0e4abd1d273b0358bac570dd8207803188670546bbc682f188696578a89f864242c478e396e2f458582d9b8d5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h634aeed056244205aece43bf26b9944ac112f576d218549b069ca65564eb1e7ef37530563c383444dfc67aee425366e4f6e71eaf397c78a3906a4ab4b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb8e8901cd37c26f6facc508a91ef8bf0b2af8160b7dfc3e6a200c384e88fe90514ced8be6bad0c98f0dc17a75cd44f8a0efac6771e7f2912064b838b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc36c4467b430ea35e803289b7428ee7f4986d8eae2ef9e571a74855ff9a8a6ad1b556d1b035cece4c072b7cbdcaf8d144392e818114d2a3ff65eb34da;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7df765f0d08224b841ab0943c35d57b327c76bc606da7b1b38e22e102a87bf7367eb9866d3006d129794f6ef5c43936a2be13912c8419ac57282c38dd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he951f33b1d306f2efcd53f2f002ac71df52a5f4bfd706998c748caa64de90ce684f2c55872c0643b674ef24b885d8cf0316581c58bb788a74869a606;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8958ab60d6b20ceefb6ff750e71d6b105d3e23a882e4f93baa17a6493f7c492ebfeefb9793ba49822525fd768e9f7d1047bb82ae22ddc24b623f245e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee3e473987d14061e82350a33925c0628249b4efb12dcaf29805877568eda4df178cb15f7b4c8cb409fe3ea3e335c5b6869a01f6e63bf700391028e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had9080de0b7dcc15728212f7209164259f9fd978ff106da0a7b61acd724c587fb982c734e3c2c1488b2cbe8057c12226da5bbb6497904cb60bc354f28;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h400681d032cc298898627fd35187e6845ad9639a5b78dcbc0bdb749fe9727ed2e84c3b56daaf02047c2fd3c0f0162e8cff010f5f53f3fb6796b7d5e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h488b4d64c454f8377d0f48c89c0b9d6276a49f27c36fb2734a9d3fdc35b6d5a8d5624e9d905e02b71a63e60a6f245e64f0dfd04c2c99bf0b86602c845;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b997967a671a0d189c67e95f1a49e97a6763bdd41ed80bebeda1e5e1e7f0bbb8885a644421f2d67d8064fbffa7a273266f825d581ca0b6222bd92bb9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a5d4a94be16b87366d1057b4cce504a4f70510f6cd7132e2207610cb22b0213b5a57801e216bae8dea1896aa978cc6027576372d0450ac71f9a29660;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e88c2d31efb14b72620f658c6295251168fc752d976119bfbe986ceae9234ebea28692bdf30730da315230d4dc9f045ff176736f1ed97b64c0b9241d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdafccd822cd7aee026d39df068596e76490decfd20072f90fde39f965c1511b76b0085c838e27f2438af08776e507ffb8d60a7c8e2e0e3d7d2995977e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h341319d7edfea6fd4163c53a25a80e0612e687f95579aba8a206d3fb2eadc5ae600e84e3d804c48fee9eb40df82d1a549caf3259601264dd20b513fb2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cee372cf14717f30fdb683362668826798c25dd0b55aa2183cd3476e7a99885815c2d225af945eb6abf40e7b4fb3338a6cd808ada78449aa9c7b3dc5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b945668ec64267113a58851f93020211af0d8f0d618997d6af4bbdce392f5c5b10f9453a2e9c1bba7940102212eaf7b21a64fe45ee633d6f5ee43820;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6249a87256e520d116121288a3e1d89273a2a1090d9c86c7d88f1da8fee24719b5330381c6b30dc6576a9d26e2a905e603d8d06bdb38d2daab585e0a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8042df49da53d62df66bd1acef5e07aa88e4ec19f8a2d9da361fd7017fce1b8b6a91f7638cdf5e1d6fc2bb36f857bbabfe5f8e581fed7f455a7f7bb08;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he00deea792a3e9e5c0add542b68d7aa813ea38a5530b1313df62a9e264cc89a4269af8b5df0334a66d5c5c061a6c42e31657eb1ab892a671525afb580;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99b4362255a6195ebaf73b90c21990fc09202d4086b092a1c6e5527adee7463686402367df06933cbb19cbc6eec56d8113901377ac3a08b025860b42c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h738f773f7bac9d1b417ffd011cabc3736901bfa4b948cff70ac5025ba9472a5767918537cf52032d8f36843500a66575be67db095a3c154805b67e855;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc778ad8ca7a52b5bfef21bee7a3a9a1887768bfd6fd211fbcbfe89e7b4cc61838fc874f1b2ba5492c033a2d27adff09a16bb2dab6f3b19844db625ad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8993c3323259c35eee55baf3437f43b2532137ef5276da60209bbce9d7cb73616e6922d51580dbb51acac2e6ec62eccb9767b7ebb1c0ae6fb03d4f75;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha611d79fff31f0a3f311f456333d898c2335d3b9c0c787bcd059b618ea1839e11ab3295af907f8857901fdfabf05de2f975a3a00bcd5872b630f0a8a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he919c84aa111d53e9ab7611dcb921f711310a831ae63490c73e21f10ab62ef875621cabe02e26a0379b27761971cafcca3d9a7bf3514da099998725ba;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ae22e96ee6b9c1f1637510772f69cea3bb6054ef90df6bfa242ba20f7ca78f0df2b001e0846debd1292e1af7e6ad97a5b020cfd882045e98a7447098;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5dcac79b001d7fcb26679d7f17140358920ea2f2ec033e89aa08e6c5371dc6861578114693dea2fdcc1519cec8cb46ffa9491b581283fd1faf7989d54;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d49f9f77e09f8191394d013e87a0a695ea893fbe04b5ba75cff4a8efd663d3bb5ab35d7229013d614658a4e9dc99aff1a52f09fb75765090d1e54db1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29ad32d9d696fb4049e552c563193513e272d2f41a79176d9c15a3589af78d6dbc8cd015698c0178423f7a1881c2cd39d51d485b95dacbcfaccc6e2cb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h175114ae9d9136485e3d80957265240a85930ccf5f734467ca5fa9c4259e2ae5a61352b71468701a4bc7f607929961ec005bdab1a1ff6caf843ac1c5b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2b75fb76631bd58c14e5de7797d944f6e5efdee656c15fdb1630cf976d6cc5e92d6e3f60fc7b5d57c8eccd224a1d78404eab2174fae993e1afdf736c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h894c59b366e4734020153a6652546fd591a6572057322a895f349347bea4b9390d0dc9962a28904367d84e926e45725894fe90f6fa7bddee5aba35264;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab21d3fc1b938531d259687b5451b081e087d0666b0436ba855c4b4f65db75a2ca9d88d750dcc59aa9836dba0c04641c5ad43d19905efcee2addfa928;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74c05dbfbbc1917ee38500bd9bd59d9d95c4d3bf4f051855af47d6b715712f1db22024421f4c406e725297ef0116f444ba08da2c2c4fdf7e71241d43b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4b2b303e00e91b84b2fc0441a9484c736efbf4b940d3ab010ca3d3fbf23c506b4df106cadd86bca036d5d9b0d8942fb2632fd91d631c025a8aa87dc5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba52208f3729a5ded68869a575d256f3e1bf1c5e0a989c7c3caf0da8678d147d803f720ab6f7aa87a2b2cca4e5c91503c1ff70683732e47f4addeb76c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b70af82281096e67061b5488c9f6150b4826bd9a9c2abfe5ece90c2ac7f7f2cd0ad0613c23d1079e4135b960be664a8b9067bdde76042db810521abd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11073cbaae0efb4d415fe8153ac5e0b40197b4a7e909501bfeb80ceae2a838c4381054f4b7de18d8511caefa70780244ccce92b38812d0c7a1dcbeb2c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa1eea7805d484d52e032b8969299dab052ffaf68575ff3020603027adda89c96d70c6845c1ef4631c63665ba37cbde5ab703314e9e11ad5bc16f40bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83686ee9e9abe778a9b1436156fb7908de524f1b61632ae17d11d31781259c67156131f6abf8f6fa0d7369f2b3518c5bf4330579cea52559b6f168b66;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd996bfe86a987ae13aff94216e07092a70c540ac320173287ce97874c76393649f2cad76f03ba3142b06056835fa020997148068c49f786a0a16503b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd95f4b45b2e04e1d6051b1a0d5e092cf187ddf0cbe6861f72a49ea2462901c45977f08f22e1525c36012d3752f5dc7085eea9db53c55e1a0d578875e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcabc0594ae8760922959f53accdd9a8b8394e0faff07c53b91efe195953201bcc7fa08ff1385dc26e02b7cd8d39ac124d1cf342055bb7d3ec5a99ba2b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f3f6b40e413b9ea05affeed353112810fd525e24b68e2f5a59f569baff00af2da1b6f574488fdf429f04dec3ae4f79bfc77d8dd97da041d3267df65d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3f26c3faeb81bad49075be5b39adb6c2b907a00c86d61d767672f6a8093791b911e4af88cec9f700df7466beff06b43216384364a2112c32215f1cd8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff38ad56efffdcbd4b4cc28053d954cc1a74603b99957ed8589aef043dc11189ff7d2a99f57626b5aaaba53fb35e1d81b118777f01bea9752c83d82e7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70c27b67232b917f91b8b15f99d21daeab8ec18d1ee67aff36d74f9f7175c5546e4683987853542b487bad762e8dbe1ebf51484f8fe5b44f38bc8434;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfffa3ab2f3a1a043e459bcb241a357de70cc110f6f7867373577d608bc0b152a6bfe838286d97ba8c8f4cbc89af1d970deb22d96e03ea3191bd070ac5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h770e78aa103b8ceca7606ba6ad4e892ab1efda7d22a6a4d31ca82080eaf7cb4410c21c47a69036446ba043e9b2a61e4e92bc66200d87e8cb9cc6becc7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41a0e3106cf5fe889a46d1cb5ecc7c34b1a854a99d97917a7016b2be82572f9da280e721cf1bf31e7c6871ff59852d9e42e831dffd60526de20f580;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85fadfc041912965e76fe2c7231202fa00db75598f9446a6a89bd9761117fec87389181e0424105536b9a09e3ed281268bef897dd49eea4fcc66ebb39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41af6e81dace5bc8d20b6e577183d7276a58ef922f3d1622e29510efe90d7e30f636ba03459956ae72fac6c833054dcc2d043d8487181aec86e694d56;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd52ba242cd3d7f1fcad979ebb404b59d63b2ae4dfc11d5d723d8a366efb8bbd3c382ed8ef92ad2d2ba1aa2d2677500dbf9cadbdcc221f6b04dfea40b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h873aa0b277863a8c8dd093c27d13a0a5bd7bf897fe69df4da2f0e0dafeca3e82dbb0e6fbbc5479749004c717f7e84779d2e76908915ff93f9f5de3d8b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2eee614313d408eb0a1889c06cfa55a4f45c6bc407a5f4dc011fc0ebdf5b6b073013d3f0f5b6820f612f98173641488455298c444a905488249deecb7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfcab4a782119e88fda2c8fe327173375ad398b574d842b076787ccc311ef61843a418b566282dadf94c904545ad8ec3aec9a2e96a33b57960266332d6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20d4cf7260254a916e2c0e8ed94c9c3ef3d826eec61b37a43102c2a00ff6a8468484a4576f8d300acaf19030594f465b397f3613030b4684f022ce403;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2127b093241794b478d348e154a7caafe6c1498e3272ac37d62896b3c79f7964c12b1dbcb181fdfda6776bc40a15234350f82f2ac115a8eb833ea5b3f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed7251f814d8eb9fb7e921999034ee2a589ad4293f4649a7f43408f7581ad5676725dda3bd416aeab6830e0af22daeaa306d8cacd9779398004f8fc6a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22163f1eddab298523906771ec6d09bbd3510e8553a9531a0f5f1eee53c7bafcf182a90702a994d9f59ec38fdd910e009de970b45f7a5bbaf457accf0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a7fca67aa6c88b9f3ccbf57545873c675c1716ce6b97bed23dee16db838d17f3ae971eced1d893d46b4d2951228103fb4e7a4c7b5f942aca641d2a4e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3a0ed3c81f64ff08256af420b832e23c27a0543fd471e4edb043aeb882ddfcb07fa2c71469417dab33b15ccdd831a0eb497d09c5ab9d67478710f525;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60d1727b5341b9a2f0a341a95584a957d3ad938663348c112aca6af3fdcf8c054f73a3fcbe9fcf5d53ebbb586ed336ae8e41848deec3332f12831835b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca13fa7f8ed2372175d9791ad0710a4cbbca9b271afb97436b77be082bffd077025e38e4867dff762664f57fc8ca70465a4ae060c8e0e675dfe4d149;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24a073f8d0d0c5b062c91e8cf672142be3b28b687faa819aee532e35811429b2e76f545507a0290a59119261c4f2a5f22d756d7410eb9508b4ae79241;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdab44523187a3e457e338cd218d825176349cbb7e8c072ac014a109569364393b4adba2810bc118c69de37c352fb98b98177003d5aaae4701e587452c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14cef6106513a3115a5de917d7f341b20054ef4ae18f52de20dcf5e3868d0abcdc2ab67f8351671cfed112ad5ee3d201938b536d228cb1fc55644c4cb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3987cf656186b5d77573a5e91be79cacc2487047b1bdec9d419b93a32344324a4d8e660e92d692803990c19297cb5989b8e098ef9c6ffc08015944158;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb02041890246ebd984e72f26ea65af315f08896f21031b837d8cf70850366e9cc8b764cacea8143b17c13a944b0f82af0f994c908dacd994d704bfe11;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc29c168dc3d9a2601dc9678f130c18b3ce85ab9789ce2a9ba70c6b4def1eecd27ab2b2fca674faab665bb2e20e3304f9d3fcbef2b13e0aedae9b2d45;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d699f126b4da0597ea640a6d6c81e40ff6a9b5eb0f503442e7e0f45e85888654831a4a6086f4b2cfe1023731742478698493d050f8627bac8c9b73f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51557bce512c67b432839bcccce1a15abe0e5637c460644d6df8cb12e1ca20d6604bb4df40e3bdbec11664441dea7037be6a94bd5c1e79ba105f45ce9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8bb95f2f2233f39035f079526f6da20ac4507504ad5aa32d6be562e4beb59f58d53505e363fed8ed8ed7af077707d497e2cb01927f6e31060af65ad05;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h859066a24c7fcc3302068f5fcd70d1486ba9599eaace84d6777e7aeb919ade85ceb1a82720f60aac811f3121b772d7baca5de47fbfe0a2aa4501a4400;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2c9180edf7d602b0ff425f393ab905d2e30f005ca693096c65230ea67ee599da840505be839f1249a8298fd41a7e678d3f7f852fe585a451e1ae1b1e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9868ff0912af3e35b27f3c66f839e18faa63129386636db6d0f7814a4ad366f9492638974b896a1e1bd6260174cfdc93ba21744294e924247fecc96be;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2cf7b3782b3dc85e318022e61ef20874011147e16ca8b4e36548ea66ee03b5ef8515f90bb720e053f2550a529cbd987362b736b10d532cad0204cb893;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4adc3bd875d1bb7400a3dde7f324b34f424b7da25e445c21ef041b4fa9a0c7daa72728688d5354e4bc6c3eae85a3ea6093ad3246dad087e26f65b4341;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9bfe566e0194a62732b6c47a9758a0e3b7fea62caf80094774c04366e143dd80ba73c334836a98b8e00d69902a076119ab650ccbf8ca33a72c396f4c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89d80e335b4702cc4cee99314b29abda6f61c726e0b37da3a4ca254142b87880423322eb04c0213af7ce8bed254a300eb76046d0078e204c5eb2eba5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2658e9918113b1feb7c30a7ea399c58d0ee682557ea2509477f6d8e018ba45d93af5988a602c5f53db8af652741e5f111f430fc74d904e291e13811d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he015b2ec975d98e9a6cac39df405f9ae1a365f0bda54c85f10c0634ad6c2f9524b37fa517b2ca0a6cd2e1f163e6b4748f80e6dec1398a82beb442d4b3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf621ad4dab48cfee375ca1fd531f2a6fb38b2a9ef90015bbe6eb0820b365913cd236a0f7c1fef4dfb3973c1a29c973ebfc27ce7e45d3bed4e91978214;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haffe92a4828b7f8465b21ee1710583b99eb46587b24772c5cd4f0bcde0f40265a691f07f9aa6085da1b10779b621fba4fdfb78a8a0cb045bb7b576e82;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9c2070fd3c39089a5dddd1c4307ca77679697b68f8b51f57edd087b0f02bcf918ed47c21ad03f44e3c38ccaa3e7c320d20f6feac63d0eeaa10cbf643;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5847d4d24a182447864e4a9631bc0431bdb2ebfb168b12ac2af91b53687889e9337b8d84f0426708aa09220e300d46ba1b6e758ae0185a17c4e2358;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8ef2ad153726b8f06f85c5b294c80f672add58d1432380397cb0abe681cf1d2a7defc685d59d47c8d86cab61abb7dcf6f3653db2ef298e96d1441409;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc2a0b047d0bc64c35790b00c86887926d53c22bfd11610c71ef83a016240a8482c6c57eefb8a52a31b744784c6ee33e36e4c7e9b19f34de9423e572e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc897d8b41def0a7fa8c39ed62138e22c25a54343465c1e00af0a06d774b7596c090ba9435ab059bb2361af141e8bbd6d6172071d31e0874a4f7cc408f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1b09b408bb1602618795682a10a153f598dd59779fd67f848c20d7c8738371e7c8f69ae6d489b9bf44ea30dd0084e6bb174820db0aa8f4e2cb9dbc8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h727e7e5c2993db0aae965697501f1e01b5699c0068e9b41f18ff91aeda5a633c31cbf5b22972d310f0f199efb0304fda08e5c604bb924a7b6d7db6e31;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24527740e9238fc55e1fb0d0df644b7518a3c8ac8c1b32b87fdc7e8f1ad3016707bd486c36562b25b397d1a8fe5087a9504a733937511ddf647ee1fd9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17984e175af1f3d26b741e3e7853d5c2d3b26d95ab177d37557d38e7215873ce51e8ce696831fcd763b2b13cd96fe755ed1846a5c40b96cb8e51d9c96;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he8f9c3493dcb4c8804b6e6538f651ba9f28fe78be1800fc923a2bc170c7a3670396659fdb95c9581c3e45e48f31ea4ace74c9d14ee63c27bdfffabc6c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11d6e00841b25dcdcf7c019afbe73b77d8a9cfc8298974ddb87c2c9df54e715b65f4e40b04a0726fae3e7f3ecdb04a085f5f5e46ddeb0c512b11a0fec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha451bb29d5300a004c29332892d40126ecca09636ebc888a2c1b87fa62d7bc2ebe5a02fca49d07e8d41b5a42a0bf0d80011bc283c6f2eeb38296b7148;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8517b3cdbfaae7578d08d60fcd86bb7564e13dbe8f6b29a5c954184936a8df855adfc1952c48314445123a58c07a339eba308698b62ab3e674463398e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4958b937ffe07a7bbbc5f1581730bc46b2c948824c0ea9214f6622613396efe98597dd97d4e3ab49a5060e889d48180a4e2438867b2d549fd9724dfbb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h842feeaa16917c0d6e70affad54710a57ac2190df8ef59397ae143a733fb0bec3b6af4a3ebc3a19b81b165b82773e1155308ece143987e9edb74e5f6a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6ddde9c519b80adf131852aaf196e0e40f0f8b3f7717c77a8982c46c23932406c6de4008d3ec171c95beffb138393c92eb9840219d93f9faadda07fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab3a6bd2cfe016054d252d6d9de794b936dc9dfbc3dfc074800de99f871c655eab51c4e99572f86dc0ce24b397da3f45ad1e538e216d654784e04d5db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47e11805835f187520a3553b04802ec0d2f5aa402a0ba0d26442f53e6249c9c71598b7be9cdaf8a851a0e81d0b0044a30ddc4627e3d4f7c3e968cc377;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4f20af32bfea534192959adaab1d2c2e3dee9a71b6981ecb766b61af949ed2798b2d9b59611e42126e9d8165b6c8979a059cda69664367a8c78a54b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c0932c95dac9f3dc1e223b27c15c0604bc8850d866de0fcd3b1362ad14391fe8d6b7b33f7feeffa95308a106a2995af7a40a1f11e6bb36f10b6aff72;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2bfea8c0a86c5fac6ff42e10bade8e5ce0b1469702ce8809f8547a3f91d2557c2e83de6e6072bda5d8922edd4f8c29303178ff8314cf20d704a234c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ef7fd57e221d4c2e8586dfd467831a5ebbf48b9bddacf4bf08a4f48e9c018015acdb0dd8cd26603f45e3b6954b568a181160c2ae694a6537d100da8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4357ba7a7a2cf099e7710f995bc522a35d31cf9eb9ec504b5cd2a0ebd621493ea0186be8afe2c355f70fc7e435319d0592fb22cb5b17acd458ec2d4fe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4852bb455c1fc4155bddc221743f74ef34d4bae504a15db119f9263f7e74c2af21319599cf914fb081362a45c08b9739a21981b22a2d175b5058013a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d96dabb8d7686720fb9e26fe3f21b5bf49655710d67fc378d2fb6193c8ecfa7555eba7281fc66ad49be64010d7c7978f927fff78b0b4d46f4335b0fa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdeed433d4bae44c10f02df895c04d740660f40525998d469c75485c1af466a542c24eb505e4a15fe01fbbf32310ed8d5788c94a956087fdee540031f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e030984e245c5748a8b4971dfc61f9b020967ce797f5bec1487bfa7bbcd4efb75d4217ba6f5055614cdf7a0f1af7a92c1ab435d2c05906d809b4ad3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he33309798593da853f47c478daec8d396de1ff8922ec5c30ec48c79cee32f370677e9ddc40cb033683eed271ba35de0895eded8f75e34c6afe3b35248;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82b0e176ee850049dde42c7d9d9d0f34d863fea1ea3e4d2bb20c3e5c161aaeb75f8f98ac5cb73ab8b018eb4fbff613c01c26172d58c5f26e5d32aa1f7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6eeff20a6966cd393d6273b24cb284b2220c9c71527f9c5a7c4651d900edc3f0ac96138437a28919b070cf47b4b53bc820878cef3a6f52c337fb027d0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2568de6c62ecd5790554bbabc2d9a1dee58dc7341591b64f4aab280454b76f887a09e0bf6168c8b7eb91bbe6d2e8b4606300c66f366b40cc39774b984;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6e741603b52f5b96783a9336408bd97f5356640a6a450e787d91272acd80cd42eb8ea176936e8d9965eac116ac40735b5f781831bbe7c7289e330e13;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9fec1b2e55939e6235deb57d19f13659d8dd222c7b70270004aed5550057c5d7d4c0d0bf96ebd8a05fc2a15229d17912af1e826be3b43444b1b102d01;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43574e527da3921f4e28a11cbb3ae42ed983cfb6788b09b84058e1a75886851ab8769e8e26067835a80fd2eafb184c4b4d1f330d2ff5dc2a0133b4fa4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87a8e8074da9ec47c11a2f7a715185b9cbe3584ae3e09a51dd1a0e5342d1e8680249d7d89423db0bb7101965e2846c1aa0aa08b8c54632277ec7ebaa7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95d0840aa86da6dc537780d2b2c31640ef194e798a484af4d611ce07c0978a26077588146dab1aa9d437cb249ce700cbbe77f76f324cfa7bf38cf7240;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e89cb3a03aa4c52ad9d692c5d447719aa4c56e8042396cf0d531a998326ab5405763052c213091525d75b45a35c376b9d00a7fc4bfb896536b76c078;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57fc395c6932035e1611d0c137d54d17b660efa39854f0c5af985733b6407d91a5d66293fbc1e7a5dc7b11e9aeee70dd2d210658f800eacded681af58;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0f6561c6fdd8dfe06596f6f3ca84b2d2a02aea48351c4d354c7007951c55fe88c8918c154aadfff787e73281260ce6b6419d2091feffad6aa6af2fe9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90884c4696846ca71f7cadc208ceb0e99e7efeb531775d3d7c8a0b62fdd1c99a28e9ee2dd1f428bb80b26b00eb2493dd5920c36d164a9af0515bff77e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5659cf178f4bb3b4f28d872ab0c20bb0d46463a77967f0ed1a5a8fdb892844e2a73fc263a75a1240de777d2df2b46ba282c83e79cad2da4a4cbbfde;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7314421fe668b937a306af1c83f1e3aefae18dca9881c3f9da175134ef6fe8c2c8e6a279555067f0d8cd59bc6e7da55a31672988f81e8af69be6af5a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5195c50faa5293dd205cad0e6e819978a99a506772c51964431c78f0e2895a63e1035a8a122d4feb17a12e353a757be2f9d0076654d27133b969519;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78be73e24e18057f64547d97db731a341236ba3666924684eab891ef10b1cfa2d706f8ff4e8b6426093d1e4b7dcefbd6eb59935f40c0da405f126f123;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0f6db7c22066c0e50fe63fbdc34d7bcb00ad015b4ef2b61e6bd2fdf10cb2509de9fe6fb70288eda7f3d6c5589809008e82c284b177a47a706721580f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf9f1fb967e9fa035955057418effc0620426f51b1f3f9457a4dd2a35005f8390ed284c7d833fe6e993696e03c02addcce0bfca1710778a3dd12b8e78;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f5d28925c06097bc9c14d509d3efa15a5e9f181c0bbab528bd2db4c180003ed48a9bbf617b6de14e7ac20940d3bf989c41503e10ef3b44b61c36d387;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81bb9b32380eb6537ddc478e3a0fa12968e0aa685b16190077478d95e92e8e688553f43fe979271dc191cf0a1310b1d110e6e5fc69e505f8b4bc76cf9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ea05f522ba3d04092cb9dff12abed4d408b6a8e63b44ca6834e25da9aa5c9393b4962739798edd94a327947ed27d5710eaa5efd3e24e03b18ffdfc31;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h165e8c525699efc9d32fd0ae438c5428858ed0b4730167b5ecbcc8b05fddfb223c0648f89fa37bccd796194ab73e04a6c558f523fed6c7136dcd43419;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e26353e3fdff2169b1c9ddb567b1307993d5122c0f164d46dbb5f11e67fe04e1fe80fe515680aff8880ffb3df02e0d1fb4114a272c7a0725ac662d38;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d2e33559d8a1f4ce87eb0c0790d7dfe8866fa8bb160c1bd0feac094d6816302036f46cba74377c32c2e51135c214c169c14eec7be5975373ba667a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h567a7bb242b5869a6c388bb4eb1d0ee363155abade841f692334ac9d422fdbe965168ffac03e77dfebbeaacae7710018ee3ef87140252d54db9c39fea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a46a193aca8dfe30d7d49f10b51506c050e5329ab25efb9540bd14b5a234395f68a23f4b40d48ce2b3f542464ef23b6264e588790e3a28f37bea517d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0942a6ba820a690afae8297c3536875104ed9d9d0d50cbff2e8f189f59f1716c9802b86507d479bfea4be2ce3563811372d6d3a4f57575469c7d19dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had9f01f7b8624bcedb5b885ac91a4f78709cc127b538dfde5eceda90f1f3dba8726106cf102ff3d0fc9ea2120f8fa41b143487081d5c860fe134c4538;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6852061c33474b49f08f0102ef257a38a555e9391daa73b0232df5faab60c4d61bf422d9dc217185cc2726b4bdada8b2b1c102065adfde0183763493b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e3a78e27ea4ec5e3d4f7a21c440b3aad13b643e4453aa12023708bbb1e632352b4382f2c4f4e83018e989fe3ee1fd1d5753789414591add11bf810c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2fb957cbd50aff5370ff48de3ed848822bc9f7e31a1735e5f4f4d4b3c06d70d2126a2dc70453c13c0b85bf8a327937672e58e09b06dd28ae0d550bf7a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51b879427ff33177143061760dca9f164af401ae401d6fdc564a14d7a5cc705f9b48f07deec9937596af7fcf972f6daa08faecc5ecd6f9c41bf1b840e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8cc9915322104147e96be03bf21f8ed6c93ace4dd64892a726c1fd638cbd165dfc99c60129d5d3f2b332286fdf08a6270c0eae0b40d49c6c61c5eed6b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19222c5a6fb13a65628131e66ed8faf4b1bb4b2a8a326aa47dd8ad096b05343f22a53118ade2d3f32e1be44359a90c61a8836ea54ac26ad2ac6c1eec9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9dcd75028d1984793d4e2210a7a1797aeea0e68b58ff6894a56809e1f9718fe64e8ef92e668be36df2ca354aeed8467e730560b83fb860d619a47112e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee25e961f2fd6abebc06228aaabb3e605b3e11f6245e0d1ec1cb7c1cc9a1d18e16fbcbbe7a6c007f1205cc13213093f8edbc9c1962f21f59d1f880d53;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc2ed30b062847ac600dfaf61d2f9ca3c82969cb8062aa53dc4623d47454c17ed322354e7bbb1c8afcb1659245418ac080fc063490e3845ca213c10cb4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc75f4f807eae36e851b4f7be5150489576420108f7b5e48a6c4766adad740cae82b13970bc8aefb8995a6135fa07509ac1b5a2e00b5249d9af74fa496;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ca5d393e003b84c9f124808430e18c47099c169fecf52fe9032d01c29265e88e4bc7d4f0ac36b806bb3e0da494a464378ec6b9e94266c4c18c6f63f0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f7d9781a5d502faef09f82588dde8c666b2193383b7e839aedd8111a483048b44048e7cab2bcbeea1163ebcc219b3a8b566165ac1f69c7147653ba66;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e944e0c2cfc407dc423e059868599d1835fcf7a4914fe725fc1b9118542e1fc42a0d7baa4c8cbb12d492d7a5c9aa6cf354a20cfc436a4df8b3c6b2ed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha353dc6068a35c34f5effa7f68ad7738666c8d9534ac99d1f7c07343b84961cda03a7e7832b73edd259ee1c7375c4f08338d93a174eaa98928de48dc7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba8ff73b16e34eda933a2f7ab0d357c3a00c8c38163fca52e010fbdb848974a19fbaa08e96beda78c557c8e722af54ef89bbbcb04ffcd82ab5fba00f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72adaccd5eb40a70d544f3bf88e4471192ce6fce6e740a73907ededcca34692702eda5ca407175d2bdad43f5737fed9932e090426f4d1b7742a46ed53;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61a9b4ffa0054363a9fd093eab6eaaf4b71154afec84761effbe008a07f52433e0f72bd35d4305f4f588dd634344bc085cbb21aef3df33dd87b54464e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4545701e569b6d22e4e6f0265902db3fede6d9ddef708eb96af2a7fbfb712660a70fd15f3c418b582afe8f2e90fcd85608b91b6b23ac91a80e58a6ee0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4e50dd18d9b46b9f0bc9f8b48c8c9dc4eef552024d8aad3e6d53ca3f0b9066840e3602ab59d0ab7ae8887efd8c5d5e5ee10a50bead744a62ac0c6e03;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ce8c96aad1b47e11c556b9e564304af0749196dafd5e8fab0d4499ccfffe268a301d6435d72599403fd94da9a691b65a7e32f85b107964b1d6265911;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h168c9c212cdef40a43c3bedbc997f82375ff9bb3b041d0c247f8f6d14e5fcf6088d701f6ffc01c291e23eb467428c8f34cbcdf53721fdbef067aaea8a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h550a734ea1b814863a334f13b5dc2ad6e1229c1c18c32df4942ce4ae996851501d89eab457c8b0e011beb6ca21f4d24cc8e285c6de73a6212f472f022;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2e0ebd1e0725d22807d86d98b30fbc9fbeab927bb5e3ea29599c673496e26383420af9b41dc7b3e1185e6651cb036832d76a2c59bd2f5206cba67f5d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc136491316f20b64aa2764de725941b40c3bb098dea23e92ec574206a27d9523e05c303218f2c306ff8d14acf1a497e9d81a6a54c2be0649c17dcf5e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35237dcb8e4c477768255358c7925829e49ca859152d62061b92b5360e6c0c78ab78453b94e62c9387e19459ebc125803a0d643283f1e23faceeecea9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf21970ef4234e77432e72be1271356f8891ec5c373b30bfe8ea7334509f1e995949b83c96209e1e94ed1abae907664293cae6ef3ceb77e42a2227bbc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4d8bf6550d086c3c2959b8a970fa57936c5bc8073db242d805a6156391e8695685fb9e1b95efcc1a604f21d082b9ca3c95a6216f9b89617e50c3bea7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26373e2359d0fb2d7572901255abcd48c4476201e8f5c0ae3a35ea8c177150b294db80072f66d31c21f777935b6e0e86e9fbe2394d1ac7e2221fc93a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e6064eb5dd14f7f590a7b6b93e27219f50b9caa78e4718c7d0eadc2b18221b8533b6a8bf4e2bf1aebe71170b5e10b9288f2b10d43bc9912fc73f5264;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f172ad5681c9e9c71c2c7bac64d5acbf159ca439a447f57af0f2e178f54c68df587630b9bc90dd6bbe226926cdaafe0ee228cd33b5bf3d7632738f19;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4dd954c4b7771b6a777a1441ca7ef6ba64dbd751cd56b2f8bf70b8a17803bae9f866863dcb802f9b1984313da0ae0160b2df1b74458d766009dbe33a7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h373c3eb4ab1ff5c189cd86efd96533d4179a0d2e0f10c4c2a66fa935c233ed720e0066d1d8a6a96d817c55eaa825ddefa302ed36f89e2f6f1df9b69f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd10823e795e06d528ab68c7126625dc1b4df9c73a8a11a6a2793bd340a40bacaf8019dba75689f5cfd5ddce61d0569bf6740e52073e39cc15d222dfaa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78ffc84dfab3e3e06b782b211575f4f7016f4acd2d6f1b73e0bd6d6c052d5dee7be9aeecd72d9c4e457f3c067d981f1140eb8ecbfb9d1773a187c46f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc84e9a96e4648c23c317ad22a2e7eea4f1f3553f63656b44b5d918ffb963a81dcf6dad8601fcca68ca51282993a7506a4f4d9b361688cffdc89ac0dd2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92fc57557acb52ef2b143055ec784f63bcb11d3bd612183b61ad3b74ec5d7d5e02a7fe55ca456ec3dbd6042bce1795c8af75013451dc0c09f962567c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5983c32ab327e37ae3e73fa48d3adb559d84fbcbc7e5b94110629f9c635fe3eb26a7a3c4e998b50cd65fa60dd00582dae895973517cc98dfecbb797f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5d6dd1f453e38922cacbf4fe834ba2b56da0705364409e61c67890b5ab7c1e80aff2031bb95e619e78c1ffed646958c3aabb7d284a5e9a11a7568d83;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf34336698cf788e5b432affaf0eb3568640fd782f0ae6f80765912c7e7eac265768de0fd8fed98c62f62fe095d017674e777b08562ec0fae9953c3d1d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4c97d0206579b6fe354f94bb21200e6c742dfede85e575a6085ca53045fbdcde6ebe4643812faf7b1ece11e4f0350122fb8d9ac2ce733158b51ee02d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha256a124ed6f2f9f6643aef3a5708d5ad90d663e308be01de0579eb9b1e03abe25915cdf17b9cbf6b4127a5e0b53037f1c33a8524dedc4e78f93fc484;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd02700c19552600fdcc54a2444b2759bee0ba6a146be259bab27e0d8fb60284aab82f1d09b9dfd76748bdb0a6abb898007af58d3852d434edac9f69f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3529d83b7cd68cf4ef31643d8305704c60ee6dc7689f3b825d527d58aa191c18a2db7307f2180fb9812fe1d5baafc735c6ac4d857aa0bc059f51ffc9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha6708f647ae8e7ca28910ed5bd51971c3b0c45e1ea9e5f49105e7ba7b0cefacec561b2535da8a389cd34a45369828b94212ff2504bf7884d7d6223263;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4af508ec0dd06581ee0c7354fd046c9dd00395bc7f37166ceb8aab90b0166376ea427930bb17cf9a13c376e877e54b8dc473cb2c9878275adb1cbbe66;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf13f90feec9f21aae8c3e9456fc02635e953d0ee3308390ead3d94d6dd17ae1e6dd4e6df3451b0bb39ec13cb0876feb22c7043ae20c15659aed9a4675;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9688f560d773543e06c7315a62e3326ed8edfb13a9244aace8c179f573a51f05aaa4a3c531eed1d6db7147c2055e4ada9be6848a19e64e17e84bc8d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6e8f6eefe5fe79a9472d16da69be5a3402657735e7ee559e786e61b09b5d2c5b240806ec2c3582644361432bab5cfe7dc1d830bbc0f7555ca2b4647db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5360efbac4bdd0f56eef87b7a7f168187aab45ce58cf348779dd410d67b03904a6de14ebe340acef685af78f7050a0da3ac296fbf935eb5e50d7b5b14;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha54f773c4eaa247d3978c53b63984057322895b31f92b3cedc8d5299db9809c09bc01f67db51d62162a59e0e0b025ab1775acbc1e7f08c6db88520c10;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7807d8817e1d8acc01cb4eb81979bdeab641624b8129bbb7cb7678ea78b5127b51afb20463747766bfb652bce727da115634d2c9be83002b0b215a07f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4be92c0be1718b9372fb516d4e3cf354d57fc596d659405819502ea885ef9a40603bc2968439a744b2357f1a2f5a14c5f5ee79391b7636b3730f8dc2c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he1e184c276551d4ea130127da53ade37ab9fb39408af05041947f17565d4e6a0c83d947d83c372df3656c49e2fe1524a23506466261f2a0a773b29133;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd75f3cc0fb793624a1b68624a1630cdebf3a3797745f125d9f661f6f18027417a7382cbf37a24d6eb5bacb2ad8e82bd1116817e47ec243e75dbc81ae7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3510962a57412c8152da85c7a68cc61402c32a526abb3df90d9fa58a18a99d68f22ed467fe6e946681718996f842e9a1d42657bce5d9bcbf5a05a781;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae11499d04f0c939013cdcb29b26094d11b16f15f000d9952e8e47dce28176bf6c1cba17c19a865b7506237bd807c0c446088aebb48130f84e8924f2f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfbb8fa7fc674053788be40e8e8862af15b1775d88b94e49d22501b8d0e8f88f955272a892fd9539fd7347da81c0d403a6db5c1299b92dc76e12b6a986;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5472586b4ab9b2dbf378109a22922e6044b32ebf029c0eebd2e8ce27ad1a6c48443e793ff4848725d270282ac428f38a430df9036ef40795bbebdb816;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27be8bb90195065bbaf67e55fe4d7f5a93a77b29631f3045b57481e0b8f3a9fbabc804f5737d6737e56eeeb7dac678f832af94d714e1494944e503740;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd5d0dbd56f556dc81681aa61dd6f61895479de7d5d407fcdd41d064e274ee4c2602b06e954d0d52ef1f761a13662b41bb94e33e8d47729ac10ab4c105;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a3296e6798c979866d731f043ed74be6953cd4ae30573d5087cc5eb5b4cb99a9c86932c5ff8bf41bdcba6b7a2ba115a312628eced2482cb44d05c297;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2132aa8762cc430a1a8186f7cd6a8fa6def1cac7b66a18faf251e3ee66046b7def1e5112454c5a278150061e4b5fb7aea44dbe2be0e0bc829e946494;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66ddeeb68bfc1c5e541bcec60d63eb3173e2d95bec33ae27901d54226163835844a307ec1162a54e88490274ee9cf2bed7aad68b1f8a204cf730886c6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0183afe54b7c6d5c13d1ac3c57c7163071a16e2cd50cd996b448f0e89ac8d4ba5ceaba0aa4ef292fa7ca683137756ef35528b64f190092264d16e5f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf15ab53d0fbef56c38ba67bfa77c44dab7153ab627285825b8b73c8085c9ac9ed5d2c24f1c16b3e21c654d01bddd00f7a1aed95c8d3f79b097e02521d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4054962419f80898ad08192e6655e6e3fabda8cec1d26ebd7206ae6125352c9ea985e1e30c517491d74d1077922ac00b932b09b05b770b4c08197a4e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc699285e8f3c8044630501d79b4b83e52c9e72c72b04a53c24ed38d1eb4905e455bbe3834324540892efd0c4702df5a8ed9773d7b3caf47cfe72b01ab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h357d0702edfea28c9e8beb413d9ab7d7fc4f8002e9e5a1f67d06e455d0ca3de875065cb488bbd994128b414e0b1f87dd93f2c0f90b5cd437ecc65b1f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc799eb4f236c938544f7bcaa2b50ce71c94cc5d0bd716be7bf861c37ffea600cb90bdb5bb5f83833c8a87dc27c29474596d0f55a7dff407a3d1d3402;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca3e2af120853744cd9a25ee16b03ba6a1c0cf217dbc8420f076d2315d49ef8166df6cf890ecd12941279e752e441a90acf0c27284ad8fe7d2934ca72;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26e2497e1f5f9354f5693bb0cd214325c5adb70feafda6bcf8893aaa35805675f901af315b1071ebabf80686e1b4d18d5aeb9e5d9e4263f03ad61eabd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha099bfb396e4f78a1063cf8ae8e2a9608a7fc7bd26a17afe83ef0aaaa93959c1de668fb64d4240906492db9abf6ed9f6ddb91e0059ebad746e15b768b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62c39f2fc0ae49a081f2ed09ad1be161435a921e6a34d92c6b8c121a7e7ce48270c637446c9cbf2dda599ed252bdc64a369679e5380ad1f6fa0be35dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8937d8134e6bb1060df812bcd29da2521ec033706f85d594fa23fecb1e1c2ab37f5413ac485289ea4cdd2066e5aac8a57db3e7ebc1dbe2ab07f771e4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6dd78eeada86800e360be8b74cd511c84bd097bf5811a071c4ed2f0adf99899d7193080fc5ec020f40020f0effca07302617d01ec9aeaada2095d9cc7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7dc62ac9d382ca26eb47a367b9c6ad35da82b02591059331ab562fa27c8bc4ea117c7f9ba988f7946affb20a8874ea9430c7e7eaac4012656535206c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50efedf387617e8303b9ff2f6ff6f0f303b3a163c1552a480d5ec641ecd5bb252e081b228d0ba5d3ef7e34ee4450d7d09b48e068bebc4bed4df7efb64;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5779db36dec05ffb109533d814f057cbd3a395450c93bec6281e73c745df881225eba8ee373b19f9a60a161e6ed1e860a2e83104a86571ddd4c49931;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h368fc04bae4346d56c4d59dd52857d669de8b081cfe6fd38cd745823fc27abad385ea763cfcde745b58b188e225b4eb33d5e5094c82e12cff87d9277a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e71c92369ed96da65565ba37d981df5ab27ed72ff0f744a02bb4c476a549e59733e95d8e7739feeb8c87f724b51b7b0d5558ff1a287611bfb913c74c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85d47bcff83a2d318e2033feb01261c54f8b559fe343551df7876a628261b9c69d779cdf959f54ac540bc10ee25958f3c4b82990f5901c871d4e6a48a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h455167bd0baae9396d797c95426470836dc077989ba0536fd19d91cf42c56672cb2020d1d41e8143d7e3d7f5efb80555a16859aff45e728112175656b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18e04d152ce6dad4dac59f2f06d819846cab3897116da297f27e87be6ab6877a80a94f8ae2e75b3fc2e1fb5af0caa9d50f65315faa95af308a8a8d7f6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h412f3aa72114d11d2effb3134cf849c19f963c62c4f231737b58c37145eada62c4e1465113fe06c1fc73503bc58cb9ba90fbb6e5272b93607619398c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6bc364e5e697a73a8900172900cc0f4ed9401efb9a046836e8fadeb77fcad874008fe5b9805d989a008b06dc07c25dbf6a13a74ca85edaa5d19444275;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ae06f1351c8be6e513a8e0ac10e121f22db0b21a01266e93f689c3efdaaa0416b6aa7de1b5330bc671e1e96d9ba8770a6ad1eee7bb680ad2ab09575d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha48fb14b857abe857c385b297ad820fa2a207163f52b520c52ce4b66a3db0c753b492071b39f70293137a38cfc751ad71747533b9863af225039ed448;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd72804d8c02b7d23b4f83bb80c8d025e3a53fe4705f56ba2c3382f4048d115f3b13cc99dd9e0613158b958b324474d2f01ac8c7220b9ffc2961aed546;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1af8f59a7c9a29778bf1f6fdba8adb6a387e4c18a67170591ed4d0190ccebcfa5bbd13427b1ff81e98781b0f86b2064bd53870ebbde0cbb1e8dccda61;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2794715b76f2d76e1c80e6608a250d733cf5b507fb9313a589aca9e23701097e9fdbc77dd7d908345061d6374d8b221e712fd8afa65338803b138b1f4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca9c9ac8c989608dc03c2e291e932c37d4be168c00577d2edf66d8d71d2009781fa454bc5bd33259a61fc7eb8a3f7a8da370af38404a41c388fab7e3f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf291b1cd4c5f4eb82213cb916e7a804cfcdda0b55ac8ac1d256d837ce3deea3bd273d8d1d25ca0948bf0823c6505d74196ab135e0c85ad6050355ecd0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4eff1471d4d6810b2330cc636c6944acfea003f80ef1850a6e7c63f5885b6298add33887c3166acb8db6717af1281b7a9d53e77d0536698b5a5593542;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61cdd3558a53102e3603c104a21d1390e5182fd084c045c1d9251acd48696acb7c18cfefd05bbe38ae97c926afb065d48a788a4235c17efe9dd0497c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5540c6160ff1e78f577202e32e0f41c625b5bd7244cd8b15c2e326578681a93f90b7e7269b9dbd8e23cb1fc4b458a25f78000420711162fa4097ed826;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94fa46a635f16e18fa474fe81297e13f659df479466f7bb19dc40f1f3ca5a3ba61c95ce10b7bebb053fa010751f934a2fcdc02f1e711d0874609d833f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha08fdcfa4054b6a5cb46a4c5f1c96c2b2bbcdc540ebb35652a59e88ad2c9c8af5f377af87d7f9f5a4146b0c3acdfa5d625f3313182181ecdbf9a043d8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e7bc3059fd71d59a1b553a9127fea5be314a68b7ac4b63f692b5ce331d9fa7d64666e62e3a84dc1b0072ae94e5bc09257016ab32ce57b2e13fe03fd5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ed6959213cbbf56fc20ba32ab8c1547bc69c6a12faaafcb80c3524d81efba37223bdc5226a79dfbecb07130ef9906419c4267c40e78b25c8f1e74ab8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h668d86411dd441d77aea636bbe599c0ea8b24614ae8c77de9b9416ac68d1556f4ded5d0a0ef65b1c36861e14c74a00f33a9cff6cd8440cca3b65c7980;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3cd4fa0166291c4f062a1f347c5c450ec9a548952a65a42b8a27f8c9646e10b74fcbfd2ff69afddf383b0f2b562714648ea01997d2dfe878610ddcd3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10abc9cf9f9ea0b43fd025d1c83face73beb711eb87c2395b1027e3c593aa105094498983b325d44774900ea3611065e32a5a204439cbd8f9b827f57a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h24b3bea3a1838e3e4502134660d602aa3484ad4e354477b66ca09dfa95820a842923b58c0d116a228aadb04a877366d66d98868d655711a274325cd0a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8bfda66407cb25f4e59e6965902664b136cbd9b217b7bf93c706e12f7c212d82390f662e0ff1e1f3095284ab2fbb74a40603bdfffb3f1254b1dcd2b13;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f9269a95712fc5ce10577e8782affa96ab7c5e172bee3c3daedeb03de70aa509d7260dbaf4c57663840b378520b76019f958dd8d8098f0b6d1758814;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5fa619a10b820f308b3a1d9cb13a9b960d2ed28dec4978d9004c0e12b53dd4229d8c792a947d65f752e02c4ce9acb93db2d594f8e33b256211484200;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c0321b27b686bdf3ee305d44c7aa51275e4dc79b8e90686f6306e530b542c33aa4ada6c220b52a28e4a8fd4f0b3770823e38c3e9752b2984a3f825ba;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6e0c682738aa937aaffef8253c9f6a7b519f5d82335f2b9be70296bc4300bcd778253d38101eb35418b3ced812da95cff45f95b3bc228c2fb7df5552;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h982a4ee0809820f88d4db3254d3bfb38fc1762f1beb4f7778c9515565e2011bfc370fe9673ee2ee69eadd5146a23683cf15b0083955a63b837dc852ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27b3baaeb5f024011e982c825f8b28906d5c270dd26b249b70a5d69ccec0ad4520e1a97d8af0c1064645532cc61568b607c3e078cdf8aa6f60b77bbf7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e38bcf89a3253d9751ef3b3f70229efb559002cd3656beb93ae84f541c4954e77070f7d703d5e4396cb921bd5867fe32237f238046b25cd278b690a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68b799f47a1a616483cd930cdb7b4c24586747806e13d7c692b3ee5144f4f2e28cfb4b27258782c95302cdd113ae755c50beea93b6fa07a8eed09bffb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf544ca86169f2a9e4b3b8f70470556b07e0af637726af3cf6142dd60af8ef3e2d20b535d9475a7b3e25d95d08c5892ae38da51b42fa65de9cfc606d8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf1756e0e1b31e7ac0acd1f7174d266520bc62e09539a4e1c4dd13cc42b9f6c9f1f36236635ceecf8f07522c0eb7b86bdd249d00d10c04ef8691391877;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b6a37110910efd8f8f6acc001c9f550f352523726cb16571b726bb458915249cecc0060b83c7f7a022407279b0921d1f0a4979742aade94a0b74899d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5969697cb60c31faaea43d12360b2484529999992a6da36f673b53c384464050dc4645c21146bd36447c3bd81342c0e5de7f992ab22da048a3dc76263;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had43554ce99286da6cb25ea401cdf4817eb5c2db659f0d8cfff372353225e9cfc4accb200d91294c17922f58a69d60b3781368cd79da34449897c7302;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf034a1ae3335cf741c9438271178aabdbe2d1224468042287614eb9076aa43e9faf629184f426dead77b75d6f56b65d840480b31a6c26f9dbec614c85;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f842b1c05d89f5c0ef6cea481a4fb5bf1bd8855258894459b4eb139778148d318acb3f5a4d79252896e0813e5780323c47622e13e610670f85bf57bd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h41d1a2591f9bde4e7d7d2c0a4794199829d55cc717372e96a44ab1979a00d61bb0798c99c810b9ad41079eb6b5753fbdfd3c340178af3c3fdade93e5a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5978735dd54072c17f2b82da59637f97999fbeafa939c874ae7f99c6a22aa5a307cdc0d461ecdb2857188ad931854fc150c94be50a67f3401cafd4652;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h439d898a4a35a8cf853ddc594b73c3d8f272dff8cb31c73d80e29322b180267e4e88c1daf3b86f7f56bf9f43829baac34939e8c472d6f1075ad31b1d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h188d8db2e2496b40e6bdc2604fb8a4ae0c3141419362a9d682b80325547ebb6caf3923c44c8470f8436c2fe95b5973849906a17e878bc782954422d7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedb564086d686987126bcf63435860cdde194f3aeee8d554c6344f41190282febd76c239557fb43feb026a6a4f1e5e6e899e9636d935e5b8ef0c7d30c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92cdc4965681a7da37aa37a87a9e95d038ec026a0baeba9aba58b6aaa1e3db0fc0ee524255543ed974ffa9427788be784be90c041adfc6f77ed3bc2ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7190e37efcc3478a6d6baf731f5698e8a75b9b4f5b24688defeb18152a4becd6573f2c619f366b270bae04761dea1d9a0db82f14a105d1a88151f4788;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28ddfdcdb771daefd1593904e54a2370b58b9e0b240eb74f4e13d0843bad593068a0f9351a88b0482d02f5bb1be742390d733e8a77001b05e82a13cf7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f023af2733104cfae16540f7f3b05ec734923d69433bbe45fb43442dae181aeb8e93defd42d721334c7f64140331f537c4f0c01378658aa2c2a8da0b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a08a7dfa12f9b2075ba104dcad25b1b0a3245033cc3209d0ff9bb6492cb2f17541393f500711a9ba1d9d61704fa264fc389132ecbc238b3afe468572;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ec4755f085dec8adf489e8c3fbdebd1e867ee5c24e03fb351521fb06646bbf2df4f44fdcaa2e00ba345ceef6c604d3fdddb80be36897b7fb21c997fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae64e8bd3e986b5d01a4603509776ce642e3b26ca754f26e216aa50f389f3c91ed75442e5047da8ca2d2d52c1bfda7caa9d6c77a755e3a85e4190fc34;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heea8e896d6d2e72bf2c3c9ea2c8f1818f6e87aa035faa27dde389a2a27a29f06a74fba527727294d6c6449822b4f38811cf5da09ab13fe4987cfaf65f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fbf710bdec0028f2f1fcadc23e09642206c4f591415aed5083ff5e001231a7d0432563f4d5c884845a07eabfa83c19d88bef05617eb84a72b57c2ef5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc60c5be54e1077326cfcb9b846d8eaf13bca6c7b8626a1f29bf7c4dac84cd198a31819e71f9d7f944290a5174c9a711d28a243fe4ba1225921655d0ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2df8248a1bd445300f5e6cae1ca5940d8ba4663a1e1a8abe6046dbe3ef61eeb797c8aa0ea5fb486d1a37174256bcaffa2d671ac2c96199e1f90a1b363;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf138e91860b38438db258c86177b25eae65ff6c32d11554af9fe9155defbd6fc46e2a2172faca37472003e78c6d01807679df359c84f7571fd8aebe94;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f7d852c3e8e443bcba07c859ba3802b9ca0fd241f2d20eab3d2fa19997192d493984e38df6253cb95595cdef5c68a8535133ca1bbf18547a1e53f029;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2de3cdcbcc2e08ef3827f3240651e6d43eac86cc597fc7d8a3ad0fd001d733dc67f523200823d7c2ca4c59faf8dfd53413adc977c8aff57b4f9382f5a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd3cc66a45225067baa40637a0ed36ede02e44b38db09fc087d5f936aa4cafaec8946a2a7cf2de15c8d0504b0ac0df7a120485c150fac3928edaec15a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92ec784973f01b89dc3905d603d7212acf3576d7e1971356a4fc88875878c81e6742b5f5585cbbd393a3aa7904a2e25c2b59fee94853074f3859e3765;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6bd85c61fc1dd6d16ec8fc077dc7b39289475a5e04f9dfc4bff6f46496fdc5d7b61b895bd23ee9440603459f700cef96d76bc1c3b6838c04ac56c3ee0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h720da66ea56ba8da1f82b46a9992082c141bf7f382b081788be37183c7182ec99a10416637db47960ded297c911f2d516af458d3daa2a5139f2ac2955;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbaacb295272e7f5161e572c45aee5f013aeb650bb8487dbad5266e6424a76ac9b6b6d9d2e721bf1046c20ef857fefe81c7fff92abad5f881a32abf983;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fe225356fc1dfc55b3011f2ac43cd09e6da26de5b8538adb95b7b6df7f1d1cee56c74b37230c26355859db3a40640c3af3b024982a462c0540751535;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7809c3df73e9f330640ca05860ec57db0ac3f0199ed8c51bc8d44b90274f47c9087f99bf519de8870ddf6d1c025e0d491a3f62ced32898391fa68f497;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c1b9b9d8661aa8cb5ffb230932dde5452cd8fe8449df5ac6be6f5aab6afdf3fc492da27233133eba295c0a9f7ac9630e12e6f3ce23aa896c29427692;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf76ecb20c3ee7a57e82d05869af328052c1e31b7947e71fabe93ab40d51187fe15a22f2a3f7c43db07986ae75eb0729c2086b84d8a24c0dc203abd00e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbce31fadfcd5b2956cfd2ee10a21d5fb8317faceaf416228bdf03417ca1d5c2dc3a83c5241c79be20e0413fbfeb0dfda5b3c3fa8c032ff34a8447be9e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h618fb4c2ff44b49f2449d12a23bcbea119df37c928fa6729f11cdc7beb6f19357a04c76c1640143de9e2a0dbafd97bf4316ba5475a0b5096f2dfc62bb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb379b83cb0e403f406233b002b3bc1ecc42cbb7a2a22d03533efbc13c6484b86ec063c84e361cd3533b1eff054cde6718b4799961cae4204de979cbb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4389e3e976a6fad63e5d2bca0c7a762c385b898ce564ac47e01a041c626667b1dcec6ded81d60ff04f6e313c0157393932c33f05b6415632c5a83e76;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he27dc726490c1c82ad81d2114c5241150df5370ad0c44b669ad1aaa29e87ea67465003f752880125314ff6270eae7498f826a039b66e631665ac6702;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6871d4151d877d6e23368affd747af99b657fb84f1ae7e960784eb2fa9a19dc41fff5505a08fe95b49689d6dfdbb264dcc19e8429dd7bc18fb301ddef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ace6366eebb0c4804f998c2add511fe5d6648dc3aa48cbcbb11adbf4589727888ccb6ba07a689d0040cc0e71ee0e51336a72de4e0cd94c456047f2b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a1345617a2b0e9df4dafc14a1d3840b66273350330784d74da8aacb3e57c84b2e047bb0eee088541ff0b954b986643afd2a9e2cd69b8e42e624b3c9d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53c68593d91c30ffbc7243616c1f85ba18432a0e6c6a5bfc867b162f485efd86e58d96889d4a8b653793f9cbf0a32054139f06198c1dbc98b354d50c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h711966af45ccd7bf96f61444d06010b9ac1493b677a78d2fd3314a494ccbb95e8cfcc972dece4a1028a643e0c261d345f1b8e559ec1feb75b01771265;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h110bfd2e42f5623499c3d38e8cb0c37e93b3c2d3cf3184b25b54eed3126c0cdd3270e629fb558ce9dd6a597af960294514798592f81445739504c11a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h168abfed2e5fdc7dcf0b92ecc994c1489b138f92a13c50245278f9cf6c427ce6a24600e181a33c9be0c5c0a5bb171024ed4159c0a5fb9cf58030af302;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9907faca11ce3e869f51ae898c59b0e6001719b221d1a6a655a5b7106e3287b45da29213f793adc34562baaf91ea5c63b33090f0149e07efbd0a891c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8af638be12700937775c6cbcd0004868ee51b4286e9460254dd56a356b29121c66a4998a620e954d2d8a53bb4e61d1d8d35576e3a5c6d55c2c76cc860;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e842ae70a5d3c8c7fce13d4a5b25dfcf6d0b6b3ecc7e258042cc8aec814299f96f44abbb4ca30d14f0b10382b4976d9006e927d93f641ec66ac4f15;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1fe5c1beb8e697c83f0f928a3875f7088f72cdbc82edb400c6e3a853bcb3ee4efad40a20a5d78de6940ba07ce2f49795e51077f350658db9652465c4e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f8aabae8294e4f5ee0e2b38cc3726772d7f3c9898dc52c2293cb858792e76ee2fe81eca628d727f8adea62d3eed4d72b0023ea84db25ac129039ad3c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd11a29240dc30e999a312e1f405992131b016325cb4968f39b0f597f139f0569a98537da2d54268a86bfea2d9d7e5e96f79fefb2bc3e719d714bfa91e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf14f7917ccf4fbfcbf7df267f6772690cdd6a613f3b0a8fbb43b452fbe685b296b9232f904e922b0f7e05912d24c84ae015fce5b9eefe1539d699d83f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h386972969abe902a8e0ac8ce0ae655d601cfe338df09f3c69fc418f21e18c101ebccd93362f93f4d957b0ec4a6527e6a8da1da160ded52fd9cfa73a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h559fc579dbf047a5e2ae0836b0bdc1cba2b9fd587bce70198ebc26ce59abdf2c40cc1e6dfae7f711adf7da6dc0a56aa700777e8acfeae8cbc02d918ab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha64a93c550281450fabcf4013cd13afb8b13e346c28700da07e94389792f54c15bbd84a2e8303065b600e6500d459cedd305ed5761a72694708d7674d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a4da278d93a6643ac946f51f28725d72fa260cf94ed6e09d4272daad29919e914f78da0ca49a9847828b9f60d0fc7a061828428d14b08bc8f3ce0c32;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9cba33292ffb557ca119681b0b2214de54e73ea905e811a7d450e7d84127cf28fc70293e16549bd27876cbeeb87affd19c96c8579d4a914db79f29dc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd39dde7e0e590168ab3f425d61c9b075fbbc397fb22009d2d2ec8390d4545aa6513a349584f02bbe1528bdcf32fb1d3e26e9a66cdd50fd837a29032ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bbf7ed8d694d031e0b0571c23e9ff55de9af2b8df2b85ed1847eb83ef253ebbd10b4c6ac51fd6b33f9e2e728e32fed8f232cc3ea0a3f1459a9b6c37f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7c877b1d85fff7364ed695c7334297ff296054b49c29963e1c20d9e0e938e268d5a9efc9eec509b6c8fc0f50ce938ad1268086eaabc35dc63ea7c789;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a1d691145287dfc1ae354ce1d28b024dab51ec8f261a753f0b604399ea1a579714a0f270d039ad5b9b46bca3132f73b6bbcc06e7d91c08e91969ffd4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20493e164fc6ee45a87935eb7550fec5fa4c25329e1bcb5df0e75fed7dd039fab8d4ad6f307a1ac89d871afba3533f0b4ebc0911e18b5c4a1001a9924;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec5975d4fdfc9cf4e110ce26fc498158ebdc8d83c98cd2c10460e6d8bbb66dfac02b9f5108126a6da037367a1675f523dff1383f0cd9992ac3948bd2a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h421df80cfa6fed98cddacbe8ce6288cec4310c7b568de800acdefad496935b17c50de2b98fa36756f9c3b10e0d89966a9d27131ffe7d8a9ce281a8e72;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fd8822859f111f24c37903d60d8d0b0259d21d1131a2e8fc88accbfc31c759070baa54ef18bcf6ed5b947e443e4393ff75a5984239c4e08807e4f53;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h679eec88b8b2b39b8b2cb3a04913d567738c02348eb362bfb084ce8cc8c25511e8e2523aac0fe7f25085484ed8aa3c7814e58b9b343135e5fb808ac9a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc378cd302056beafff581a2249d9276e622fb71336e7a0aa972cf6bc8c8f965a1b50c966631f4e1e5d353531746b666ba77bc240b7e4707f21503bab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55fa17a6106a284cd2ea18fd9a9abb34c67dfe4feb5cb7b48dbee481a66c1e3c5394e8a4669fb4b35f1016dee0105470b1cdbe7bdfc0c4713324ecd14;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb251fbd6c4c2ce3754b27e13ef3e5ace7e401a3c94ad9346a4eea790a2527fe321937aa0e36fe4254224af9470b2dad0db199613b1bbfff584c87788a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83a9eb0bf87b61c1c55aa99cc969b2fd9f124f0b24462bdc7d60bc9c7d3b0a89d2d49dac39957f54555c74e1c19a651413bca7589386ab3813e5e4f37;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66e177147f743e200dc6e85dc5765bb4cca58e3f944cbd0ec2d289e026c0e834a48b8862765ccbbed98fdb97fdc6caf47672cf33d9e0c7e4c03e9bbb3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hafba671d98ce945e44886ccaa1efb158cc7f8fa4dfdc323feb13f9991d97b22f2f9185b46d9330026bc7df67ec1f4ffbdeae459b2fbe2e60c4d3b9898;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e6f7c175458a4b7a03f2457eea2242d384c9f0818e80bc94c5e0322c7ba47df255eb48cf3f4fe41467e60ee6bd515d592b8e9c1fd42b2ebe2e3a9f14;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0fce6e1bdf0a471bdaf0ef4762967b043d6de63dc6171819bc1d42c5676b83ce64bb0d05db489bb2521843188e55cb7522ef38748d0d9b2fd58ac13a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha93dfdc1b31422f5e75342b23d0bd9a8ed66fa9f21d73eef7398d9c39cf84ea85a1a143802276b2173806d9018fd4c90b012f729af769ac45533a1215;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8be0674bb2f5ee75ba77f3b8f0d842dc7f089f9f90ec5f76f73f91e2958c34de34f6fa8106222e6041d74dd6e8e4c45ff766521105a3b329d511bd223;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4913fe22a357c5ac363284ff9929daf3cf91b43ce44f93127119be1cbaae91c6c683f434b7e4e92ff296400a47929949e0a4885c43fd140fbc0ed129;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h845da17629bc6afefff34911cd716b0a40a6c71fd5d52e1a4711d21c9a991bb6e71c58391ac8abfaa1980f3add92f25433baaf4057064c23ef95eca9a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4947b11906c66ea9c5ffae0674ee5fe5e6165ff8b635d5906ac3673b9aa73ace4e933bc91a22c4dec618f571a05f6d4ea2f6d94182205a3fa4884aedc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a3f4f5fb7602e62e62dc0da16b7f91edf2c0396e2b413c74b9bbcab8058eefa3df93bb6b346c717df3aaf513db0c864fa091e76fbc8ce646efb04124;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd018b928163e1b371f60cdb0661d6e33755975c5444d4478c3415b976bac704c56eab4c7611e8268ceadecf47d7fd3107062e2f02ec9ae06d14c92158;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80286a3c555786085e38e8cac4f5369bcb7e5ab52ad3182e1b4b086ab4cf3b64876c85f13b549b184a9947d73e612ce444ff07a79e0c16ad017e483e9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8d2278072a4e9a117eb5c52e6cd9fdc06383c1d4d2d95cb632b28d105c46a7a37eac8b5e08587cd1d4ea579224ab037f4407741344812e99b3bf08d4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9b04d1dcca0486488a555ea1ac03dad23c65c9abab82f12e27eb0b8dc39057eb091e59a3f720fb96af57ebc2385ae67882a90cc5504e6e70d4dd0fdc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b1e83381e4cc068c6228208785e1fbdce0444bc3ca37d0cb9808bbcc7c5de81cee090dee88b9f244a80c53b4e8fe52bb9533cbc148f2ef50d4aaee84;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59cda02ec95b938c39cfbd2ecb2f788a95ad30180209f45780840777358f2122b698c5e9f472b4266546415bc07f02a4c090b3573a57ba37863478200;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75aec7b08b8db7f98879196784a3db5fa6801b244a2797f22617b3d6c7de3cff6c51b0bc3945c1964bc366372cab4624589e141b3a6120762efb5faf4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28c4697c7da153164d9db01661530ca897e4a5d4569230b3b5514c2b78b3d44a3bcf0c5b66651c77a0e2a16b591f26cf6fbc6f50b527f68b556192a4d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h914f50bae9154f47023cd8d5f7352dc317f052614080f11a5f5789f278d8ad3b4d800554547f9f1e5c5af7010b9d3a3bd134d08ab1c49f60094b9d69f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2da555769f17906c3a86376c26ae96df1f2b0cc06498d119282f0cb482d8c96aa10ec1bdbd09cb475483a3c2532dc8a26cf8ea7675a75bd293ee5f2ff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea75dc18f34a1f057b5839a47c6c0669d1c4b39192a98fe00f9774847005862aa9f15224ab7df79b03077bf40c1cc650bc83ebf238620766bf8207668;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb65fc8513bfce351608fa715c5cffa4883949a6a5af6619815ea66fd3d0fc981168e4e93e49266b146ff4925ec6a494ba86fea93310b1d0af6bba6727;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fcb07b1c7bbbb744025a53cdb03c161210d4ba76868fb9e7ae5679011719a77a761f4998cc4895fed8f3c985ec7206b448dd9b1d2eaf31a9a72abaea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbb6c63b5a608d35509d1aab6eebfbe7531e3ffe4c28d9c892c929e0c381ce9ec5f8d908034889efab7026ab00cc8a008a871608521c35dc9c4f9e13c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30bfc40326ed27df2bd5764c97f83dab02e473e9b1b1727b5e57fed45ab00db2b13212986a40d122245b1bdd5dd752417bdfb44d4c2c46917f667537c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd072f068b5ab70ab18d96d0dba4c2691169f8b6dcc00c7cb825aab486311f73c428239a6af121e9b25cf62f5fd9a4dd6f98a61034251c120ebbf0c4d2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf2df70fc00d1e016bf9ae7a2777ee21a3c00a97096d2ae7f7b600ad9936037e4d62ddeaa505a419985e215c0e2070a243679d6b688dad5a571fbcc8f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ff95893bcee02de49d39b845bd4be64b8a34d2b65bef4226fc3d9589c0f2c746cac66bc80107ee2a70a980a51dbe543e47008498c8603f3617f2c30e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1939d0fbf428216e91b9dc34d84586ed734d69eb9a77500a8091b4dd41d43b5703ef399c6f3a63099f74f67d0f58bc31a84067b23823c9b984a1a01fa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2b9a516c7daa64285e32088f7008ca3e342afa4beffca0df16f4f26fc61930832c84aa04fb26730a22967c6af846cc6bfc46ca527419ca98ee9370a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f1af2f02eea180e53641d9d3334f5c31daca1510d54d8312c807a6ac319f46fa7f3eb1cb8c1129359ce122eb1acec2334365c0a2519588fc0ec60d04;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d2b2edda0000827e4716f5b1e13cb2dc3fc606b53b2aca51448ee9fe8d8c7866036184cb2fc60b11e6e39fb948ba60446dc7227b92749376b100e586;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0f7c94196c86f9059670d519e9c1502c7330708b4efe33732e3e1963cea034860d8d4a12ee86e5b17ff00b5d14ff8f4bd6668d5987279f99add695cf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9921fa379b8af322f0d4148949ece54bbb415f0f30c4167f61714475915d61f777888884373b6a1be21537a1e209174767e67e7e23db7e4aa6fc962e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4a9ab4ad01d65312dd7704f29dc67d021741f678f2520209498dfa2de5d9d7be63d92c773d87aefcb8676220a1eb9ac4f37b9907601a71a14ffdaf2a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0da91fda44f6eb57e596b2596448a2d4efb428f66ae4c72916d0f51e3dc13164c64f058f8c7b4475c07e90fc2c0c7e9de86bf58a986cb098f1b6ebc8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69490d8957962fc1edc8af47acf2b457cc322f6f570fb1df0e8cee0f3d42505bc5c3a835078d56b631cc171efa1ff23e9414c16be4add471b351331f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28c85b6bc1d344b04c7675c2820f19650ac83825666795678accb0033a3b0ef0fcf415d66ffc86f0544618e3f96999905d093335f84949fab2e5e7f0c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2676c63e6f161c753e1e2f433864d68fce81e11114f6479c26eb221f90beacb8426c06d21866451c0499df9df18d65cc94660b1171eaba1f73b1c55ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc57c6fd640e0f4d4f37169014fbdf9ffdf9aad6fac631bff028308d0e6b7ba9185501b6dd5987de2bc2fd6ec4a361224f8a96be50d39a747055c4ba38;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5daea356454a622d7f0cbd78dd4da2ae6fe7beb314a432db48bf296c4f85e15aae0edb3ba72bcc4aed390b823044e3657c70ace7fb48b8ddff01b0753;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3ed276c32a7965403be6bd3a43af55883382955ce6a93bd27132e5ebde9fc61c1d6696427f2335c203aef7cce4d269d9ae8adbd2bb53a4756d2792d3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27223ec4b46cf96dd2376fb6ec22a46e670b1e381afceffedcabb6a32c2efa3d678978b9107ce5c0ea3a1fc107cb9d829234de6ab6a6db1718bca6809;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h528e8ff884a2e6f24fc7acfb9d7a382db3295df91083a43c71ecc53e2487240fa44722605e57e3d9a666d763ae60271f84f08d627f3454095e6426eeb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc26b93848c3fd035e612584211feaca4c32c52f1e0a800a8c20201e00e72f9eda51f1dcc5565a109a85b4aeb558a7867c3d808c63aff2b7eb2e18b29e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e719cdddb94bd6f8f36db68585973066135996c45b0e98a9845dec2b7c2a620e4429ae01b804a0b21320df7c0f9a86727705996ea6ab77503c5f76dc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3cd0c072441df30ddb31f23c7d67e3cc25af542ce8c4ab1953fec24f4fdb12b17f3cf1ecb37b9be42f860c18b10030dab3274d502eb45d54f0a361efc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63eb753c38c8f7a30e1fbe832476081561afa69a4a3ca76f0779483fb29b890845fd8fb498594b990b796bab84eac45f41623cbccbfac31166e72ffd0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h395a6f231bfd097f62a79111c5bd0430ed11aca6d3437a96ff13fb379d1558af33e2b4a7307e362246a604cb58fac087c290380ddb061c96fc250c690;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31450d1790aaa844d9caf225e74c55963f215836a894dad9259cdf6fa0441cbb5abddf620d51897ba569fe427d751ca03daa9208358bc85e190afe67b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha182f2f5cbb48665f154fa002cf5a0a48b93de14695e6856653c96d087126a1ae443f34f80b2e5e500d2be46a8c0b6de162a3b3359764de795394157a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e5f158aa0ad7f04aa160eaac83290e9bc70be109016fb3b74237b92ff542f22d0e72181ab527bb9fcb0348d0a91c69235261edc6c1bf97911e225778;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h753fe3b3308e1614ec2789a2272704ec6c03b056afb25f679217aa7e1e1c88dcec24af50149405664500294955e26a51edd2f251c76287f6c7636a3ef;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h644d8a7a9f445de1c68b8b73cfbf3b8799270c312dd6a5b2fb8747a832484fa2f33dc22edb2a32e1b992f2f779a3d26c603ec1e81e72dc6111409c79;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd351d9d1f7e60e12becc90596172dfad24ec20acba0d1915e0b57022a8b34c0fc5f588e5f154ed62f98280425c0ec3d5a3509f12f03eff5347be50e19;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74ad663ee93c40ccefc22356c1e1635415736797116e349a723c38a07babb739a1f01ac4398af603309b6304209c37c60195ff7bb37538cf9e1437a63;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1596ab872b6bcaf4ee2ff1ae5bb0da5fb261d3c41e4439533c52386d5e72c176502829067bff365c3c2c9c4c33f9f69dc76eb2981033cd03c5bbb4c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9fc03c9fe40c8e9ba03170a2c356fc003b7a4aa9e7f9cfa5bcb108051b7f3f5643345ef703c941031fd289d15081383b80455ea4fa62ba623ca92a4c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc37067b54363377746108df8fdf4954f790bbe6b5498a4bf7c37b56a6a059f1fc785bd8fe696aef329b82b9429b6f7d57b7940e79454042c60faf88ce;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he37c5760fb2c4da435b7c3b67fa08f7949323ceb7625880673a8cb6497cc63b42be7295f23c09dfd7c25aa4bd7567054ce65073d299038f6b9afc94e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf02488f59727fbd5e4dcb36f81fad61a808da8807bf216406e087a1803f7b76cf7870f51bc7e45c298a19a494cc8d2567444bd0edf97c917becf7a332;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf70712892d097e260b56fe5f595fcbfa30b4f77e8ea03608f10045a3bad535dc48794688af2c84898ff6c64248e32ef3d3255c657a67be1850121ae00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb12be249fac7646d298aa68cefa8551c721855c608079996a760ec71ad7b1586d77f4ac293f23ff8b43fbfff1fd346eac5365331d0ad471dec1f7f75;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a362b30b359fa0c856ec2526e59bf990b2c06919e66bdd41d7b08108ef396727c7222a215c113427d99b834d6830cfd0c39f822b8173dd75e365d87c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51b47fccaf0800e98475db4d7a5b765adf43619e7015912fc534ef8130d71bbeeafd4883b5679a3128363c01058b701446a6d6fe4e78976f3930c6b75;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa5c964becc846ba726a2416e64ec98b13c1e8c21d69d937a257b9719daa60f82297716cc65b1009c956032ba188f77fc082221f170b10529fb2b076c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48ffa7cf1272ac311f914862d20d7b642e12f379eb7e75ccb863434c53eb7c2967fd5ce0327a5bfd441d4fef04de85b3a16935bb6c07038c7ef946689;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d9894d561600eba09f8148357f5b0d97745094afea63127ec2806c34f981c02465c376683cac2a657c0cec872be3f8cf647880a84ab667232958e309;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h183e3522a28d79cc43a578d7d2cca15505306ab93b39218ea7832fcf19fc082c6eb2b154caa15e432fad6b6501c073b4fafac3012fe4237bb47ac8d4c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae5a8bdb4856e60bbf864852ac8db2be356e1f2d4d9d1910a52a8575d93c2558756af2404d94179fc09565f14f12983c1eed11852d045033189d77f28;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab6315ac22f4bbf601e1d347a7bc32e0f3359170cbef97d0e48d94911e5209bdccc022c47d44eaf2ff2701aa9a5c757fac78273ad53c636727d79c967;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h953e1157103c1e3a976cad0fb4572557d13a55b70ac5fe273f94a746ce163c44ac3320f4999a380de33ae36f02168f402083321dfe64c20744f248bc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc07a3ce6336255bafae1e365189549b0ab087b4cbdaabad22a025d3159ce7cfc9ffa50ef14f75af212309250eb8d6d70384bbde2344bb82a5a8247ef6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7553504cc7b17ce95cb01ceae7e26ab7dd10f6e881ba149078b15ac95590124efc9b4afa0c79be9b433b7acdf037374f3b52f8d198b9caee19a18f910;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97ee40d59f7d565b00823eb3d33078c80c562bd1b31c7bb7b7f9789f37bf943ca9156f58d19c934d7b0ed6c78844caa5668f8bc568c7a787a05c45236;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbec817df3a5323e2670ed1516e58feda6f5f4a71bbf3a27adeb370075b70817af972be4c7fd99435c55b971e1ed49cd9cf259578683ab698700e757d0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c71f3f8f7c4e275c6fd7020b4cdc53c22943bd69564126fdaa8c494e764d22f36e4c5175a16383975c649d0bced86529327e89c92ba9b59fd684cfc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdd6a8e5e3daaf17bc4572108d78864e96ee48c4cba0118ef3d3edfa550dd40b8ded97d9abdd2b330f9e418e94f1020970a37131f66b56f0d4650b148;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4d6d55285fe802deb1e04891f94e164e496454d8dabc93db8cceeb44f5c5dfc15299833f761300218ecdceaaa5ffafb10270b811d3a2d0b2eaaa3940;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ec6f1e5834ec68b5531818d5163b0cb870b3578047906328806f2597be8b1589b418ac391410dc1bf627e4e34378c616c741aa97a98ff115b423d629;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46ac63b5fd6d17a45ab363453dbf9cf1498b0ea9cd1a91f62ea5c7eb95c0ab260432081ace7ca5d7fdf38ad6984bab1338060c22d59be6bfe86c0096b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6331b1c3fea0ca1e5d1efd698728a78f1ddf83ce2b81243cd2e3aed4ccabb23340ae0847c033c67ad2739c50b44a485e7ad79223da428c31ea23ef310;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e87e3f49ec64f315ab98b77ef76e27773aa118e116d948e920cdac5fa9df1f8937dca516069a7f50fa17f7450e1c1db0be9b3bdd4c23fc5463e702a9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b6c7f7ea40fd0385250d3014a0137f539bcc48746af041dae5961a9fcf0293dd6ea3aa6c04e5e6d2f5cfb17a0a598567de8f099f5111f32ed4df707;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf391381ec025ad35591938376a2c77de866ec4da6eaa3e4d7b501e6789d51c5f9a92e4aac14f60be118ff2925ba9466c49400e6e229dde8dc692bd9d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35b8b2f2e4678c863e995cf07210d83997e95df7d848e6aa01861b298f5aa5bf243ced1fe73164728c5930d0c0a3c278df50675573d14ed79762ebbcd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9a1066a1551616d301272951f430d8df403b03a2ccdbf1aebb2d8b7e8b5eb796fd30368a4c848f58c5f1373c619b7673c0ca633917b25c8b09f2e3a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa294c487d16f2058d039572022df9f17e8b0a8f7ece3ad4bc406fc641607ddfbc08b0a2311c15d1b3dc904dafa6ecafbafac9eb01465e5e8c57589b9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d51cab2cf589ad67f914e637d57b84684fca689e16ad1a3d39f74a2d6218e9cfba18dc7e866c43a0fb38cd52a714ad8c3e19ac9eb08976c87837bed3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2bbe6fc55bf80d7d85ca11dc91831ad512dfc1d302f4a229aa7fdc0a12d8ba4e799cb56e5a911cef50c360538a5953362bdec8bdaa5e6babced674f35;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb76a0a09196833b6855f6ef7a6803d4d7fb8541f9192321d2dca66634829c080e90258ed50bae1cbed3c8bfa868758a8fcf531911939052d1c9e7d54;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84e485e4ef421cd84cc6693121008c71ce9e40e0308e9fef1ffdbd2a92ff5d59366eeb3b4a9edbd8e480eefbb949b90d2096fb8c852ca730a4bd6c91a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3eb56183c7bb42a85dbba2733753ab4221f1c7b036245714c1c824a7380d65df61f47af5bf2eab747191a2edcdb4b61fb75f6bdde4967886517b011d5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h858cebdfda74b5d0498edb19be0d9d62a497a7beb9f6f00719cbc77469cd9080004a81f656c9100c2ba34d99010873a58c54da9eb7d480445dc35528b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ef03ddfe5d89cc4eacec158bb441ba5b194f2121e6da589c51b0a36b74ca1d13d47acb9c258c9087d51641c259cd2b34579f2b41c4f8cc5b7f4254e7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80604341adc7f22f59cea034e45a6048f6e2063fbc3fb82182770183613930d50c679bf152e98fdff34cd819f226dc0c4c17dac65c24e6fe33d002813;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf247f384d5efab4152795d7bdfdb86bd1f8a3c37b015799fcc955257203e7c5da62850f5b1b8baf55283fafa5d24b1c97bc5ae27f3a20eed558191c4d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74120712682ec3bdf1eb177e1648ef77504a349982a66ea6588a8b39dcc9055da45e9bbf10f320f5ac05aed11ec263d11a62055131568d235d5a7f0c1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h418ae548cd5c0949610137e79d007e5c0d2d560127b5a3af2fb5ee697621bafeffc020171fb4fcefdf9e3ca69ccc2f4db15b5a3e6452e7ea848df5fc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63ba147c32cae5d5890e169095f74d7822c3a44888fe282a676749fc683f415f4000f07c4978a8758d87b6a5faf5866edcaf9b10808a82e06ccc501ab;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb33ca40ca8d43a0f962f905c5f47fc26d41b9891c8965d9d1cf5143cf24f301e208cbe1f39a611df13279a55be8fc83f923483a56a528d0cb3ccc96;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h750dbb53efce48e1f23ca558abd912c42ab6f445733d9ca25e982ab3865fb90deeab94eee0d3489121492c2d83bc4c7e2cc020d377de79a50ec138f0b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h397a27eb62ac0a363697d56ccffa4777e45682092c2279c6946cd4c1f53a89fbc06343712440852a883a4c0e7973e035174ca4f0e0a63d16daa70bad0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b1122f649ee827788931fe5ed8d04c92f9f8407489fe7668d0d82f1db1d425b61e6233d0c8fcbb35ab83d7b85e75e3c1a3288c3563436663c74aaa7b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0cc4dc7a298cef9aa376ebd72efa0a794bd5712f8a0f947feb1bda4b890ab5845322f56c2e1d9e212df15743d120cb0b2d9fcca46c38889aa3f72c6f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1edf062ffc8a564da4a571fa8aed096450f102bf12d9a6cbd9af2c31077532df7e7d0e9e313bb3454aee99d73e0127a0c589c73cd37d287cadcb9bdb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f6671cf6871a8db7d915406c469476ca1b599dfbc29eeb50953512668ddeb38683f6f246dd5ea19702ab369c0913532e2479429f5c494a88f73043cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73591e18b5ad77468a72cd57fc46aefb7eaa3401b7c4aef0f62fc6270fbccfa952903b046a0ef0ebad2177995cacaf110f3317161084998cc7481ce18;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1bdcc6e39d02c4f8ba50090536ef885e5dd09442684851fbf48fcaa38cd8f594eef7f26c253a87281e885ed5186f0dc7bbfba016fd5ca6df045d9775a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6da44c618e7ada365ba347dbd9837b60e562e2594b13efd9f5519914450bf77be42c91d1c79b83c4f6e0753938cc5c5be276550ce0538680d6443c5ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61b2dbdf43a07885963d1c261067e58bab4595310253022930130e65be79d1bfbfbf3ff75fd33b328ab1a68cc1dfbe2a3ab7770a280adce159b37bbdf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h340dde01b0c57d6c7f099c2f04195f3594323badb337e653ae47147ef332bee60f417ecad4af70b02bd7e50d04703b2f45eacb1a21897a65f8f71b37e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19b8a15e0b9fff509459f2d35b6f8bf04774fdc6fe07d5ce65ce5e7843120b1c2e2a288b196436e0193b83445064bb7ea45b796e25a5597bae690388;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0be270b51a7199b0afae3c82792380a0c1c7ffafb5dff5716630e33f19872434ea538d73eed5747c6a84b19307a11957f3fa38ea5633c59a186df41;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcafe09bc90b8c057025d7072837bd95301ab4407a7f631251b45c31b38ebfcc66b15952c17972b1a3c905d482c891d07f7a9a9eb8b184b74f64b64f21;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdc546da14aaec17e1f8cea918ad119b4aab98b8815a6ba66e3f0b02966aaa6e163d157e9b667533a1c2c3cc8d139ac27c8e4105125728080d818da70c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebd6f3a8cb3f12c425ffd0d5275f35b38220a4ae5badd79b5e1f7b1011da3609a58d25648a09bf787e526b8f3ad5a9b80689c3355eae0c7dc748f0fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5db3da175c47a4628b54876c101a54904882d715f9a865abefdea6dcac85b6fda5180023ef0dbffe140ae92a1921f9f6396a12f9933d544dcea52556;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61ff5b95f0cd2cfbc76b6de917f40d8a5c08193586ca64ef286d7df576c26e2233846d7cbddc444712c647fd59e3cd1d548ed4932615fe52316d3abe3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4977ef9c36f8f14aa5dcf1550cd5a3e4985c71e66d1d5056669d687ae8738dcf8145b3cff20ff7d0bfeab1fa8c1c4c50536f423b4518c759bde33e0b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed5aee17c1889b6852820de65e4f1527de5df3a6ad19c5309139bacc5258983fe2bc4b9f7243e03f8d806834e8b8caf538be9e772f433ac2213af4864;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc905d7205a460e500c6b3fa148a1d1a45123c55382d73142056deb573320122be28143292c91e67eb72ff33da64627f0958a5453f82f751a8d1b458eb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba6b6202e12827c13e194a5a63d323c8da170934c3e052b56d666bd057a146dbad637bee7e34ff899ef1d63ce66bc125a52f2b20aaa63da65e1e5a3ee;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e45e24ce5199cf919f6fa7ce54722788653eac698dbb6d35e14f1da4226a44bb671a8b7dac6fd2f4443c08cd9a65de13b06d80b6c480516ebf3dcba0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7e060ccce687a8d963821246042ed923fd37eaa86fdab08cd2266b30aef488993cb38c5874e765927280f4216ddd16a7d625a4c1c7d239dd7554883;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h241beb3036351392df72e2b7d4b6de210c89c6fd4f59f4acaf15c54144d8cb3af5f44e427f34cc8b0a752e61316710fd56b123cedda6f1169a0eb8ea0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10452c28b668d802529ef2ec71d46aae9d880a91cbc7e9215e84c145d48694a71903c7cafed186985801f9b3a73d98560855158cb95bf244ac2e8a3bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19b70e070508424056a7ec348543b1539b51342c8217b1a27f979fa9528843e7553bccd7a82b008c209a7ccb400fbb25bc045c92f611176d770acda3d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b089458b4e2b169f5be99c2558d9a8abbf7602f2d48c8ff6b677315b935fd476c03f565b06ac23b43f53aa8879e00a8d87d3ca830e813c9a6368c8d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc81a650b585912a2b030d0631b6994d30213febebc14805bbfd2f6a674b7fc954197799a6a404fa7aa1c6d2f7e7b883fc9fbabe9fd8e0a9bd24036b5f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bb5e925075fe8c06f254eca79a4cc98ffe9dcf18497d712d416b8407a572932774a7e93fd071cd2c461cb0d658798c76d0dc767c7947b1df9e2d9385;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6347ad6f54660214dfd95e332f1f2c13114deb10078e5003dcec3de8dfd25e9c21fcd6858c0d5806cb27e99f42fe764b528973c30921ddd9fd0a53aa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2c6f9d9d23498e117ae8bb05803b706e3d22a105889ad129a69904770f580e0beaafcbfa70df01a074cdcabc20d05b0408a84b9b979c0f07488474;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29145239be12f58117f9e424435f4674f4014b88c55d6f27d79dd8f461317a5eb2bba727005350b8c18cbf10a7c1edcfd693425e0ae0e026aee953e1f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68dcae911083064ccb0756a37dc4de78c366fd7c3da6465429630a0f0170a4d918b05e348248e6acc1d6a9d158cb6cac1e37038684be86426d7f686fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f5c417bc07689ea34b709b5c65f853e764d413b8cd2178975dca1c29cb601e6e05f9e226980d34925ad591587367bfcefe3c1aa82fad395d9e460e0f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae8650238a5e45bcea1888c4e8acf652b861faf205737ea937de7bc464e1b478b9ab969a5c3c4900a4c64f50655763f3c19ec90c24f5debc9fde62167;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h291e453eeca251ea94aae321965a7a1e510d76ba5edc39327b004f1978964c68772c3c4d63433769326b9903720d03d000a3ef65def941f3bff86939;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb70803f1ddf639439a59f5ae12ef5bf107d309fd1c70b0b88efff528f9c6c863b1b5dbb007d7304c5190223f63d9576d44b97cbecab0c2befe56d918;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30fd80d9930a3f74adf423c3e6488661a48a72150e86232ce0dfa787cd4ac43d895e3c581f7a63b320fa1e1d075b8f1663e520e2d8a49b1a807694aa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1d4ad7cef838784d11ab6e256fa5866b5a3a17124e1cb61c6bad09ab2e94a0e6905bc34970f6c5ccab24fa6afbab4e744d9642f854c53359a4ce9239;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he42f918766e4afa07330505a2cf90fa68bd6b66506e110823afb47f594880e9d32ced85f0d71c791b124646298d2dd1e6a5a3a42fb88ae96b449cff5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5136c56ba0787f200b61c7ac723f8259e5399d8c9ebdd16a6c0916bb2e62f0caaa21e82b1a9a61bc5588a937c2e497d07ba5051bb1b71238cd05f1e5c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9974707133cb43a0e22ea48d09215b4da32488a97fa2b9801ce1ec5aeacdf70f2d147e15ad9b2edf4dec70a2aaa91ed71389f2514cad6b85764aad95c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6bc7a89d36fe9b18b4d939eaa3a952e4b54e80dc079a6d7b17ca7654147970161d3bafb922dd9373da658bd04adc62f18d9fc141a09d7d5490c2f31ae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b5a5da9be18a05acce481d07271fab5a6936eb0b4332540089b0dc8cedbb2e4db466033c17b56ea6f81a792c74b800acc7aa540f41e00ca94454e8cd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c3e0858e43d3c2768becf621ebba2806528d8142fbfa880bf00f34665cdd43d53eefb047199878eb3e3282d3a884ffc42606707fe2afc97480d76130;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88122a39f367da487b34c266989f36a2a47c7f04fe9d19b8b29dc2e5991abe4669541fccbe834a5e2bbc5828029bcc4468f45c616649e798dc0d023d7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h285c91f0048ef694b77775b4ad84e88273e8a0920b24dd48d7b56aac03a929a53233212edc97fcbc4e57cc0cdb7a46ac0f09818b9773ba99f264c2773;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h782347982759e3d2071593c3e57308cd7598681e57785c8b410a70be11832de28fba70a9a7c43dbb2326466bcb95a1c42810b642c775a6b535b9e00f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c3099cd352709d3704eac0d1896285af234abf6d2003c645dce1968154b224faa12de1d735643aeb6b512721cb9a217b3f9b37f4920d75c698df83ed;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87504aae452fe27bdb4cf928a3ee7ff7c37760e76e167a05d3718f3e428e05f03d58b856c2e256280240fc008370468d8a763fcf29621290bc636690d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88dde5bcab43ac69199ed4b0e1b0dcff351333d5150255a38d515efc3ef820baa0eac9ed506ce3a19edf8ac2b976975aae1480b9c0361be1aca314845;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3e61191f389628ffe208e61d65d222eeacddbc5d9be0098aec362582c0a1f13cef1745c0f8dc29d253998c79fcdd8eeab37e0fd95f2d11adba00521c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c5d693befc0eda9b6ccc5c7957e9c05db361cdd86200c51d9a449c1893612c8d3fe42f42521281a67bbcf34dbd2c7357749c39a451d7aa3d83d8a4e5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d6f8fdac6c13b55f213e69a691382757fd83c547fc169c25a6decce6dd15e86d8dd728fe33d27dc953fd7f43678eafb6011236e8b34f3d511aac563c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8557668d36a5027cf4971e0dd2dd9cfb69a374d5f8ad64999af56e09c4b49d0823824e3e0c85fb826e0e38dbc3547d915c990f1b057367e7a05ac329d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1aa0259123c8b96e0d7fa84a4385574bfd4c8d4911c6efa367de9d66d851e9ead813878bc8806ffb2445a9c9f0d50660859f827a28c841689731db443;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32a9fa9e9aaf9a9f1569ac31c968cb2fab4bcd29f8378230c38166064106f71042f96f460aa8be9dd0e7b7c2c8a9fe76cd272246ec2c0622f315c7fb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53a37ddc98f6f42eecb6760e4b7c6ff759f83112900cd808b14f23f25902f4d0f1cc179543901a8f5b84e3a8db8ec5cc5bd09f740625a4e2e5b5997f2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51f74c6747d5ebd2ad4a889c32a3f7ddd0370f87f60c95f6bb30aaf47d3b4847c572c9681b402b7344750f7415f491805416020abc5889a570aac2667;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf163e5cd4198495b1bae5b26e6e2c86e053c8f1be5232c8d102a8c84d01ac41ae878b84413e49dfd21852af47c67c5c36ec9147f5c64112632cf176a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99cde37247b35f59a9a4d2403c0c8aec3b9e3bfe03078c842acbd2d33d6da9641419e81ab6065a36765b2ac71db0471796bfe71898e2a025f7d2de932;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d73ed1719e74112306a11c714d3898d526bb858608bee199a9ac8e21f5f7d8df9ab2736f2e16ef43653ed923ef779f1b6393ce688eda4c52c4de0844;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa911eff9a7186c933b66d96f185c7c3ad7452839e4c524b05265aef9a51088770d4a87c2d43b7d84d57cfeb31e8aca4f5bcf45cb1c7a60fddc3f4f41;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46ab2984f2973462ec67079853db36daf69a67a63a083fdf779bdb1636830178217d64c3bcab48360abd302aed9bb198e4a6decaaa8997fda72915228;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e333922c08c4a851f8bc595e9c5f9b3d0e9108b1dce7ffd079ff7ef27612ea8c95a9e4201d62e975f34c24d232000542a4c0cd33fe99ce417d0efa2a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3af7606f6ff7544a32f3855c083d1dd888469d18ed4c33cd3358cf07c6ff0e3fc75aee060c2459d5b882e283996a359bdab2c18467653b8bacb579e7c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd36700ec0db654caa0fb34ca48e874151c35d9657fb9600960b7d5dfd95ddacdd99127af6f323d4167e011e0dddb579eeb5e0a0da428c0c6449307405;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e56ed8a10b4d5053a582de8ee90545467d1d890afa94fb20845100aecdc47b7905dfc327a88299630c88f8b81093cbdcf121e9594582bac4a6b62db1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a8488d3b4a096ce2c3ccdf50a89e6311af141515584d8086e7b40b49d8d5bf8c0b441e35920273c27f1c077a5659ef5f5e739cd0d333809a8babaa05;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a012ee8ed4c63a4b0ae593706184319dd76da8838e863b6db223a9002f1d62f3e9b6b1dd78e39487f66a8ebd79d2e27fd13fe9a1dfe8a4183a916bd2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89fa633d9f20734779bbae9a120c08b50ff75b10d53d8e814fa1f383f7fd9804578f2f5713fc2b1066e501d1f365a984bd3f6097aee5d3ad4fd5de560;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h450265d4de8556ee0cdcffb72ef01d04ee6bfbb38084a1063322da71ef9c049e8a9fe8b41454e7238a3a9fdc25efa0eca9844c0bc43e7785b9d5f3ed3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc275634c2156b9b2cfab9340df05edc85cb9f4b03d59716c5a8cee32351c997e03bbe845931606c76a3b4f8013d6b21582d6c46c011718542e2c26caf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1ff4d7dbd8dd524f78d7d453172d5eb80cc28d6a3ab1966ea9cd797e0e0654b77e9b07908625dad0bbba89d19ac39448cee61bbb4215a8e4738579a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h803a4ed752957cc5c8b69ff44fb52094246ca289dbe30a7ed6688e8ecccc23455bc92137a12e94c1df0e07521e1765383d366b2edccd1f900c32aa3f5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b5dc70cefa5671d3b3ff62e892c4222c71d7b43df6ce7168a100ccbd12cc1b9cd8fd1c6a41fa2dc894c95486357e8b8d8839d54f7663ee23476fedf1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habe59dc630d9d7884c95dea37f603533889403a67f375edb7d10d06f3d5dd6c02d84d2d0bfb7c6c599844d41adcc6eeefd9a8bff523113c9d1b05d1f1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30ecc10335be86cb1bfbbe709a585ca49e11ad7a689d7b333080209762d7294243967500988fa80129e5f21bcfea74e9dccd6710f84e3f926acef6f48;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdae0a792bcc5629803e15cc1ac61aeb3e668df87ca6e52ea2f77bf0c4b44b8d0eca5cfc0d545fd949e102602accd3ee1ea7f5f9ba7e61ce40d52c4eb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4068627908d30cc33dd543f0aa01beaca03c5d198aaada3f9202ef1f20d901cdd0a87eb85439c342ba6a66efb919f2612e35ddbdf86f2ed6b87c86cd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h492a017eb3dc04864b012c66d295a8add5a400afd541a8bab816d637c5349389fbc9f83d8f91a5d3702fddb6660c33f2be362e739fb15d222dc98918a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2e9ce7ee41ec37abea72e380333ef52dcdba6933cab5adf84a1d327ce574fba5ad7be4a81d29afac79c4ab92fc62ce56f44e300f04e2eb4de54dee5e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h929c8f204db71233ab5cd2579ae927fa261a04c3505ff91edf97fd49fa6bbe6b9d649873e75af77f04b8c58e8e6d9400e9222cd98c8dc8a2a2f652a0b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60a4456d000df173bd53040060841ccefab58a6653cd618e7089bfc49570111003165bcbba13e476cf5770c18d9f2cd1a7bfa66f73d0b4df43607d97c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hefd033138bcd5989ca2637b51fb7b0a35ec67a373644221b52b3c96c9655c2e6c1ca537e79b91c933cfe68365722f0204175111a331bec31a095b329a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78d8070016ef2a62ac72c94a50129d418bfe32358452ecd6c4af98d3c66150357e8903b4664a85e3cff40449afe76f96a0a1700456ddeee93ca634bcc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb098d20a642ae3109dadc8f4b06d2188509d9934e40298144f8871c75761ab64e1d4d254dc6cb9b78859351d356b38997b7f0df917e1867e11e561dc8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf526ba1d7853765c549f96493f3b4956255eb3569ead431e2a6098d2d9e434a0d7bf04724e22e288c81209ed6332269d9acea2322049bea807ce669d4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86832a47bddde63d7255bb143040dcb68866ba26b751b266f150f6ef8daea13e0d37cfcaf282b61a239ac287ae16cdebe6e28dfdddb2a5747644466b1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he45aa933b15dbd9569b189c222ce9609c9dbae9b87352764ea2b2fc0305204d24e2534ae2648e8380976f75336e9d8f0207dd2570d233b371f41195d5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78e77f85f847e0c1db009047d91e11e52c7db93bc1989709f238540a55b21c8e24f9a6d3e0c16a06ad75b58db023937af6e5cc6441be3a50f822309bc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hface1a94b0244b7f6f45758be5527d437cb0e8a5176d1863e348279402503dd1e909e57dd48f4880f8ad21b23e239382420ef1e38910cf0502cbff587;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h748d8a5f043391e2833e76f613ed1de5fa4a977ef0c35a96f4761c36999f0e16de1210a14971c1868490815a88c9723babc148ec38d18e07085730721;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8cbb52cfbbbb5266f50fd2b532eba439f6080fd20f74bc954a2c2b6eeacab0a1b8494a2b0bc3fd3c58dd79a430056a15ca7bf31ef4b9001f069646f12;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1c93f83a29b3eb0160e35532f6a80193ef3acdd33e3503d9ceb26aa928394321a1ce7d8828d6bb41e8bffdb0d20d9ef92d657de118c8edd67f4d3b0f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbb63e36880b146ec5ff8897a0c2b9d7a009ec993235268fd25e886fbcdf009efa8833e8c9cf42c82bdbdd92b8ea9a26e8c95540a07ccf0ba72b24379;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4b2a56536f174bc1464b8beb1e28564522c1b191f46f9ad8070841095abd518a12faf51a7969c989b4ad4044b651132e70c53bff247963843fafb0cc6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6677abce91e8475ccd9103cf13ba0e61a86859d9b7c90cae049d828414c364511beb54e8e4072552239572171d14885748ba655816dccd9542440cae6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4eb06e8f2dc8d075c000c4156f4d516a5f60bec7df0e5a0eeafbe3dc0c3ff71a8c0a973c0cd3ade50b5b7818f02ab42d75b150336958bb32a5bdbb60;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6f870a5df058e3577d522b3e5fced2bab8a0f4ad1d918937ed84db705ceeaa7aff9e7ca9baef22e0e4131e09a8b51f50040846937b12cdcf448b2e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h244e040e560392b69cf1cbbe122e2d857dbc5b33d48dbaec295c6e390fd5f7e15e13dbd0a494476b614c9f4b29517257aa1e67e025306ad79ac59c8fa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5822aee2f21dcb355df02a22193533eb23c9bfd4c72387b62256374857c107974d70be9eb930f96565092adce47b8d7ee0b1c20a491cd46cc06f5201c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he83bc5f0688797b7d3a9c5803131d5320dc9a40ca163603fd5277bb9c52fccfc9b5298e862f92fe767b9c40d841962d7c83e576fbc4b53e78a1e0368f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff66045eabaab25aa78893ca080a7459da4964f2d627f1931409855447c9d0e03be62f21b8650eb08d86c375c5e91af2d537bb8f75dab6751ed0958c6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b0f0dce4d581fb8c61fae2202fecf1ce37f17dc538494f97d77da91d8b3417bc1ca66c0f6bdd48fff279776c13e55114bc1d60e7443a7e47241b007;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d806a52f21aef29d8f29856c0491720678e7c626ce5877742b87f2a634fc7ceafa472698dc21d196767dcd0e7d54064784bd79efe1911dbcdbe79116;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h81796f121fc90bfc3216e46595620bb652670016ad19007a48051a2a92bf3b34c35f11052d08bb85e8b3d32a0a104f5eeca248fc29a64cdea5238805a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hafabfb0b4a5983860e3e52993a6292990a4daaaeceadd6141423df730d07069f3bd820da6eb5cb174b317113b9e019aa10d7077e311ea508ef677dde8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f4b1e8e0c019b19424dcb678f4e0b16ef3f8ee4cbaea015fad2a03e6e8bf6e998be6c40aec1c760b4c8d7d70c9da98b76e1a518ca93cc809a7b4c6cf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbc17d904f03107199e88b1b4a8ee15c66aa731846fca199179179af96c91604925b4c90fc22208dcd001b6d3cb97cdfd629f8150ba88a1784a22b7a4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e5c563d0c588e1b976f69ad4188408cdbe2c95716bf39e1f5c6030f83bd1db0ff3496f69ddfa232592076c2a7fc0dc1ccc17ed38275bca6283c62aa0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd07ee9b2088db60811bfa318d6097fc29eb3b038563cf512f1440d8a55089e7ce88d7b405febaa45221d29d1a202c6ca3c86961c6e602093cfb3027d8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76ec9556021ef9dfc49c35be1a348ee949f32fff366df153e11ce39942bea559f657342ed0a5daa2687565d8b778e339012be71d1b8376bc4fea9ef51;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he14d2d850ceea30396031ada3d1fe8709f60132d11d31face68cda8a250e8b18b931ff44e78709304d4e330c81aaf1b4fd1fdfcf83f9f9a8994441d69;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9999c7b963d20c13f287a23f04c4f7039efd49260b1e5a6d9080348fc038c94e6fc9238a531f16ac237e51691d8c3e958c7381f96d5902843b0b2d0d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2b5525a786a40bd9c88cde802e30806cf6b2376dea9ce826628271991b28032c221e72401cceaa79f830fbb39e9c300d1756446bc4bdad373b1c382;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4c0d6478552aca03052562fcc4c51a8426e49e9d3276c11b9a26518728f0c29dc16e501771ada008f3a59b30ff424193d8e5842675c7d6566ff124d2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6311842c474c7426d758f342fec8f9a0c5406765c824d1f5cc0d0daa8dc680f78ac127852103877e97d8d775d302d365948f82bbd385450dcecbb1eb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8eada0b74244ca5d962584d94e59172d25b5ac38ed6611fad2d03e40b0545a7a95921c913903839f46a56ab0c163800a63da12aa946e2850b8123293a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15e7816a5d62a4fdfd2382e517458ad609a88d6ea0a1d5792f77146e3a769e9f0e232b725cb221e69207814a295d85294e3d98dd8e488a0c4b3850d3b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h14116ddc74f5f3947a21de84f2e4705e474537e2128c361334ac9a6352c556de044ecad17aac592f3d91c37d360d2dfc598a4524865e2b2e983d74cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27116ebb57dbab54c9a41aae8d56d9b42100fc6fd4aae23c3c13c1ce0aeb9cb84c5e12ade7b757349941bb720f5450b134116022853f08cead3ec3302;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1b19ef983434041535dc3c4d2ff50cc142db89e65dd0c5512a4751e57b6efe7e2f5397f5cb1ca361f0e6c621e9e68af32078b06f5327a7e5e8a7f188;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4043c6bb6f94a1c28615ca4c0f1060a516d051dde51953368721f09288897de15e80fa50bba7659261da1b6b665aafd01c0e3327ffb699eb04cb24b33;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc066feb1d530f4a04fb2633e36fa57142c47a2371470c7099924f624d4c897ba51da1d810e44dddce0441c6aff043aa73e1fbca7ecdb5a210f7ee5794;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae2bbfb8e926ad4c55a0d036dd623612d9d71166721319b63f4660b49a358f989820cef8277f7d1de3b4a94b2e53821d54e2cc21ee4ae94891d279826;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc45725cdbdd97000f8e2ebb966a446ce21bf165093c3b9596c4ea1a41fc1403bee7f72158433152672cc9a801aaf7d031790ccdd8497aa5bdd197cf81;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2a228001ef3855983e64185b169d575328d2298d268553931e774d28a2938ae855d46d613e3d7f69c9d14b0d2458a9802e1fa63772d1ed3a35c968d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc0529394a9ab92aac082fc6dc19a15ab0953920157b588dd3f1d1719565874b9ab89d55411ec1b65ae9331b8a3f819c38d09fc2f8b4d9a6e69da858e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a157eff120cf746d480e03511c7c6681848e608740d2ae2d98cd7f03d9cac0ea30f90a57528645d8fc17d1aceeac269f84700202df74ada83aa54c70;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb6c89bf37f4e03b5d203ad101b660e8cfd51156d83610376cb70eff056c0e81872004e15ac51a1a5d3bc79f1c5aa8eaca10abc4078776d60c97242d5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdff2ff5a3298d9ee9123db5ff7adaa55cea7a83a80be5cea48ed732c7784dfc2731ecaa5cb5e50be070ccd31be0284243349d5934de682845f99caadf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0c309039d15f2dde2d62feb338bee59329acc13dd143a039f63170c31d603c8eaaaa5f724bfe0020bd3b2edaa59969c48d3f871ae825d1557bfb9dd5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d9ac2292cc873f86caf7e33ad31ca01f90b8d3c9d5b9c7eb4054a4b299607ef9a9880e8a5e57d0f714b612316cc29c3866e3ca44669ec2e8ab4d85c8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f3fbdceda8a9f3d39e45379c140564e21d6be039a692fccf51d7c60b09dc10a0f2ded7caa410b513e349247e346be811cf6144c1e6d4f7d73bc71b8b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40e9565ddc8287bda657dfd0d840bdc1ad5421274801a3985208625e50468d367ceaf480aba8189e51e4b9295e3bd873e4e674c6f8aa677abf652b1a1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93086025dfece80e64bb640b3a062c801eb68204ef55eea03690d7ca6134abeeab7e89824265b7e3f295ad01e7b674da4fe2b19bb22976fa81a9a719a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9db002971bfd1a156507a62e8d084fefa098d3eb9e8de51e7a402808d0b7f1712b863a1462f9039d776f86076053de19a000d656d07b4196a50b2c35f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h565a45f508b35430b523713e63c8d98fd1646c5308226766a58a89aad3d43940a8113dd647a5d0d660041ec0d415f6dbebcb60e5de10c9c59dec426ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72bc9771049bc2ad41404275b085af2e574e4bd46b70f4a3eeafe44397e2abc8a4b2f98a694d7853aafffde4788ca7382253f0eea2e74aa41ffb3fa00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h440d2df09caab07278b2a3efdc75b278ea484a9d34315c93dab12323bcd669e377a9b3b2bbfd4fd3753a72aec07ce9f7821efd5f5a7afa0acb3707360;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he11369723dd827b1a712cff625b180d5a4215741a4ece25c6e26595d0d1ff35117b9d873eceb9803e2debbf4ddd7a74fdcb56b7bbf393959785ee924e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h583c6859109a36d8d886af9b874f14942d4423309d4783d5f99f64b5f60c58889453f243180eeb25c98bb8f3462e14e9281a8f2f082807be13c1c714b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc61f019ab2a5e5b7b7e02b4f9730895380dfab8a01d11684ba5ce7b082ca429f6dd9adbf46d5187543bf166c62f0cfeac25c1bf9755042585d66fceb9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26b415b2befb7312a0d8516de8f158e3431c52898d0fabbcea0fdba06bc2238696eab5294fb8a662c1a9053b8926feaef54ec229dd46a431b010b3799;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd86aa5ccdbe534f875b46313f46c7a4d8e6e098428b88ea5429482948dac5615b91755148c014dde353271cbe4ceb78bb177b28ba13f189ba0eb673af;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a474f495193fc4ac67b69451b081ea90ab0ef9b4bfbb23e7f3a0bb9685c6e5327ae7c21639e6326e21a88670709d51c7f5327e73c568a4019b8a008a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdc356a189c66c3c099db5726e2319babe3125b7d7762b0dc1afdde345816e056b14487f8361e2a380b18a2456c649ce6b42aaaa18b40176943781af8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4b9522387e1958489767ada124c39e5bc079c4219d622c5bacdce6187c716bd194b545744186e3d4ca2f876f0454c3b268b854ba550363b9192d26a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had1eacf3e4369f838569ea30acdb1274333d3f249f93e3da30e83d8e1b0a776f9db8cc3f4eb03364ba58af25ba963c32e42fdeff1fc2c042409ed1cbe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h566be999e5f7d34956a4508a722ea5907de1f00fda5bec58fc83f22cf6268d7d2a8b963026ab416114b70bfef2492527b05afe48e7108fdcf35faedb6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2279a6bc7dacafbae4f902a406c915a44559fee14543abd9b922e2881d2d43f11b697180568b9795bd0366fc6bceb3e6bfbe33a768cd8ec47dafe5ed5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6fbe0774edc3167fff346a5a1d1653c5f127ba724e2a55f557071d60ebe4920cf88dc5a3c71f150f3207dcd567a6796610b3d8b40fc48859ad270e48;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h652f40dc5eb0bfb0d64243027007ae2e7c7cea7c63db0e15d90f11698d97d77ce1b8958688b808e63ee1a14e9df79350a74d6b100fefe5e587fac6bc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd746c396dfdcdc3f3397364d8009319a71102a1a71297fbb67b0486e097bf48d6559184e1dcfda7461cef59a22f468ddaa913bc1620462df3b9c95fc4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd87b0bc5bf94afb4d78dbee8f85fc9739c4089dcbdbf96613a7d493366d536753882139f16b711e76d97784eea4fde02ea03a5ff0c682b024ec9264;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd69978315060e25c122992192807135714c0e6dbb02be247c178ee7e1987340a575275796e98323f3239a18acde8941b67d5332b812c8ab68998aaa22;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a72d601e15353a38defce7753b1ba7603ccd1796bc9c795ee252885abb657464b3b01eb95e9f3e6777fa1daa875667f9e4637688f71d6676d2f973e6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab77eebb3d5a35a7152d185d26386a2be204787211543cc4cb3ec936b265a237f12b4627b2d611df5bd1a03baa6144963658fe700fb8870c3af6248b7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e63e9e158e48a939bfe8ea16a54326660d416dfc3d5aa1afc5fd38754e98cbb09fbc1899d7ff4fce7c02d589e0976d99383d03cf5667cecbfbf32340;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haed905c88e71b00c894e568ecc854ff6e4e396e7964cc59d571ba0950456ef1e483d10b6a43e9b2a86ededd3173bd7e34cc6b809d3488167be1bb398b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3af7920bd66a3244031093f0328f962c7c09a68bc74787aab478ff013c302e05be89fd731b9028ca2061d20c82939d39c85de23df874774e05bfa98b9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha331f787b2804f4dba9305f694839d9f01ba9582eaf929c1d9f40e804bdb92ad91ebe75145e5868b3f7425c0a482c26d6c369061e1900d0652f9c388f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2cc9cf0d3fad44eeb83f4c60a6644e309abe50ade525ab915ff2a53d413c83702fd5c20d0fef78489b990777cff2cbdd2615593728c0ed2aeaec2a332;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd782b95a8607a20132522700b879708c2a8c668c014647743582236dcb386d09ee7106a6eb9e8feae6141d24cda95699fdba6945d7aaf6d0436be1a58;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98d8d39a566d8cad95ea4f2b5f2b4b5821a933103eb8d752a1c853963afdec726002edc8793cb76f692ff211149350594344317d67d18a598cbd68c93;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5376cd48e81061f23f09d4a9e1acaa789f3b4e1c11d81e882c3623f87130f4596de1647169ab6c4b25ca140e4153865db2c15f2d967d67378151bc1f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h637b4d64c446c66a1ac198fa8a74cbfa37fff60fa98f9a9fb0551c1d000504f6d1b024add96548bb9c82620d2ddd17685cc7be5768a21fe08c4c49900;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha44e8e95508f8b02471e387257f4c1afb81904e2df212b440b4e373e6fe3b27e969deea6521fa5b2bde86df6fcea2140dbd767c7561000c48df79c2e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb2593042ab25118d39b8627bc33cfb50a312a7720de4d4d9d0563ac5970205af561b4743c3688638a284601115472691ae80c794fd712ce3315eee44;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ba18501bb8ace00bae2ad5402e34e4c8f0e88b07be6b3fbcc9bfdd3248e46562ae381d1dca2e68bc24a79ff94d71dc5a9087e5312e12b26bb890461c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ada307136f1a7de7a58515e07478aa19d48411caeb2a8c14c2625e4b25be6e7a57776c5162578292b0ef79166319da2b824b95a23faa22c5d893796b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ef488f7e357a3dde6326d13902da576c76939021939555a39c3b163e60801d6a51a895f93e7ea9956b02e85331da86e5eef65c8cf6328920e2983bbf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b9aca0960cd7b01549a3039f93bb4d103804ff5c93a950d0d80edb6b98725f30f10a70976e00e19fa03f9edb9c9010638e97ea2d91e0e117550bac5c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51d592df099b11553c66f5a55d0f7c715aed4178b87ab5605ad81b7db22e26c12fc8691103ba703d45752c3d62e279026da90947af7438658bdaa0fcc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe48cebd3b3966974e213833d1b7d2afd5d5b74c7459c26b957fa1e1af37822a7a54b60c64a1b7b75a1799151a3fbe0b86ee371acd60fcf1758fa14ae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb41ad110775de8ea996e6d7657a89a91aa8b2e024767dae1ef2fba4bcd657caa203fc6fe777d525c637ef50f4a57f81047eeb6d94cc0ab21ac0362454;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e4d4299af3bc8a4ff51aca05b6c03f1af5d04293483c7f0825ced74c8eb9debd52ac787894f2fdf62f11765b3a7c1e054cb44d2c4964501536bf8406;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93951584005aaa2ebe27a473f9dc448605131bfd2847ab95dd4a021e68a4ab38facda184f0f90843cb84c857bd90454241e592ff46e8ac2e6defe259a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h931e417784bbfd9ca1f234cc34b1d552e0e5276b9ea5f5f33e01f771c3c18224f9259777ea590f2701cdd467cd7183595fa2029926b12ac3a17ecc986;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b8c54471aa80334a672bbc9ea0ad57f339280ff4e9c1e6d89bc919dd0b3c11913d39e115b79b2c2ab5835831ce0368c7f871b516489d74224753e85f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1369e965328286a763ebf283c3db1aaa8774b0edabf0e0ad5fcdb29c44b4f0629843d5c410ffa4ec9f2cbb021a200e811c917a2d98ca8dd89f0053c7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3a93aab5d18dabdb32de69053cdf1620817660258c0615ba1ccdea2ee351ca795db4be44e5d7074adec07a4e8c982ba9f39d4f352e4609d6a4434ada9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h704e8d9f43c17683238d75ec052d807548752d3a519144b1170fab90adcc5ba01a6261f68d82c38a425d0a1174134636bc97314a4e81ada1364912539;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7e8d2c0455a47af464c7dc729e1a0be3b16aca421d6fc35b406112046d818810bccc88ca5fc524d92f710e28d63fc45ca7ea45b30104b5132cf5d14e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6be95146115c23d9c914e61580e5d77e66ee5fbe4626d131614779874e8f31afb0fa90567b00271829823dd2eb65c7f125a3b40e3ec9672122bdf508e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1f2e3c7b2ae6358f4572e841776c8ffc0fc7d7a4f40cae6e2c6030742ec5f5f6c0be8e8f13b843d9d0dbff5491415f6432a369bebc88b6b0b15134c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c5eae0a909eb8e215fb95c8796d373abc1bd5f13a5a6c4b5b065bf7ae9dd3eff5eaaf0f262eea321f0084c6697d5045c602d7e51570e9790519679f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3cd90b8eec212e9725d8f88e78c37bb884febe6df90448ec3ccc9b6b9c673447dbaa727ce6e64c1c0ff98f3307d54c798775890a3333cc33e9c72e9f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h370ec191c2596a5aa975b3a5cdade74b5c449c1fea3c248b531ea313b667146191aeb4aa2c2cc87259d202ee1f5d31bdcbb356ebed39512bdac49d560;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e23628b08ac1d1a267ebaf59952313361e699c78e95905ac2938dd1719198a8419383a3a392db5624f86a628c02477233b2eaae6fc836f9d85684949;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h82e951c5fd37feca16f0e74fbec7f65fd7a77c7fc637a73545612759eec0a344623cc145686a217e0ea478c4bcf6c965d83cde874eb760e2d7cdac56f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99af3ef51e3438298466fb0e67b891468ecd315119dca6c3ecda778840269af1e1b51fe53505c042a67ef307c2629cbac8d99d3e8378f42d47bbace04;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7340a2f7661cebb3058bd8a1ffd11f7acbd07a24ed6160b1b39190a20a235132a26bd5ed01751f5ba418b1801472a7d485ac94d18e2b7b0a49c40da64;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdeb8f074101b8c7f5b6b1d7a55aff80b0d68c3858eef74024b2467072924989edcaa0176d9b3ed11954e7bceb0ca92ba45c1112c6cb85104f955212c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e509c5439d9f9333095575ac80ecbb22549dfb0fdd862b722124673fc45cdb59290dbd48b97af18f74d8679d1827c7e41c79a02096177fc7b01ad90a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b3ee723c7765decc500ac45a28beecc0accd65fe35d1f6ce87f3d08452e0b1d1289fd5cc830f423ef726284f8a20dabecec62712068557ab0c878ec7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf75fda98957a504798a2a37ffadc216407a691ffb5817a7ebc810fce90599152e593ed942ef1950b7c15b56d14ed196243cf3a00b203a55705c55d212;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25f6167f247983cab004934ce0cef6a8c8b145d91b45783c8a1022ced1408d9a57d2824ab7c4be40b986c4d8caf266b3ddaa20823c6e36b27f9481130;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48ffb38ad9a3c7af4707b1c896750beb42201958d39d3ecc6d65e7cd272eda8576a3f3df6cba889a648d559ff5ca991a1cd579aae6f17d91f58f9deae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1abaf77cd34f4a4c78108008f41ffbb2dbfed189be741828c064846fe36fbc8a911f38c6381a0c829135135932ad7605382727e305b60fa00a4ca7fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdfd4259843cafa5877eead96ae629fd27a904c401cc52737f557b66dd051197239b1a0074a01635251c7c63ef1363be639c9bff6490628dd45e7ffcc3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96d82bd888029d4315a40922297ba4fa0574b88634deea76f2a8f384b6dd2585f98f2a7bf8ca546823481bfb200c53ddff17efbd50a6f968d8929139d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d76bb4f75fe7982505ffd2395b284e868a6b44472f525581cfbe271889c62cc2c8f9afdaaf770d251a4bef0c0c7287506087da92d1bf2734cb4183e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13c43477cbe13d3e769b2dba6253dcdb880338e6344822d2ef1aac0539faf49357b7e1a51b1a15a55d38a1f73c1231db5e7f57ccd843cf24910fc6643;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h397741f16221391af4bc953da4108a88fdb58f533b16398f7993dc826b91377f25c7e59f53ecd200eb59f46bab72ba3522e910db2ac41523a14d6718e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1e853aad1b8bdec16a8e4ae138c08efc0c9f6ec7eca0612669e174f52906e6425f19555c0279c3a1010227373a74b52ef2f8affb704d5b238fb157a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8cb83f8279058665eeb73da8a03bdb23f4bd09abec1d559e35b4d77aa1b1e59de9d16bcf505b810cdfc9af2da93a9bf339941bda22fddaeae70aa4f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6003e718baa9841280f63945e7b73c6e3a134b92f8149f2d8506e07a1a9180ba6ce9325aab0b3e2b81c49e69a57fef606b533a63b98030b27ace27a09;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31f11d97d5b6cf311c2f130cf6e83581a8d472b348b6ed311ff2cc40e764563328c3e36dc099d1d74b11fb6e25899e692a9071d0d6c870210de219c6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57ec4b30ce8b8949079fb68fe21551b8cec1c5a11ba00783d6530ce2066c2aab2f5544ce05f1f41a40ffd90eccc8fbb39a7bb58545dda4f06caf22a9b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1bf1d79f4711f462c9e42eb13c8dc5f9c65bb964d7dbba0a15e2594401553b5124061238b47dbd1d6b9d9a32707cb13660d2abdb3ed4bdae298dffbf1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2777539c6a63e2a6a481609c8900315cc24f559ab01f93b604d373bbf704af5207899aacceaafee42365cb2ff5dcfe6776f01c835bd99f94ee5ad2593;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc60cb42efd1e42fe5f838f1bb7046c104624864c3e3c6a35f4f98ba20d513521c18c98d0924c14dd968f37f9a8209d9402ec1b7d1c15c9415193c1069;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h644afae753a47ef7aa25e56b410ea0db73e9551cdd7c0a2cd6b3cdb8a572ecdb380d395dbb29b03816515405e588529f8b547375e4291fa700e917002;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff9ac8f256fd55fe5e14441856a7c336a56018b584a020efa1f56717a31a34cd185007a0bd2e06b3c5fea27fb4aabe64a2ed0a7e8ad3c07e4dfe9d19b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha65d3c4b5e7e75db6f2239b543e7445547cdc60336cde1ad1ff1f3d714d968741cf165f25529443e180e3efea3ae1f267141f87c10912b90c191ec546;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef40df5631a6cc6c01ea1778561e1c508534dcfce8f307e70f4cda4a4903b2e9bca64be1b0589fa24707e1819db39d7840c7ebb9329a59bdc02b0f890;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b97aa6f12ea0469eea587ed6e777be739dd54a8e0667dfeadb32bd7674ce0e8b77e876968ea768a6a6b2a833696d0250f9b11f99f294a5731266fe61;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6125046bef1b6c3b4eea82ae813d37684565872c401884b809ec07a3215ed77508aab7962e3b45b8db62e8ba8eeb166827f0536bc24cbf6b87b02e3b3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h619fd743be8f4194febf1b83003fe0c310ee6c24144f08f75956b85a4f8bef8f996a1aa09ce4c78d237329eb76ade995dec43e2b9d68b48f5ca1ef59e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb9976c349e0895fbc70a4d2b16fd086c5580a03f29636c1010696eb2fb42865d0c3067ce79ab88ca8073d7af41052d24cc2022e721f572556a6cdb8c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a9cbcb41daf66fc07506ac5de112bcfb48a6112353d5022a5e4974eb31c16a8cb4b8a2111d7f6e8a3e3dc6937b974e7be0df9e16e16d194a3e677d01;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hafdcea8c272ac84f2470503ed27a227efdb0887996c5c13efa35c3b6229d591de58331ba2a166d3892f80bbf6cfbc03c32bc7ce38b229460f003e4f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56876ebb97e17480147d89c49358ed6f897bb65033c0faab11a2a2afb37b83c7168f8920fb6cfea37c0a8c6c329479bbd469480ff4aa5caa9b66119a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89a3f970c588ee0beb359ff0f4678ed98d1f17fd9108df32a096ec9e8720f99c88e179626d7f2a417866bd3d74385e99c59af16e22f0841c2ddf9d7bb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c7290de5fa55d9c107f085b46a7202855b25ecf8d5082453af9f5eaf0c9030229364bbe383d634d22deb70e259007f4873ffd8e84d65279ab78e9ff3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84d520d39a790e01cc0369d1aa0e9c29a6de4a49df9e53af131b034269ac3ea6a5c120a2f480a7903f6141006252137ca4bc2e3eac3e5d742d11b322b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c1f6724dda805c577473f2aba0a348775bf5fcb92189be51cc5356aa2b9263b391d7b800f647de50d08a1136baede62fa397a9c0687f143b10d2bd17;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h528b9122deac98fd4c41b09957c61599bd4836a410be66247f7e233e39a3a6dc0d501e6cf263b072b45f0166248d54104aab3cc67808b7a9329da6c12;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37ee6edd1dfda80f68f2c1221af6a04fea6e5330aa9a8832055a8d135b0e9c64cc541012b1416593ab659796add5eb6d7cf2a15b21f184e199dcd8fa4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h935325a553262515f4fb9aeb74841374fe3f0238228f1fd7e14b3ad7466e226c041f93f209d79aae4bf0af8f3aa2ad2056055d7b4ab1b91182f3e64a8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h430fd0bb22f3e735cc29b5e4d153f70dd0bef5bf05bfc925a8d80aec1a6085926a3f624779beb27f62e4c225db24c57302f75b87219479d56d4fc2ffe;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha031cd2df342052c2e9570628d955227b15faf088854212f29965fb08cd97f9cb5bacfd9dba3307ecee3f1e3efabc70bdbc0970364e9f88d679593395;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2fce467307c962937b82b9073300b7fdc0b7c2b58ae874f470282c3ec8cae64c7936eec17eaabf7ac3b336751239450f22837ad905b8e6b503e725b3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f49dfd931347dc64748d6f6e20f053a49d1f8e7401a3e158137fd62e95af07fc67b56c6a46f73411a4fe1c1e267af777d4f6655595a7f2abc76e5e36;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ef3b2cc77b532cd3ada388c7b87dc258b924a389b1e75ea07cc6d155272b57f04d07be8dbfaa53c3a633eb383e5fb63a22b02929d574f51a1f2f0a13;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha54c1a3f0087e7fb25d14f3bb5e79505222651521aaa6828c186b59796aa8fe51a107197fb84970f6526a4d771ed9aa010356dde33366b1c14c92f1c5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c825fe31bacf5c71ebd2b07501843c2f2b153b0af52c70a620a151aebfc204f8908712278630cab6e5c2c5a670c73eeb7ec0b217f6469e8833bcbf17;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e41b110b4b4756e5ba6e526eecbc14c93b29dc5b871506a13031fd25ccea9b03982549b7645bf60b3729d76e30ad27b8babee1e939b7a32723f020;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5cb04fa0f380176d2509cea18ece2ce2255946be636376e57c02a9d7d3909841d78fd9eddc3d36a58b97ee1b3e77254a8850d516a62f57006295bb64;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e9369d25838db16de15f53c16de96d68305020c767b8bb1cac0e49d6537043f1a172852b039f35c90067e7a271217d23296b11095e5e8636ae5602e0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4259d8d3bebd9f279c60d1315768639497235aa2af651944bd8863a15b598bee3af6cf0da97cbb8f093c5d7897943ffc42482a9600f3198054f167aa;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf35565536d8384504ddfd31039a3d7d46e44f4bf3e29d038b4bfede2fe3546d23e18e9a6cb97aa025490bdf540b168e8d2f3f68cdfd594d6967a68ecb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a2e41da189df4bdf126a8b71b8f9c577654c7f213223d6e15278bb6257c834f922fa0b0247419e4b0cbded5cbbcb365ad5b88c89721f50a601e75e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25648649466c8e7355160a481d28f588b9941cab20d79c1db048bfd82f66fbd9a77e9b7e90d85b802e8e1d2e0f1655df02524a441690d776470c26865;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54f238e57308b6a732307e860a8c2263e3eb39a820c4bb8bbbda2fc4afdc91572b8fcc9d0b0e26b681d3f973f93aad5fc4d7c910b3daeaccb0feee7e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6805f32c20d79dabfae5c60320f66ff7776e88c2be25ce50366076f4de7e994cd8bddc02ed38aa8697664b1021951d3257531fe5f04aec244bf932a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h935397d4f95382a97a3e36047353457151129929955ddf0d92dccae07372b43fb880b24e516467f522ed639a172902aacd878754b1ca0e78828d5d845;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ec3cefb1e1d28e22457acc8fe9ecf242040db141aecdd6fb0b0849843607ff5ff4de1fe03dd0d6084c2bfdbfbfe8d41eaad34f5fedbddb7e1332c63a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c6ff3e1c4b6a3d5c36f1d1b48eb80b8575d27eb11c0d668267bce4010b27f4f87a39027368f7cedc0de52cb01767f93628b2dfb0b526f71b9fa2ee7a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h22cb614a6192ad4ae57035f45755dbca9d9d584b3ad451dd4b5680959af3f311d96b9f41db79813a20c73a8c9570c7be72991db12b8ef8617620b0023;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab4e139f914f5b25c3436699658807c621e536b30891eae85afd805a244057b70acb7d77de5d55d961961e56cfc94d0681cce59b4bc1375df79232851;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ba8f787a5d95d4d712801b2d70c1c7bef6040e538d1ae00e5f826f5d3deb5a75e6de50bb056ca86bc4a38d25999d15ccba19a3ad66e87edc712c1f5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h212d28d0216fd8b7fcee1370c7914e61eedeae9ce2c72b5a2ee23fdd3846a337f65a2bbeb40dba860556a0e2c0532a1ecdfcbd4d87471114cff53e462;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d03118283c42e60ce11f9c8bd9834c645b2d287b636321f841d3d9e1d8c42492659e9694600e2c2c21bd12b77c68e181ff489fab22b65fcbca46c90e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa4390b2d59f517ec09bc0d31a37d25a87c00541d8c69d2c86c55aad07ec38998a6d9c1f74b9dcdbe0886d3c84c1f209c98c6bd4b9638c4656f105e8e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdecd796ec851432497d3ed8f4204f853f9ad91c3e802d03f8e009818b528c88f4cbfdc5241f6a417e88ad80cfd4b698d9de5722f4c20479721c1fa3f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h427a7ac2bdb0968b268e71fb670bd8e2de55005aeea4b9c3121897dcddb68eb0ccdebb768e0b28e3ce1f99a66638de3a987560463d0502a54ba60e1fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h431d2b489fd502c05dbfcde45c112482564a5d10fe423d5e6dbb5eaf2e21c6f7263833d85b3da23fc14780211f2bf4b5ae3bf15daaef632457d89691;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4963bb7b8d48a779725ca9cc2c5403ba2dfe1d96de3c25477db28811afd45b28e16259cba8113ec68dd0906dff19aef76d63f32adab79058320d2ed4e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h828b0a1f69d4d3df1a62c12c6f20ea3011b5757cc097b39e55590b7c2259cea41efdbf9c87ae51304fb515f0c7f73070567efbc61634d58704b2ccc7d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8f4b77dd702c98abda24ada789ae31ac196ba7b94b6df65f404c4a182736e2a0b2fea73c0c46fd57afec1e9a83ff56d1322a9c60d37d5467609269a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ab13555c5d2d6e4d9fb04c37f26a581166b7b752964e68dea224d0cd3928ce41643b9acda6827a364f971c08804cdc3e24e416687bcef74cd47c1c09;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76f43e41154a5f99876b978941f642ea1fdae3c53ede7306f6471ba6be8c42032261142ea1055f686ec704f3e4cfe4c15404be565e887769c8a6d39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6be6292522574658eb4ecd5d4fdad506b1d0a182ec52ffab18313b78e8fde9bc3a66a485c2fd59f7fe3fec6027cc9a39ae3969bbac6b0c0390109168a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc77c2f6504cf75ea5b49ff6e8f8de57861b638cdb9965fb526078ae619ed0527b8fb44c73937ad76cf29c7fc016c658bf630bfcb4b7200815cd70582;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h572925b26bb69b8816aa35ffe498ff3a6054bf9b5d19801ba66a3c3a8485371d45db58ffcf4692c7e11e4fe7e8e6441ac2ad2092dbb8490004dc819f9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5432b7cc0be7df69510fdfd5a99cde6a7753b67cd077ae25e50999988b05df7e227b858f0f2892009cec0d18b9ab3fcfc4fe6ff7e6089fdb617da52c5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9198bf58f0ef227ab87516f77208612602e97030fd0ff8f8f7f746b9039b0e004446bf1fdbf4bef52668e305a00a4635d5de921d538c88de7cbd012be;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e3d47fe17ca452025b7056d0601cbc5ba78f3cca01a6e7c533fbfe0228338a29695b8be541af4264617c3a9a7470e34a0f845f122310e9eec14f1097;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b238437c6e12cb6c4476c1a17f6fe2d2037d87660a6ba512e0b6bae47022c86197a330ee65c62d46ad3b1644f8ce8369b565cf07197b1feaae93fc17;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a60de72e545613a0e15de96f04a8a1a5e290f5dbb451ff29e32c9253c86b4fde9b3320aa442ff63ead08d886e45255c317c41911a79ba3a3486ceac3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a47daac387288d83af1339c1c39162ea895dd3323441ab32a864a1835322a40835e230e109a6869fe91ef1485370f0b3773abfd16ecc245607d3d0ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbba7088fe644d006fef5f0b376b45f21b5c4c221f4513363e55b76f99bd0222cf7430b3a4ecd8065f09089e710f4fcd6eb53b8cd95e6efe71e90e07e2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c180bcc149876c926f9aba53273a733541e44ec3341a06dcd27843b98d850912ea721c0df50c4d6b0d44ac6db38c55409d32d201487b169fe68f7be2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d0be3a2dcecb4bc0805b875168347c486bc7c4d696665e783cb5035e71cf37ec6924f80e6557057e355efe9ddaf6069f48507a80c687e32bb50eb337;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h285bc98ab6650288e58f498f0090f6d7016fb86068ad5372af327217704bdb18c4a37a9a8a0fc2a07f491cbc00f621c1b7a41f716e8c0cb4d50f3e35b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf756575fc9ed8a69037576c2922af843f07975d5819e8577385e4f8a38be3bf448953f192e31d1998506f2c0be5c45d128b167ef599f654735c48245;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcaa5c1fc101fd1c18f35124a26669d3aa42d5bd9aab036afbb3774e353919de239f0742e8e140b941a505fb5a8cdf12824cca4bddbbd7f1f8ae7aee86;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h38f9fda6505c5b867087f2c08d8e8b485302e5bf4f02f50f51fb830b16b29b261b17b433778335960645ef3d93a9c18f9484515f729e23ae20fa11e00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2cae6c103103c954272d950d3249aeb43cae276dc713ef190d00a539ca6939a32b71ee3e70dffa98a75ee4874f9fc929806ffd07da2ba55404877e3d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19405df505b272097d7acbc1e600d784bda5d29d0655f6e645127c3ff68b51893919c51445e8c08ec8943e1ca271f585ef67fa87097268ef09116e227;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7382adc7ff2dc75197ceaaa397c29c5fd958fcb1642086a09262f0fdfff31db6d9522ab141e30c2c4ffc7916ab2277d6dd7e08b8844fa47bbc44a6c71;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b575464bdde39fdbead0c5dd5ca97382599dab0cd4e1cc9d2d124acccbd0f411b39c0959eba05833cdd0bfd2650a3b95dc997df84bea5df413f9fd54;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86b478cac3d34c1008d00bf29a0e0671b0fbe23c9fcdffc5b5ff9cc5837bb433f715e178de01c24bf4d8ae59b3e0073dcebcf288446694db2b9e9ab02;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13d6ab1806680dd2df0dc0970a3f8e9fde050c7e85e9ba6d1bc2db09ae5b240fe1661f84cc2f65ae817b9d8aa0c5527afab90a4d9b8e413f73bdadfad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4925804e95c1a37c8379c3ac3329fa5a9b15ba8162a29fbd8977e060dc8497b8eadf5a6bf31cea8941139785a7efedaf615356115ed6921264f2b1c7d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdac41a065a9899476b6e78a00df8c84aef87672357819b1961a40ed1dbe79bc8e813abb6d4955b69c563acd077688fef0ed412278108f4365e4dbbd13;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcfb0a09f1496e92ea67268d561069951b755148ff42930a5d70715856b0e551e9427da0b68d5ba1832a320515082055206447287fd119bb0af77efa67;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee9a91580e0a6765b452f392796246f0c203cf8f228e507fef8307d44357396fb899adc724fa82aa06cc367a282b4d43d92002b6df982f4f04caefd3a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8f760b57fa79804033fe1e2d2fee702d69cc450e9deea26ee351eb5125f67ffe2afde4ad0fcd6ed07888f1b7781bf9a78f56b60eea84db4878cb8f71;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc9a8ac2a25515fdc089253cf61a299d957c58b46626286c04e47d2c68335e6206ff60ebb0e59f264348764c1e1443e8381f5eda378f264e5bd9cf766;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf64edd20ced8bf44f154bd910e6ad8e3500477fdefc9e96302115b291be23fe70e197f6f99bc1d651a8a676003029b42740bd8c91b1f3bd8417379591;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a3bde433358e3a6a3bb3d944c9b5ad06e197bd08da94de3d4fbd5846491bddb3ba0adbaace7759104afbfef314f8943e70d67fd9fed85eaffbb75d60;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0d435753e2beeeda848390e502f5b836df2cd7fd8326ac02144bd0ca1bb941ca75bdb323b2acc69dc925abc8f95d46b254c489557d2f86c3b76c818d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f91a46ce504f20e59bacf5806528124b966db73fe52b917d92395d8f64328bd07dc07d21c75e226c78aca83221d9e937367d37dbedb8c21448dda8c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h896f01bdb155398635b2c50c314147d6498d9ec09a41c566eddd0c837e9594868c3e556b7a22a3c030f4c2bc363e1b000f03ca154456dcc6782f7e7d3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8130461015dd80adae288a143103c1b245820827a90afe5b396de3353cfce90ae48ca058a24b23ad19d33ae1ff992c578330f34fc46dec39255ecd559;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha943406c556111eeceb432c39d459789fea000d988508078ff8d84807aa15fd27ad56ae3232ff2737f94a0afe9dad0b8b71b73f36f2289bd01894c09d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a80709e1aa7ee4b28853ba71cd315fd08ff1ad41a3495228a3cd2f98767a0f0dfebe0662974d1d16bb130561f261dbc40a7b7d1878271cc2b98dbd5b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf91c1ca919f95ad7ea07d9072bf5614303e5b27dc090f9cb0214105baa0dd7b03bd8dc5bdc5926bed19140d2de1587c15a28c854685c51a26cb921e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c5f4b31dc09b43cd60048d4e8829e5e8a894c0594b1dfe177690e0d44aa8e267df35a72474ee1c8400b10c24ba8862a90b696a8bdf63b83c7dddd735;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7556a5af1ba53f89567f02dbf7164e65157d7319734287a21e73e2ccb301977fb4ed205a9da15405273b08f52655ab8e8011c6f0b315f37d5ed516c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9b8e5df792419961f9344d3528befcf48dfee1fe119c18378cf0b752d4c81549db606d945cb3a522058ac341998d810bec557cbb68e508ef91d1aaac;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85356c5f5c95195d801687070d4b880b81831899df84c76496738be8f7e7f03097466ed205753adde1b50cc8517ef7bd81a6b90227a670d254dc76d6c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h959507a59ac86a19bf08e267f118d231bd78d350f9c192c9c377cebfb1d9490d6bce219cce8fca77a171d791e11b8f3f3750b1e1f553bdbb1a2c22f7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e031a71d37ee3b9989037a89f5886409b3c2276d3d8d2f87e5ca4efa96c4cb0eab51ce69c801fa6bf661eede48cc44d442624c1c6c91d9c27f0a2832;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf61cc1ec90e371969cf9d65cb0838131522751ee7cf38e857b2b2fc8a81927df094875c5614cde770a369c85e8027a301bf0e52375509890f81d5ce6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h800217a46e75a4cb41d04d21745251bae35a81cb39b23aa7b0bf2d8bd6aa53297f1418ec009e11285deb58b2ef625028400ffcfc7197bfe5498b0dac5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f1672aa7ba13366cce78f6f3cc1a1ed57043c5b8b9a92a458df373e2f285c5c694de0d2d8ded9b8f6da852b0c5c5addf6a7f242a5dcf0e86ad9c4bae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b62b5f8023d42dfbdc9915dfcc8d23820fa3ed46513cdd6548fae339e5f7dd5e5f0f8f4e103f9f45b0bd090057d6298af23891f35dd299b44fe58052;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha680f8ddbd5f1196d412ef30cfc6451337e86c5516b459339d5cbdd671373d16b6d1fd175c9e4bb557630d91b00fd2ba86efa3d5b4aeee0f3b6e7dad3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdfe154cd09d41ce18f22a78ee791c5deac1034a61aa532a03e2f98114f5ae9b86d8180506ba7b0be8338340a4585070c116ff5df2e6ada54066e85e98;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd063877f5b22a6d9440f79ef5673d71e1ce0086d3c597b864828c5694493d7ceb52cee9b8fa993b40e99148e669f83b2eda68ad31ea43a9b3e869b7c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84d7344af36bfdf2c7e22d904206751f949e365e8c3b62ef345eb983b9fcd05c89de518efad2f7fbd510022a54c166b4c04d518bb65552a73d22d982a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb422192e0cef62b78522c4275657f93ef36035a74e429eee03d85640c55d36c1509af0beab6b49ceba0eeec08414445a24499f51b246fb2379d91cb32;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ffd44958cef6a5b4b43312387de578e625b9b3c269a503418708b7aa764dbb46d98719a2fd45ee1acbd003366554699bc69fa4e6aef3fc5ba5864bcf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6de64cc376a54a403c72564aaf6771d02c1a3839b451d05e93c2d7b4574f22974b6b4a24a453af035bbfa6fa10583cb15da66d1ffd1720a4509b83703;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbc22e5e0b0b8054982814e29ecd696cf8866fd508c8456419ed1593aaad4bd6e46ae18b335c37d47def66551b33c301139aec90b670ecd47b3d95797;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec6eabc3fb84cc0bfce651e801d3354ff471bcff57206d17695d78c604a3f8c786c5b4e9ced49ba0e00626950310396ab4f03e04cbf021f8caa620fd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4854b59eba5bfa0f4a99a5ce3dd7fadf1ebae9876ec8415b75b77745f009696491f3600ce0dcb2cd122109e6bfd4868781e835780bb67836cd270bb13;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h634f38577ced5ab498e19e58978f908a4efd79a4a535081bd9de5c6a24e4f36c9f5cd8388a87ffc793f58765a9fe1034c4d39c1b156e553ee14ba3517;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed8ac9648d56e068bc2339eb4775dee147d3d54b81e94060bc8279f0a56808e7c6c31fe1e987189ced0f28e8253996b9a23a1095f4f3be7f0752b6e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbf7c5bbe16063b2527aef6f451bd02893c3d144834344e112823079b4430e3c566c24dca3b4fb7c5c6d7340a441abbeaea32b8172b6de613ad0effc72;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcc21074ea760ed8461535cecd68d0960f79e10f9b51bf451b44b1a7699a1fcea2101dbb7be3c3d0dedda6a4384b5da26202f25958c5f912f27043e1a2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35e7aa28e1d2fab297f9e0acd4d4024e09329f7b451f48a249a322592a8c647dccb089abd50f8556474e0ab34c7af03eaa30ab1e68f12d5a34af29736;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb7a80fa35d2a400ee135a41dae04acdfee0047ee5ab7476f3cb31022892b420c3e17262dea1c3efbce2c42bbaa692134ef91f5450a77c32aa3c16003;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67a35bd0e719fdeef06f7440a082d40c5aa7a916b5e1081b357e13a047a6fc8ac088a2995308ab517cea84b14ca55aab15a1375b05fa1bdb313d8c6be;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f0b8ed65ab0870116061a583d5e0cafa301ffbcf1d011605b369001f1d830f33154eaaa3ad877333757fa4789ba1f4c94346d3ef4d6b02a2dcfcfc86;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52d4d6fcd49ec858bd44adff6d2caf4029c2fc198291531ca9875b0f7f30aa149e7ef566cf3eddcd67fbeb0a694797ff853a2e2d76a218a3e76a92a6b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65d415c2d13e91e4cc623b51638ce053ca532242556a67f5f5815de6f11a574086b5cb3ef579f98c8fdb2cc00e43404af5ea48f48d88a221029a1e993;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f507144f817fc97280831311a0102d2ae402a194afbab1d3ce6553bc9fc0ee9e2885a69ffed7a3ea1d430fa162d67e3e3e1b0da99824de85dda6fc8e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa091bfb80cd25d2a4038a84df8bcb62e9b2d47342642fff07497c69fedf42be43fdbb985378bec416f9298e1df687d1b0078010a5955e767fd866eae;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84853322d653ce11e7f366c50172fa0a686616bd55183340aeffed600fa4123f53aa0553393faa9d8309c8ad4306fcf14a966de68486500f33696539d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed970378742b8e042ca513df6b51e8a29f872f1d9b7c24b99f91dfdadb9f0f3f15c33f1867116a21bdfe2cd54094a9249c3353fb75c1c8e08b5b14b65;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc143481f9d8f900e81aebb87d17242e3456ca5d2783530a1d23e726357f380d4e0cc70e7d1cc00f74268dc16f2ccc95e56fe974688e687f63bf2f0346;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf941ee51b08b4b9cad01a62fa2b90fe435a20743776e9b88044bf93b2542af1cd13c89470abec49013e0d0aee817b07e9f36aa1bd91dfce8c6391dc3c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd5efe468f7e02017d893ddc93e25fe4400a809fa61486558cad9ee07d1bd8441f111ae278554aa397a8ce8de98d6353382007e16ea3bc8f9fa709a27;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf072e1da7b29a3bf0f203c7ac069c272c256716a8606dcb77faaa00ecde951d728de65a30a702c75b385e7c2e1e08934976e0af4a3701232d40abafb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85174a1069c169e3d3d58b15ce49f4e8c24c06f934d34f7a5aa4f84389b725f494baa670585bbe0fcb975f12b04b64245704ca2712c781e584802128d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46c42ab61526bf2b7bbacaeb1d41243b9b2996d832bbaad022e4b7d3a77c044002a3c8f10c737c15fc756c62ba61125982a9e9393dab0d1c13b6eb7b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1fb706d57f1a03484a28bd1f702c493a0192f298186e1358a574748c8225fb6de2527effe0d6aeb4c548940455bc24253d945d62a6b68de28383e6ad;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9f0423c8c462be5f8e35c6d1c978d63c9e7795bc7f234df7f605453f1451cd4c09ce66a7010835cada70e4d5b8849acba2f16706e34373c8742169469;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h969811b8085d0485589d52d023ca71e89e3b43b4ec4c5bb315259ef9912810899de4169bdcc0207178239e773cd01e623e0a3ad4cd5c9e472ef4f5c85;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h295a2273c97b1e3863249d09dd1abba7e2e9f481859d229541bed9ad1a9c1d4bd57edb762ee7a4746fb0c7b95880e888f67e8df33fa021d0bd7a13f00;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f8c73c5faade626e21db87f2f05da764989429a33ac11674c56544c2b42ca2e700605d2e6fcb16dac80c3670faf4ec8c620b6ad90b2d717a2af9e2e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9bdb0d83857281122d1b8c0f9ee09acf69944ebf1a8eb0a6b775b2e04aeb61a286373e288041d080f0bddd6736b9ae778cd4dd1a1def8bf4923df804;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0380cf73b2c4eefa2e51e00f73b4574abf1ff54c3dd641257e44af04782eb4db539cc8fd08c491b0af1dcdec3ccc379cca14965e2a407bc0cddacde;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7410e1d15253835a129e5d565b220071b04c54f87027c0bf78cabd19c403e0597cb3954da7500055556aabc9542d3de3c5775a27ff9de729cbbcd2933;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8bea51c6be39105e380bf7a13d0ac89ead083aae244211d6fed8859c5bdf3483d0abb589eb32967a9634ec223950a803a735033f180d67f267f3e118;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ae5fb76f340dff0c1b667f008458912c15167774b2e051853f03b35270e0da14fe2b59931ca6d2eb43666b0cecf13be822a29023ead30cc5a01e26a6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74146892f12af4aa3ebc67043d1b69ac138e241fb2be6d69401c6745272eb70106f4be467e960e40df036b0d19cc10d6e4930cd4521aa28f5be4515b0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa38205bd844b75868d05dddba73f966339aa3665e5a14f87532b8404d8864e3b13229a26c5c93482c1ec9252553251ff7ee9556ddc8c48d369cf0fec;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc11cff64baf4424d4f7a48a0cd7327aeccfe487d4d84fcbc3dad9533485f685f0824102b47de8c4786cbf4874947eb529a0834e54d17d8fe93833cf12;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93e03a7e8164c6c67e7652554c0c213b7d63bb19c4495b1cb3b8dfb6e4ed9e6ebbd68fe6b8b18e4cf9ab216aa8fdfd3a7f8efba3cbed7aed1c8473636;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3a522370116d4c199516a47960199f85e1c2eb5dcb774bfd61356b3682974eb4b93a207104e97613af1a68458950838fa9072d01f34bd2fe444ef615;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he50eb3b00685deef48e100fd6e1063e4136c0c690982de84f5a42794876ad5e11a952182bd2a7bc314d99ef48fb3ab87d0cdb86112db1822dba9e44dd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4a975dca1058f848af74542467d201832ab70720b4c0244c32e033387bc708532d99b71675b674e5326b0260715edb20b21c0581262ac2f4d9b512565;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6d66f55ca1c3b4d448bdebe7c4bb731d4ff314e68c50fcc9fa4ecdf38dc735c7962e63992ca1b1cb495a8d9a4842f240afe2ab7c98e4fd73f10b68785;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc3ce9242ca5643f3bba939d9ed5edfa30c039bb0121ad785d9fc4bd3c19017bfca53c147678cd37d3840a0ff21f0aa066678f06a9a2d538ebaebe06ff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcda401f7c4266dd9df257c5b2ff2bdfde65986c67741916a8c55fa547790be1a39495d88153d6c34396ef1d9e02a6eb782a810823c38d27e4a6def04b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0ed4356a72aefcc1200972baae3f8aafaf65e89a2abac70411c33dc6123fa7ddb58e588259bc95676e1f93639d21251049d835f01ab82045cfaae350;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he60d29802f663ab268b8459cd531006e11ec80c9697cbd1f30255f6746e2e80a84adfa7a96209bbe2466dc36cd9b938f60b883b41b5f7eb3f6eef277d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hea3231080698c7cda29d2f54ae70a89c5b8dca4822b62a739c0661ea6c02feecc7c4e92e25773bc53726d284a4e90d8f11be14508094ef23df850c0f8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52d0ed711c357aca6d174cde193f2b9f0eaee6e564e2c21295f7befb57ceffcbc316531415afbff70c486c2f9d2248a1951fcf9e5b47b0fb64be8a62d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8f40b188299247e941339e22ea3f51ea2f12645f8c9f0bbd42a6429d94a27e9e0b85d54406724fc12d4c1d4dd92e88a28dc2ad1d07bfe459de34d3fc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f06488fa329cd3adcc8506d07d926a3261484cab1ce0d958c7cceefb53052e7afdc157e515be800d32bd5acb3a4513c0f4d5b4a4b58ec67f64aea4ff;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha58512fd3090e507a6e8699be03facd94318c639c087f18f812a4179105405c00079cb4b48e4135f78b33fcbd0197df886864fe79c619061d8be23108;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2163890d46232b38c17c329130a04c9053ab97d8212af8c22b39bb7102629b2c80c9b3069647358c9df08605093dcc1ae2754bb09fbffd7ca5fbd19fb;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h290113aff5e00f8586f5949178e56e3f8f74830e0505e2a4122e2006d2f4d99a0690b76ff7559a0024e4b26f1ee04340ae096064ef51bfbb921715ea9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48dfc293b39cd8ac9846e0216c24a1c45b6e654e03526759f4d4118329af302ab2ffe0d0de2df1f1cb5f1c08de4dad17c9daa09e1f1e6e3b3a8c4f116;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h522f6a68f7fb4a5bf76827e907f42167a2e937b9bc0257dda393e94ce32f3bda24900447fe043b2fdd616d794017a0b029f07dccaad8c607dd0d49d30;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e59380da96bb9cf3fb06f297f2aa35cde150709e1ed0261d1e4a4a5268b906917e454bf9a0479f82c59c3470ee3feec27bcec78d65f1170d8558b828;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfcd64ca734b3c5a61b46f080f3aa334303575d73f641d0eb30b92ca2eef1bd71118f80788d1c4f819d8b31cb20b308e179334ff2cd402709e64aa2221;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9786db7502d20ca5d8ffa392dd68ffaf2d4ce0d553929c70fde08ba885e0d3a74a9d208e392e9cdc4ac9dbd1b324466dc95eb6e06acf044604c9393d;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71f75118b5520e21e6df09dfdf5b9797f6c176a2f6d32a12e7e64fcc584762d0b11d0f284c43ca878518fa7b8d57c847688c1bd1189f15ec84aca1642;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6264db2e7054c079e6b1923dcc620d55f381b5073e856c5dfab62ebc6af83d5b13a9d75038167458a16560e3f92df8a8920d8545e60b05f1e0736eef6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3e5abcd947dd625fcfd09389f4d94f26a30c703bc5b743dbe66be8813109ce034affb8b489cd7506b88e411a050f7563757df7eaeac0d4d60879d88a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he04b186d0378d7b0b13979e1be97ae8615b0746ace0c1f13db6fc9720282feec94eb9d90d862de7957954d77402ca3df58dea139255af74451353a6b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80d0a9e8a4fbd752e76566bc778ea638b8311595f878c9b862db73636fcad769feba48eedddc32d0fbff69fb4b54353ad72193c104f3f61c64307796c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5b38b122e2faba2da20dad8330a4f17fe84a219a6d827406f21e7cadae5cf26b037992f35cbc57c79d34e35df30fee9d39d9b2f02b4b16003384f375;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1873e93deec4003ff57bc1f8d9000a1016ee06bd7622f721d76a7559a6c9cd3a233a16f6197928e16b3485bcf93fb3e77e5ad2b773b1a0ae858414edc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a6ad9c50c19b1821d7c8b08cc472e05f859581f98fb19d0676078a46b85b8752832fba089c68a2830e8bea11ca4f6d02b6b66bd3533d46346812ab01;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdf4f2b7ecce6258ed48c1ab9ab2ebdca85cc9aa685d7eb3d32e72974434d363454679eb8495e33ca0d3962b438874d2cdcc340ff33adce35a9b2d5ea;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc071a6ddd441534e323f9891ddd97585b791a05d975d0ed491f31af08d59db1b15e8fd8ac2dff68c6185fbd318460a370ebcbcaaa18d50141ee6aa8b5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5b0b62ad941c1e331934895ae3b9cb222487207ae65b878a0d018c96e04affff40774dc1cef277b27b89659d961f88d6daf5191c5062be57ec809b04;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha14b682e14f5629d7b4e4fe966bf6256294df35bf5404ee43b72b7af90ddb24e4275a4cd655d233b31fec6368dd08257251aca16f049f239613d5bd39;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79c43dfdec83237a9cfae9c443a1dc01ccf55eeeb65347bf6f8fe6f9a792e6a20ffe6b5cfe4d2b89cdd500b65c4fb54aa8ab6198472938d8dfa77a8e1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9ca6024791eef4fa7b1df053621a1cad294a03fd9cd8f8c1d9bf2fe0b7b79c46fa365f44061514c2ac4f93f290fd321a14279ebc7816607f278792bf;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d2fa04b6cd31cbf0fb42a63afe1f80a4aa501dd2b7491a494b4f5888416de3156da0eb210376200229b6403a4969ea0046c447932fa21923000b673;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h676ed229afa5fd6e7ffbffe4ffcdd2dc8e9eabcd6ef6099b865b22f902152ccba7dee74bcae4bd1ddb289a4978eaad003858677420965ed50e215f664;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf092176f91eabd4a188c897a42d12e0111682501d7b040401466cb0bf06a1ebbf9b7d25a1d0e931014dab1419d64fdf5c48d01baaa4442ab8ae95c4e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ac216a0bd984bc604f02a487ceef6a5698a54fe08bd46cce5c7e92fbe77d97d439b97dd3c57ffe7d0c35ac2710eda814c428c890be1b8e201d15abf9;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bdd3f96c61720cc8953ccab082fae16ccdb32aad8a34b225876b07a7a4a61500fd372211c9deb2fd2915b10962fda0c504aca655759a0e2a8df42a5;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h364fe75eeba6476d192cc27b56cce7cd0e4b2bc34d2e06dcfc352596a2ff5aae82985f300900c49a32c11b631df269302c97778c5358e69697881e8a3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8a67442ea655676e377c4de6853ef9c66583e17460b6a8d42e14133c408c842eeb147853902cf981db6ea76398221dfa1777eb9360c2c65627f6f298;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bcbe17f6b23afcc0fa0bb8a2cf4b8335d26fb8f0505b3f05cc93ab7ca100fc26f12d8d6fd92c197962d89a27e93a596b70cdc0b3914da5ce103d72c3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46400caca3b181063032131780adc541d0e48b038f41e28f8024224ddad342ca0c1cdad7d6281023f4f45c544d6437517164e7b362514d855c2b74328;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h879bfb749f858d746a2f0265ce6f51e1d50b459d8aa1f7516f41581a8afd8ac7d15abeef665004afe4fc62b54720ac424a8956d47a95ca2b1e2432898;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h397f766f0a82ebce10bde17f4cd432a44ef1fd16d4d918048f4131985b818da896aded220852c9f33d97462d19009e2944f094413673f6521273f9c93;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f9da131e6a3a1c4e249519cf6c2951ed22f7616f0d18f4790242d97fde841498a62e29f162de40ccf86462416e3c1520bb310a8946a14e7a2da54e61;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde8a5b6d212bcde7a48cdbcf3a27e928c0b4a8b1b44b84067b4a6d8151f0f3739de11bb5e17c6d7d64d7a640d1dbeb1dc0d7d9bd45b8896e7cf78b1e8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f5f2c7f447f40e907f320b914505b752d29d4bcba5d80e9a18fb39b164c66eee4ee8e79b8aed603dafdfd4fea94dff8608e2d6aef9491d092fd946a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8634aa9f4e83d910b26a657c4e2c1d7a30ffb32d701103e55186f2119be144dcb4683869bb952186ab0edd5ff8d96b7f102b1ac9cfbed709d0aea2c33;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35c2f87926bb64b7be920b0e18cb75edb60e0ea19d9358ddf91e8699fb11f9bf46202bb2e1213e24a9c04ef6b1c017359ac7c3b41de446d53668c50e3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0e60d9609d708cbf8a057e7804a0130ee0cc74c66498a7453322b88e3285babbb2116c2d94b318513bc48919c1154244681f48c9a72101b22fd7ee2c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28d5220ff59120fcc287a2c13cdcc681c11bcb77199314597f1f0e599d705dcc05d1ba8458c571ae3644ef49f67d18605f16f251c0b29ff3414932c3e;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hca79a3dbbe77fc12674ed60e7ac3d25aeaa942abceb7e8c8b9a902b3b437493b28bce6aa4fff6d3ee01b0aed006976bf75f5e5d76507bc90fefa152cc;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd57ca0a55975c5194c3fb82f3600cc424ead2349d5c693126151505467e2482065f340eec672ced36f95b91c1416de690efce8006354ef2544c58b3dd;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h628a39b22ce6af5dde6665a3d8fb71acf5345d7109da1360e215d927fc1beccf5d1da054d2b54ef976fabdcfe27b939ee960ed2d9340d0c9b1d597107;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31809446499a4ae99f7f71483fd89f31436d9a20d5400bc709f4ab001c472f1d8e8b6850147a74f3eb0f744687eb6c39dfae546a445c9b56e3d4687da;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d2aee291f7e5e535976dfdbd2c4adeabae977be98cfab07e2e8876685efd2f66bd390eb07d1fd782e27dcb245db01aaa941d163004203d5724ead46a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3473461aab98a729e2928ae7c0aee4cef19fd42f4cc58bc1cf0d15e8629d56950e6bd9c76518b13a1dc9650f7d53b5cddaf73add092d04501e5731bd2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46d8e6a850a7462c1256fee77a642dcc24a7cface4c0caf542aa9a6a06696120337edd9f95a321979d79c40066ef60d5220de3287f2061ece84c1f541;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbc82ec262464571087dacee293ee202fd58cebba1dba6f08b185073335f865f8cb33ba95bf3f768ae49e4e93850cc325c61baeb34bc0693ef44fb5162;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ed3f3de24411755e58b68796964b9396d62aa37d7b600ce9600f40b75d8808c1f87854a4fdc6071eb3dd4b8ea4d525eae5f83460d2d249db2b6b1ca8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52191365cdd300354731d9f530e9ca2c9ee126e0d061ba7640402989980a7ef2b255b8d314b0756173ea628b6f7e1cbd1669bc0f4948cccd5e7a7e090;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h606c3fdbe52a09c41c2e64e8cc1f7a46d786d782e5dbe7e029310ba22de0851657373bf1baaf0c09cda5f30289e047eb5538a3a5dbc8a6ce0ba9c37a0;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba0de0c9a7a4015160b2625c0666c3b081d9b86f5bbda4863cc92bca744b628088c5d92723f9c15f72ccba6ca777ebd825c7942f00ef9d0ac5caa79e6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d2858d57b5bcd690435692e4647de710db98fb1d0b11a8dc11e47bfc6acc0b02c2f775c8b310f4734a009cefdb516183db0e1dd13e8db8d8c2b7dc66;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4eea0eda6eb1415751c99e41b802eee9f934e295c0280be0ed0aba64c61a294d8196bba391bfc46f208d62e2848c9eadf7d9191e7108ca1b0870695f;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h538bc01e8a788fa24fb742072c28f2f4994dc0acd345df95280062647592457620d2ba8a0ffe2eaa85151f5387153b2b2c2ad8c4b08f80bd69e812c67;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd7f6cf199ea2abba3b9f87b660d69874a2a314165aba446c767d6cdcdfefa70285c740326435f310b708e980e65b5acfc6a86dd01e841489683c7196;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92cddbee5119dc3e7b13c403b70de6bf222d3764291316f34b43a7c49dd8eef1345b86b7dd3f905c0b9729a70cdc0cfb7d381663216f4f3de15c522d1;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6683ba20406fe2469395ef2a56c9adae0199c29239d10fc0511b3a098a90caa1f5e0887038973b3d2949cf089efb307f51dcafce27ae54d2c6895a06;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fc46cef75d97603d74a4c8aae94ea4e6c8b62eaae1740e832dff926675481469859d18e73f2f9d3fc7c5e23671643f46bf3a0ef02b7e9c046119d23c;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h418546dcd9dc5e85ec11e0def0b319c20f6d3edcf05016a9f233ccb227957e72b8b62fdcf06533a9a2e61a5fc6c1f2443e900b09a6bc3fd4607ff9740;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44886a25c2d696f3194e466ab273641d4593e2076f4b43df6600625f03f73af7dba3cc063d4b6d21ae0b38197e81b0566fa482fb897be13ef2cf3a198;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8f4a1f3aa935feb7bdcddbde28dfa03985a758128bfe12cfbd08d4ad5209b97111d04f5baa0402339534a5e6ca083f0a9731d3898f43eefdf5d8f0b7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53581ce1513116becead07c68f50e0c86ead9696855e855ae519a60a304a12f97081771c70054c7e5455d0ee99f2a9b9fba17d929386da4cd142c34c8;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9987f62027d52a15bcaa013a494340c5ccd343bdc47d7d17c34715ffd70cd38d11c64fe7641da33e2a7e50d2b61ffa0da5ac3a3fb5b03399d9ef4fc7;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74bf113520e057c65a1095665d4fe6ae3659766231691b5b1acca7228bb1124f4b30a159a287ac43dea0619205fe4ac4ff19d6e38417ffac9e1560e45;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3390ede262af3e177d6b81f93bf9c568141f36aa7bb9eb3f425d243fbd913d13b3d80eed1be91fafce6cb5138ed8ac46bbec5e962f41a4d31bee1e36b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hded3138dd8289e27cb6b97e027156b9ec6a2ef707931374bf29797eba10bfcb82125c2ac206c3e7057c2a42402583daa4d25588dc1c6886e971b08c27;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5fa585c22bd1bfcf1d2a9b4cea52f93c2770544fa9ddd373d7007201592c0c223662251fe179f8194ef4df105a39460ee0e0d0aa79acefcbdce07a9a;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf688d887935a27ab7baf65a0892e6ce2be2f777443bb6cf19225dc41c06b8b392474ed6b26699e27adabd7d18f3e1b0c94af94497ad232f4df52048c2;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a2fe2740c835b4f1c23b89c36c6327e499c990c022ebddcfb558481245e7e72121752f66b4de8e185109a47f648d8f34367095bc987bc2d399375213;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h813e4ef9f8d84a22f6724ed3054444e5cb9bdc594f9560d8788a8dc5af32dc4617aad6237351278a2c0414e54dbe52e71297f2addcfc4cf3267426c2b;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb5ad27316e07277374ad032a7938a66f59c97c11500054ba4a61435f578911d94c2987168112f04eea1d803f8a79c5f1c9d926642ab6facb613950b6;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ba8c402b5f99023b2515d809e4501a5faeae333a67d3cbed0bbbcfe2af96657fac980e7ca2bdd29a0e9de5b6c733f2ca82d6e92164dc09354c860449;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h60771cb0f35f70ee81478ffd33a93304435172b35742299cd693f52d4fd857232bbca5da5377695ad327aca70ba9e36de661cb44393db8c3f1a5a1c89;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd4085d7b1ae6dd19be8047c551cd33a458d9fac784852fe4cfa0e2f5d00a220a835f4e0fb63334a5105ac0f3519aa642fc89367ab02fa9e5cfa03e38;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73f399f34bceac816a69859db40da141310bacac736e029032ec423fd45a916d3a9e777dbf3bc047d5e09bae47126169ca37e767184918a555752e588;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55c250fccbffd99cc9c2496af94f329d4f727bdf8a4f6ae83ebac26be4c1558029e3cefb6101d63f1348e477ea858858930dff9af3727fe009c1537f3;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd545942974089e15e38696322f946217969131ac6379bb27a66bde77b6d9ff6d7afada1359d6131702a5cb7153b525d92b8c7c386e4d8b6679de78730;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he728f1d475a9f263abb22aaf16ae1a6d46ef6bd7ad66f07c0ba8e0bbed21cc8e749f6729bd51fb72c97d8aeb932ed3833a8e41f3d07a5ba80ad0dab51;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h727e02298dc26108014c347858021f5a4e834bc356edb8f522bfc65788f775b81f969a93891537c15754629d298c320cfc460ee998b74f1d20d28d1db;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb6866c7e1b9cb01f328a8832bbad1d94dcdfc646148977ca6caccdeb92d64e8e8fdd4580bb44fe8ccefa23ea77098cf5379d22feee96795f20157706;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd30f4c05845163ed52b05c07f339153b8cceb76ecf9c49838fab5640dc245700a6fd64841953645de71c4f82191d7f3c5bff4c04bf6c50cff9c86973;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd83ab369a74dbe5610e60c5ff8d0ac328d69577151a2435fb87cf1ab4b4d4dff8252e4708e23c3dc8d13e458e04045e83d72b33049066cca7ffe689c4;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd73379cbfd80eea6ed01ce3e0f1caaa2882ab3832075e438c609155dc1d212e10a76b4e7da3c273d3366c33056836122b1fbbccb8e242925e8e853a09;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h33abc4cab1f58c84c68b7d13af3ce3ebeb58968c1e5c0be18877337a105d7d196c3438711998a840cf804b443b176b16bfc5466ed20503d723b0a5f86;
        #1
        {src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7321cca4476b4093973e0c058f09156a5d1968914eeb9276a4a7d400f0d0971a9b7042361ee16111f8acd0d7d5806c8c550d401ae51eff56cb5c65406;
        #1
        $finish();
    end
endmodule
