module testbench();
    reg [19:0] src0;
    reg [19:0] src1;
    reg [19:0] src2;
    reg [19:0] src3;
    reg [19:0] src4;
    reg [19:0] src5;
    reg [19:0] src6;
    reg [19:0] src7;
    reg [19:0] src8;
    reg [19:0] src9;
    reg [19:0] src10;
    reg [19:0] src11;
    reg [19:0] src12;
    reg [19:0] src13;
    reg [19:0] src14;
    reg [19:0] src15;
    reg [19:0] src16;
    reg [19:0] src17;
    reg [19:0] src18;
    reg [19:0] src19;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [24:0] srcsum;
    wire [24:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hae69eac7ae8129126ca75d3094bd9a021c9f4e0adc0bc7bf0ff0fda7eae2366734242ad00e2b1745779988368b10e7feb692;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86cee8ec9cc52d1113d84f0f0bd22fe8f16736f7df2b2661e68010cf9c5b3122380b72de13718f22d3b8d4263cc57ebbbfe0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h422ca8c877428716a86639ec8313640da63a0d15a898fa19b8e508aa7a8b89f51498a5984441c5bb41d1103805dbe1d65d51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f84ca71dfcbad9e095bab9ae49a256a29494021f4e70c56c49086479ec3a9ec39fca5e89295f04df48519854ec98728d1d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5556519fdcaaab59d0c17269ed9983cae4d28a624b2efb0d77b7f6fda8014daf2151a21bd703803ecb9649acc76a073b0432;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5338d91ee799b7e3c91141744b97d3888f7047ae217a1f3f28ba1cbffe46b50eb28c7708ab674b6308c2b8d077b7cfccb6c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55229745c01d881dcdee3467710b4b42f350299332b1252b59581275a56de546c964ef2af9c1afd6f91e9158cefe5c499a72;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e755217b3fdb1f309b1a610b38a38b7ced06c8330a628aca69f34482a7380e0d220935cd9821cda8259cfff37c021ed8438;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf80d459da199b0ce692e7457bf807018da512f4310e9a287b6c6118c85a3d5afb8291d9ff0c30e9adc878b8b5f7d95f1530b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h307521c584859cedc2c8685e9c5c039a4234d4774004908d0f1744104354bcec1ee53e21c4b3855c362057395a32c0ac3975;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83ed032ce6d5d31ae4a0e1b5eb1fc1a5e50cbeefb64da5fccc72ba6ce0f3ef434a5dd74dac9a09b409ec20eb33bfac757746;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha4cea217865d64cb2b27a1ae47c6dde2ed6172747e514f472a4099cadb53dc29a5daed5a4fb3a31fbe6d3b9472562edfa761;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d391ac8e69f89b86d0e0eab5c1cab9c19b13415b101a68238dcc9f2b6c4c4f7f52b4f8656230e81cfa0ddced71110c69719;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ee63402b534e4d64bd84968c7af196ae92baa94509bfe118aeaa7c0c42d2c66dcd57686f0249e71bc78eb86076fa0f503f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc92bafab81bd362947ce9deb1e2024756e1a5e3b5458f7cced5b2cc26140564bfa65144261936c8304fd4f61f98e3cf9c692;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56b314df650c747305418c05bad4261e789892fe5d865777de4fcfa05d11fe6b555038d6e4855429c811b084c64201bb39cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a62adc89bb63c93feab5ae657d524ce6073acbbf38f8a243287f6e3f960922c713dbb9e92ee9961474194c9f4f6ca87aa9d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc61a7792ce54f59fe28efa24cc2cd4005b8a5c5a445b7a0ccbc99edcd4c2e90ceffbdebab64d6f8da57e235d3c499efc0f8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd75f13ad2944297bdc5c10d90522df376c2565913c32c0f028f29e316f07de7108663d5903cb73fa068562eb7497100801d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb88e8472233c9d2a0a5319cff5f218913bceaa45d386c08fe99ebcaa8bb9d3697c64e1ba4302e819551986785a6898cd6d87;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5153ccfb40ce1475a86db7b14ca1fc112c6b6b892b902ef90eb3f793163dc4d67f504facb6bc5bfd59c42e9e2a9ed3d520c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f9ae8d2edb90420745b866aa541ac3a55c313eb528ae374367652eb06b5f86416e72c5d9fe4c8e103e7dc01151cc26c9610;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf498c003b2156e7ebb143e6bb0f04912dd7842f2e65ed4c35b6c42e672f6d69196e1c3bce0ac9f4513a276103501932dbd7d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40143f24e47b9bbf5cee9143c7a84c07a54fea3f27c331884456b97a14622c546ef933e654123d2d027cc0d4c62129bf5a58;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdecf2ba916e6b00b17f08a0a0d657e5b5bace0d9ddcb1c9aa6667a16a85edd43b6b52e8b24445c5dd03ed4b042f9e1eca4f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86922a82c52ceaec392fe3dc98e06884d44f1ea0e2a5e9c649faa3c2b6b66603a4591a2b23459e0a26a0a3058b1a1a902648;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he22f3929ba149368cf25f386a0fe35f9bb72205cb67ae96318789ce66824726c1fcf8255f3e0c5aa4602e3e389c076630dea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84a2ed6b64eec26630f1a9593b2978ac50b9cb4a95215a742d1ba73eef147c5abd72e14a403129a31689da56e4b8caac6016;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2d46894179e5853ae697512ba3fe16780015c0bcaba40d738309e2b5d55635552058d1be35774f5e362d17bd5f1a686422eb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e0c250659c19704c79b4b44c477d7ceb5c42c63c678c9182961ba05dc87460f547360c1e8a1b877f5a274e44e8273a69447;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h883d5d5ac667bd03c1e45c857ce9684659aaf9cf1c20773e5684ec03866b47e57f770dbce12220050039a190dc00315760ae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdc4a0bc83097b75d35e5427caa30910f7f633b73d142c2c435d5e86fd2847e7ccf209eb880b09919d2bda3a06ffb54c7afa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66bb34f38e0d2dea68bc564bc006f7d0b5c75cea743acc3d04a762e0db5c66cf01b3a7a62cdce6af86450b852af91eab9907;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h713965f6a61f09e6ee304b3005579cefad2dfac92f9457ba5e507cebd8114723d06f36253fb9bc19c7b3aad2fd845b790f53;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e68be0b65cc70fb9148c4019a33f5927af2c1aed84ed592721e92188b908ad9ce1200c150faf025d6fc8f4228d8d477fac6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he689a0dcc9afd33fe4e9136255951ec0e50aa6699af5e2be92d866d5f63b209c32b986e853d8d486f9e09ecd4e8964fa56c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23ffceed7597dc51ffea2a1d92dc95095b1aa1d1e6ca47426a65a9f3526577e505cc7c1e88323130627db07a56fc67c98e79;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h46de2ed8774caa11b80e60ff9c1c5a8f0bf52ca235fd618766b91fddf8828d5a82d4d7398da4b014a7590a4cf45af88ce831;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha71c67ac2ca4ef8f4e383529af8c8a04e0d04087e7a23f5c7b977f966b947e8eaf1b98630943cbd7fb4fa2eb761d677e2050;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ec9a2bf3ce3b43dbcbafd56a9a982617c76f3b78b08d0f944a74d5ca4ba70b380014cf93b77b3d2cbf001647857666959b9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbc516a3c9627518691d92ef8f5a2dececda213e1e9182da120f1bd1a56fe02f2e1f42f7abb2872166ada4b28fa1b994d0ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5152e239397bef1d642823f714e254e6a7b8657c874efb904d47b11ca64bf2ed8163dd2fbc7c7a42574c4db801a49082c91;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf31fa309b316da698f4ba2a70452c66d1e893f64ce65c4ad8e7763f392c5c4dc96479da1da5d75d97c12e7f6f2ba9371f040;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b7f908e8935a8b94369b069f3fa3154ce2b7de4e825268d2149b7275daae2438ca84fcef61438055811483734ab426aff36;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9249aa013af4d8ba87bde304e05ab9932db8de094c02b7c34574098973c45f20be354997e13391cd4e7e71379cba0b4ddb85;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha424c37dad9ad501140c8cbd7074042a2192d5a930196216002a13146cc73af67719a892985778f12ac977a1229366305899;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e1daa81f660f6616e64f770f6b9edfb5b406e3016164faa6d4d5c6f4c685af68a9f661706e11074d16ad22ea7d137c37c37;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb7665717954be5ecb150fdcdd4488c31031979f4ca879c503a740f7e36dfa4be5ba264da5e7ed2be5668732f574cfe7d992;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37691b86d9a117fdeccdf2f2640ea12e35b35995a90f8bb39d58871bfe77de25dfc5e2f3c98c504b8d50f3bc4b332c9752c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf84b4fbdc63df928192e0778e8cd877ab39a85f4ccf6bcba8635ffbcb1a38a370624ebfd1f3edb0d3f8dcdf995f7aab4a275;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h259b26ce7d23031a252b2d582db9405edddd9f6f18ff7069f04d74aa0d356c191f2c69a909290e029a75b1751acb3db97159;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb699a956cf5d48242ff7fa088cf74a049d45a525cd967d9d93197c36f4b7a40f2e0511afeb339a9d6e4bf6f43be72cb08541;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h109cb217d8908303b83ecaf744277c1af23e1f9e78c7faf4a41a854165cb353ca0be1d5f1bbbb2487eda29aa6eeda5581e41;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he50432cf924cd2253b5bdc7004281d4997c934bd10ec43b7af47c6829c8ea333ae6fcb1c549a30dc4ed8152c8d30dc1d3b3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5df3978f25d5b07b9047cc65efdd7106629eda4c5b5cca506afbdcdcc3fa446d6a0f81c3b98346f96852c175cc55acc2a31e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d5929210051c5f1096f948246cad0cb62255e4f0824b57a9e710110555dfcc90c9d057111a3a5937b216744375e4c345f7f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0de766fbfcfe32b5bef7a6725a41ed92ff2f8ecfc7a9bd3a3405fa8d70cf9e2753f08c5d02e997f79c0f8b63da7defa7bf1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c0d72fed613c1acb6ee38fdc75a93bb7233a0ec2bd61813c3f9081d2bb033c29df4636d8233ff8e9962e39fb1e1a015776;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22f1c9dc9a7b2142cab75d9dc2bb1662a3d318545a8a2261e04fc83d5715ab4ffbf8a42e00fa80a7fc97fba59b7b42d743f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf79342c8eb39e3f129892e8712c0a10af6d4cd9009c1cd0548b608fb733fd3fb4161c3a64c8122accd89e9c1165316ea1900;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2ef38b858546e93ff98ecd61a04591841cf4b160ea1abc78eaa74d56f47ec6422fd2a012fae63c687a5410a292c7126880b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0f049a5eff74c0852003bd1d364d729ae73e28cbcc78d8a1989be5d93e13f72d84795e474b7c906380c0aea7d7fafe36a70;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50104316e51d8251343242df0b41413da5871776b087698c6ad7fbe66e1482a997b10832a23db14cae31a05c6646bbaea9d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcac401c535211d95032ecd3ba60b9c89a623a370aab112f293049b361c3e25c4ad9b1e50137adce2eb98404ab243a20b0de6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadb7b2a68644b40f128d6c0443f40bdc0a0023404ad1a3e8791a28cbbde0f4d6388a8e8cb08e10b5d73debd8e59ec8e5e99;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he4d3e7045946f6bb26269cdfdf269aa21af1fa3c235702eeb099f96302d561386f6572be32b87403d6e52e31b59b1340811a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc5946124f9abd60e22d4994e6a558868cf7b6b1d2863d5d1e33555d557667a1a4d46bebe07a0f006b89f407cd509636fa7a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58341f5d595fa254d35aed05400712b6828c392e01f8791634f5b9fd6b3fb60c83b0b3eb3edac626d6926c1c6a998ced7604;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha08aeacaf889b369a004bc9016032d8529f19ce93ff3f7087440b1fab741b8a27bb227dc7cf21c8bf8296ad84d86c02a66b7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57f2d9b39be3f3b678b99b8cad4afefcacc849a4d8845564b29d87169f1207c8b4bd85eaf50e9cec6a9955d331c1bf3f9485;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1fa3630bd483381d1243137713d35ceba4d6824a2b286b9124c904c8493e2cbe557dc57515a3a95990c3dc362df667a3558;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c8308d5994db57a79688ba07dff569504362a28022ffc832a2a1220aaddd2bb2b81ba13c7d1892d74d95bcc796cef8e2b67;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a6cba2f9feab13b6e5e7e6a80c6f23acc6129e03701236f6b165f73ca1033d987ec327b0d37728a82b24c5309fa8ce62b95;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2bde725d514f348844dce086497e05805748f10d7b3f982a949ae51a87d891cf633048ae1d5d8a62a0bd1ce3009869182788;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa5eaf12a970429b4f3ffc82bbdaa5144983d4fc8ddacfe8c79e5523320e701e314bf45b1928d28e2dda381d644ba30a14f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf659d09610bda9ad65a712f84d271c5eb886189dea5028b87ad9d8b6db881682e872cdb8270557e3e8ad1fef0fb5859b4c2c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde48e630f9d4cc5b62a995cb29e1d870a7ad3ed77d19d65a760c2c40174d615b2240d5128a97dc55077dd8c54672df1f6ec4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4bd2b9ec6712bf0ceb42fc6dc1e7e10c3d718e8b22963411d2fe9111f9cfe9af5e888dcaf3e0c5f0a562bf1b0d0561edffcd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h203604f12668946a841eb233e7ced486bb9aed1c3d39c044e3d8e0bbdeae1a3f2879cd43b0653aafa838ad1af33af3b0c341;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a5183bdba3a2f957a7fc6579fd55a7159bcabf5b9be0f5006487c78ded36273a2ba10e9b3335c31c4822ce71be5c1c23b09;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80b1cec85366c73183cc6bb4f7d1b811f1547cabaf45c054835179616c1e62af0d3f31a290b29b475b32437b4446973ee9f6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfec40e48b6a707799186bc4dfe0024c9ebe6107b8ffa03f6fbf9354654a14ca644bef9b7ef03c5518fb7cdd90005c35327a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha21efad344fdac2f414094426a51a25398eb78860d5a6817a98213486c43967cb4db8117220759851d43285eae2c702ec6d2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc64d966533d513b32c7ed4ef237002da2afc927820853c19ddf971c8873fb33c2d21cd65fa81fcd38182941d2bb63392e1a1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a7d0477c8f3b208b65bc0ad4d584bfd85163c73ab984cb2880578866f2353b0b618d91888091fb360892a731b6392a88f8e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1294dcef3785d85aea1a5cfa7849181bdba23de65c0cd57f53a30f86bc0f316e7e81a1c190248ef9e5859f2ae34319265592;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c2a6dec27fc08ba85b6ec95099dca3e68949c285c8e6e9f9d15cd7e63c62b709d422e9143ffe85adcb24c3e746fcc8720c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h327902585f212d1a3d310ce9b48264ecc15c31fe7b9cc05b86381253a0edb4cf4bf896241014cab01f475a4dfaadf64b4356;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e5d13a6ecb6b2fc3cd616e06a78a5d73db6f4a205d6c561220846bab7728f7f425ea79d479340f58beb585b7872933092b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haac35dc0c85cd6d4dcdd5def99b2d4213fd54d1522bef5aac8d767ed0c3b9e039147770144c9996d75ba89f45e8c19caa3af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc2a1185c9a8a921c01679ee28a0c0279dd464769103e7c637566b1c61db7793148b8ed858384215423800438fb9eb90fed6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b81ad7277010281c7fa486467de4fbe836f6f88c5a08836315f0d4347273c56edc24fe90034f1568f3e152d210c7956f5af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c08752cc64a5c5c33003e457e8fa51959a48abc5c5bd116829011eb293220b17fd2bb9c474f1ef916c6979d55cbdfa11d4e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27a221eb65253d82b905c86201ac0965ca1836f3ab9432e06b26452424625ee341e2019de896aadc3b1f343da60014b9297;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdaf7d9d6035485b56d5ee211d7fa0bc8c917237c666f75c46c108de16ec02c46844e6f0dea8c6aad0e2894fc0a0593618572;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9f6037907d9ece8a3090fd95101f8507ebc58d28355795aed376cff1a7271862e8517fd46c9bf7c2e77c6e90bff3372ac4e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h437f017627183a35a39be00810ab2a528cd8a9d7b7e711c43d7f8bded6f501a0770aa136de506caf981d18e9c27ef766a0e8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8316ebfbbd57f0a762f4c4d67625b29f4c5d7890fa19c085ce2d4fa69e49281cdc82efc525d77dd3c224323840b228534371;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f46ee558abde430e609284d9e230801d740b798ef1821f4650e495a59a0401fae55132158dc4df7dbce5bb8236758ef3a28;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7aaf8ab1ed7bf0acc3a6381e4744e8731d850ff43b14f1ce1145660ef3141e2fba69debbb5ff6608b3c81ba2d39b9198f844;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a2f280c1b2e1d670a9a81059832f3fc87b0d8784661d32223c853408d4ba0ca46a7ea19b20e75f7b5cb6166e31ae9d5766;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfd708e4ede2b7e5a64463c50428996bc2e0e0d78b96292d2d30aeadd7bcd053d3d92bd203e02b5424fdad40b6372e26df9b2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6dc2565250dfb7b492ab37b8d044d7488c65eebc705cee67ea0053ff37cee871a81959f33d6dffcdd08849bdc9afbb1cf152;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ef8f8572c78cec3cd6fbda0bb75f901aa418f2ba99716a65502dcbdaafd133c7884d9cf04f1dbf828c0755ac73811bf10af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h375e4ce9e1a26d9d045ef6db2ef95b5db62b86142ee996ba0d1528f319eb3d285d17ee9c37b1619ea5efdff338f9f51950f6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4518fbc51f9b176233ffb9494232a23454f78f20fdeaf690d2a0744fc350b3ac93a1250c3457ca3fcd8ca6cbe20a92e5f7f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb173c059d556f9f31ebe24c3ad37de0ec8abfbbf91120610e4ae9175369f62fc64940243611e52154a2775007aa16992d8c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h312aad0da640a13ea277f8b4b5195f4231d3ddc326690aa1b7311eae8236b5254a70213a8a61b83cdc4eb016b2eb0f9f7ea4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3c6315f7c51751daa99745f5ac951a6ab984bd833a9c66d854d9ba176b566f3b12bfa7c56951a15eb8531a0a22c95bd116fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45c2d3e8d16c7cfdc03c7ad442c4be2e9cfeba8a4773851147411105bc9d80d6df008da706ab06e16300963dcc6c89bdf820;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb04f626c3c234266b59213140520de815b2399f6efd5f612cc7e023521b5adf92b2c26e2b85d5240bb99822f3a8efe70ac1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea58629c5a7e4f4d859be060936f8ab4f86a18a5e1c41ed025a28ce706a252271cf1345dd88d3f59d05dd64cb19650d83962;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcfe12da37193cf06336a640da6abb5160b75ec5a5005478a093ed76569f32b48bc0e77ec25eaa4567af6809839009589781e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h71e187ce3a16556eee9045c28da4e18df72387a5e45526cad402abffc4ff01d0ed99461faf07b5117fe5e278562c8faa44a2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3008938ba03e1b7daa039d4aad2055ff6c4eb746fd98a5beb834f099ada72fae894bbc51672e9e95bc927f552ba78eed07a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff59316aef2b6386ad4f8b4e8ec56efb51fd82d2507cb9d960d79bd94c5609820b8f29905f36de04227121a890fdfae1e1ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a0cb2fd08429200551ebc724eaa7bf1d82ec879472fc44985a01cc55cefb0073c542aaca9f26eeaa35f1e29b4932a9a9e60;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5da5649cbf7de195c15ea2f3c6933e755a0ec1d9823d17b4b511cace59f65969b3f65b5abc7ee8b1b867f42976dad194654;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8058b029e49639ea6aadea4545cf403bce6abc2149e3496d7c3ad58029dfe1bb205be643bfdc5514281e5a6b7d3fe9cee34c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d474cf2a3108e809171260e9bc9a58c06bb38ba9b2ea46361b0c5a472871c5f828e6f372218d78d949ea87470ac7a1bdce5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd88695eaa22f3a5b93d8aad5e6d41284d57a4352e07bcda84bfa5d0a9da6ce4c40036cbab68b97bb1d7fee78965a1f8805d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h300ea731624d06b8a77c234f7164b5b8e59054c21d4fedc99ebb0d1d925de91951be1b39e51abaf3de343b8060eade5c9fe6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h19e9bf7668ee9a014e9e185b9445846833cceeeaab8ab1e280793989fa1293d3461f1b3d6144f84737fc15b5da4e5e2b30;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59a666be69b8885b397c2a16f62117981c566978188a6543a01bd607c3cb270f4f693f1b11218cd555953d0973e4b6891965;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf0bc2765a7bd063fa788fe829c779e55985328c266fad2fedd63c64a309205dde79923b133a2c0849a259a24e4720921198;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22be33f66ed4dc4c4ee07ab2f86aa34a88a8a5487305efb9f9ed5d905126cfd25388fb0818113b964417eb8444437733f627;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32a53c6f7519d52458d336054a1573c3a0f6a2c1760457d743aa3485a5651fc9b96e624248cca8f0bf4d17fef0313b9dce00;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89b36c6a9bcf452c2367520b4c874ff989dd7b6da96f263394f0f6a6dd22fac6b30728ff6bf9ad3e30074b1523032bb37397;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9403e3595962d8cbf34b759b78f6d7a8f0d671d89aadbf587d16b9c9b77d904af315a1178af1a3b1f8cc3ab2693108e89295;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbbf0f5009d76619b3967a2ab507885992ac870f8ca7c26b28e4c8345fa4b742f0ed57a193bae60e8fde34530da09b8322788;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49741f1a05d44b705d2ece29140b6ab0481279b8c355bde26517c0dfc3d04a476662f4802db27300f1c066861ae62e8601a5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfac0adddb44c04f923d011bf011f62acdadb23f40c06284f8aab3b833ee43354ef963c613b06faf8274923caad8b9d223651;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26cd01cef14120dcfa47d73eacfb5d1545fbc25688f9cedcae23de277709a9ecec9cfb61a59c6401511b84768fe904c85a6f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9cd169159dc9c185e7e1b6d3c549f9165be4d9696783a854a4e5ef722357320ab6a96899de6cdf51ca9562da67af96addad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a8d6639da5b9121b15e2a48214690b6f602dd1bb112aa0d154998efa691417f47d7c419c4ef369218d8edab3c12eb6a190d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a1cb426eaeb9a5eac37b9aa1ac10fdf041a8234814e99f491598c04fce90370063233380356d24fd3a60cf8ce98f17980fe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he408344b62f0f14671d1f46f1d7846e928f59c5e43ba28d0c368763d1412748981edc86804824f2291a5c274eb2a02c6ddd1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e64640f5dde5637d7de65785fb0956e4ad580d92a94050f39bcb02ab52c93b8cf25aff2a524e0fd37a4cb67ada774c7941c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b4ea91515c0057ee195a35674d44607fe706b08230015f56b8ca370feeb6ef726a6c5d319e7c2a0e3becb68e0caee8e3ec6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h631214779502de108075e70c20f8ab119d1017a9c27ac06a7b943ccebdd7c457c407398b6e2631b4d4ac3408feaca97d39f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5a3344f9cfdfdbb50e285d413d0eaa11cfe520d1d94d492bc466efbe3e66bac1356940afba68ce585372f8660ebcab8be99;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec0c6a2b9e78f847189e168fb22396cbddc5db272da024f0b73cc49832420c6088d41594180dc6d464487a1f6f19a01f3291;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6be5db59819d605f2528fa8a9211ae38598b7d84d8b5d075109e5768b5f54f4186f8f693e1dfef28e4f3fa59e5c5b605621b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h964e65ad2b11a069bf32114ab410dd45aae22bb1e886e9b8decc76f9254fe6fb1b9354d35dab7fe8d8ae2418324bca41280d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ae9c347cf7ddfca2c8b750ff0588d8dc9989deaeb1cb1ff2c53952f2928d011824be651423c37e842cbca36cc970612f68e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12e3297638f47fbbe24856a6520cdc9d32454cf909725e9b6fce1306abe1c24e8c1ba49765036ae90ecd6eb5945615c39b16;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88bdb4a192322bef894611dfc1f56d6cf4bf63b8aa6c9d63e5bcc5ef855c8a8294fa5e4a103db4e1aec7897436f4658a0de1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h41ab08279b3c8406e8bb991d636e2dbe791ca44a3ef9be491e7495c5a4893debd88d408430a41a9eaff96a3d606a12ed113f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4ae035d6b4b71312017a7b67de9896bcd8560b9716e8efef76df5d8512731730999b39dc8ad6fddd508acadc2d1eb2bb26d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hacf58fc26af14bed4a9abd8b655203955c109df3bea25cd4d1554d4c4ee0561b8651315cbde8d5cbff2291cbf9fb6dd92145;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5b4c2990a0cc8c62e6c3d014e6e198e40fe3a49b83772554f64862d46693cdff80f757dc3cc1745810b404fe368ad40dee0d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb1b429272bc1f66cbcbabd0c9eddb33e868e10d7428503015fc167e8aedae661da14850ed08a89fd7a9e0c65bf890c73c16a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h294f198290142d5ad2e37f5f6ecd787cb4027658a9d160454d788360de9beafd89cd86af9065f56f4965ca5010fb6beb5f7a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9842cd0414dd18328a70accb97706c2f5398068f4304d171b6646d2d58a2dcb3807fe0ace6d37b67aef0c7e6d077e6873519;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef9945cdccfd34a3ec3bc05559ba7852828ad80a55ae5f50275a162a4b02ed34d86525b73b3221033fcfb67a34804651c910;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h74028e74c9a126f7ed285c50432f1e721db0fedd87db5ba3db791f331d269c0beb3e373e6b8f9f8efe6849f0e0c2dc799fc6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h785f34f11222bdd2dbd6f1d1383e91167292015f68731338cc7ab964b1f2c69ea0ffce66e9da534e58bc3731d5b0faabd252;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9526869760b0aaeaeb20e30bafa1a85d63da71039918eedb0d5248ff6f95f25e937d918498bc409833971944afe2374e5066;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58170b163f341f7b792b8bcedd1136a15e1127b9dcf16ef4fd3ba59541cc4e2020d5b903125350fb3da662641a266e7975c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7611332ce989c3726a7ea336ecb9400dfab2cfb92c53d5acf813cf0f13ecdfb04db23a033491ffd984bf2f45e3e384ca6562;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h108bd8951699010eea120a95dd8f98504ee0df22e4376e3717c97cdc36943c969082b768d6120347688cd7e75a7f5cd4c6fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7764cdce27dee7bfed63fa0fe0251e28a6fee015480e7fc743c56fad4e4a35b9db089e516d713f444248eb0d1e6bcadafc7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8fd8c14569e0debae11563a58ff90803cf82e56d235ca86d046797be98ca8bcb49dd9b76ef5dd1fea533b1f0b126da59412;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef1220ab6c98929359493b481dc184caf5ccae61d64572c66f7c48d8e14caf3c1dec2c6fe64d12f9aa8541f69cd02a58ca6b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ac1876b044e67f70772ad63fe6e7f4da10dfa2e79586a95805ad26e9e93cfcb92fde23fcf907395b944fc4d94f0d1ca60e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2159086c4a76a89cdff6c9225bd21d096c94d70ca3937c54b9cd635068fd5d0678b365077681b6d79142a8403dca584e60e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3752f9d58f749c3a8fb4fdbdf20d413c7f057e11c20913a1666299aaf6eafa5aa1cd57adcc8d0868301506990393ae2be11;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcae2ce7a4b3c10614800e384f652efbb5ec21bba9eb4ac02f807ad00295bd210afd10491cf336d5ae2702977bac8c11debaa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h419661e150c33d2fc49c8a29a7ee7aedf1a22675cce110a6cad660b0f243825e6e71308bd4b1f65f152a0582f8764a0c12a2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he3759db251cd0e116a7d74a5bd4addc420af82515db20b501dcf88e34921dac7857c82a4babbe62c430cb9176e6a76acc6d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8672242340282a03e3545f27b6731ccea99ee59148e7e1fa37947134d484132e77e41b478187c575d0d75924c7dd5d9fd1e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2530dd81d9701f7e1f32f35e470a58bb513f167113916e7880335562d76b3fa1ab40addc9dfeb0acd11464b15699873d00c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e7113a7cfde95700c06afe3fa16365b2b0059f453b982ee4d3ab34799092fb751b52c825f3b73ef299aee0161e27da39c5e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58998b6e9fac95c115ab946e47683126d178065471c67a0577d80a4e119c66c7b935afea79fd320b7227f50eb6546d35a454;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h235796a89b529e43d21f77cf72374058d801f0cbca78ca12e87ec16865c466eec3f8437d529c0ed5103b02a74ac6e81b691f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbce3895b4b0e3f8aa44d7119e4d5be3df9ea2f46c63aa239c259c29e74cb45c06df0b055cef010d94bbf0ed557a32f2195c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70a35fc3c2d21b4b4a014b3d8d2ea38303b4dc08999573f6487bfd01ca0e6ae89e8b0344bcb100652e6a3caa076162f19919;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce1f714a69aae2a8a3754524d53e6fb7b5534b6c5054bd1ad6b5ed98378021ffe476349c34ae3db4d32095395046f02069d9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h635bf676df64200b8fd9529a24c5a903a9d00586289f2f8e67abae3c618e8d15c978c3f01d36542a104e975eb4c5fca32fb5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36448d0d0853a6ef267fb1e86cda272e1804eec8d8ba2304450662bbf31373289dc65615216cde7e579424e7bfea6e9edabf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23bb5ff0835c9ff1e5e54276644ce666fed52d642aacf56a14edf6177e88e8139059f039935cae127346d3b19142e6fd7145;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7feb5ed4fd633df214b162692f9c23526292fdc4b360f0c2c296ea13f5586e246da2417866226f18a3f60b8d2fbecf409744;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14d9d23b9a1dc434105941fd2c3db7122fb1c95dcc1a29b3cceeb27416278127ff9bdd5acddfd44e86bd13120e64b180654;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1054bd7d1453478598157683ffbc892c80c9a80c9d5c09074c13eb037d3f5145ed27feceb67c370b27fa170c25f4154eb32d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h520a4c3e650291baf772f99ecaca1835c5499c33c89b2b5b8aa816763685aef54fb14df8da9b90c8627fc980be0972742b83;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed69b9c97c8de5d75630de29b211c7637f284c30b09e16c2077e72c2e3d9e23beab956a845d5d87b21573970efb62730832c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ae8ae06ca25284571e96a968116700e12762d559bc1ea0635562236879591dfaad870e133df19fd0e74863c968b2dfaf7e7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffd8240c8ae9a3f3e0e0093cff1d58046c7f43d9adb5d5c7323b48705b71608b014467b07fd515b378535ef6c1ae90b09e3a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h37b862d638833dc8e669c234450c50d10663077f6b3faedade91b4aab984a07a96f63414598403bbe82095b8f2d9a80900f6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9af307307d387ab1f79f13730d9cb63878408ee18e01e52917556a6414e3113c6303b345773bd6bdc2d4e7fe3353ee08515;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7af9174f265e6d5972ff63d40104de9d45fe6dce945a1075d2ce2e1f52c5e0b80b4afc17800e39ef8405bdbc49bf0619f56c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64cdcf600e1db09ce9160033a6e30ead350028c55260ec16f3c8582c9bee4e8a71afd28edb264fbbbc44df1668b8cba73633;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf54cebe965beaab59d73e1791a92336246fb0ea74e234cc7362cedebca6fa350ac209194ad05105fb726bbc22a0790307a94;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbd5869d0f9ee2e59e73b3ed880107dfff05df1808d7c6376fdb83507e0c56d397d1433d602b580a38f8f05cb5e7bac8165da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ba45caea5da98c0aa4553fe4ad239f1dfe4472a145374492c25b8e0e70061b1e03e572593becb84c1e566b96078418076a0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h271d9dc3c14ed30d0c2d74e836f9bc08bbea5940cdf1ece200a27a5b2f7850d649c5acc53555fb585ff8d6deb23aab15c816;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8299729a79da74e8d402348c99964e354d3e0de493740d635d6005285a781544f170894c1b886ab943fa2f8bf6db0e933a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a0393376e513df7f81a036e2f7ca008fdcf8c58b00c37d31087186c31b59cebfa83ffba67b22ef4875cc1430ee57de2256f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8a91812cb39debe9f41b0fd16eed3ed545e6472bc99f1db6aa9f3f93a69517a8b2efb71e52ed5195740948fc114c91bf09d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62fcd856f01e594620e248ea0696ed8342d9c66850e6bdd25662c4213324dd331a4a5721b1b1b02e0addd66bad14171cd87c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a0ccb07a9b24c43bc06d800fec16ad4283380ff7037167e5fcac0873c5417df1c2d2eded15d4acf3677691e1da1435c55ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc23bab08bf5183fa3104e2a65f80e52d821beb51ca4a22eea3cebce08f6ab363bfcd819325d773428719bc08eadcaaa08fca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h27b26a72dcac47637580cc0d733d9d1ab9b7856a229638416ebdd8bad80ab2be2a5cf3c932ca319797f1f4f3ec135465378a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66055f8f9613f369e799eaa10fbeaff7900f609e59015f55b4e623c0096511571d83ff88ddcf427e08825702bae8d7a50495;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h836f0f6601e0a794064e277beb806f1004231c015e966a643e54dddd04d892c29005b7b54b12c5f5c0190995e0103dc2b6cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e4515dea2c1c8551babf91830bd03c33fd788fc4f3339b9e43989648bfb4128cc4a0b10e8502b76a09d38f4ae08f706e8db;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68400da3cee40ddb66bad67bfaefbff656a499c168444ed640dd0ede0e20563d929878e362f5dc5d4570a07f3656220aa0c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc0d3bad5f6fa0b146375410816d828b2a8bb5b9b54db41dc3af87a6748c7b2620bd3634aee337844b382c1f7f575617091a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hac4ac69ff38864baac51cbb033f75f9878799edc6b49f88e3d58b7a72c02447d3e6404a7554467f39e11941f3caa9c722fdd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6649a62d762c255271a16318733dbef94ef62dc03f5c1eceddc7690c9054cc280578560f8af60ffdcc4176d3b448e400632e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e053ad48a0aa2fb2e29c866aeb1d05be9e191f4efba74677ed9ffd0353009feb7b09a4e5ad7de54f968c36c79dfa82ead09;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb139eca39a7e95cc7d730a453e6e19bac00172f164157e3d6c5459d388ffa92f6a8d83d4905a8b68b49590905edd3556cba2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hedc4876bd3b7ac33e214f580823bc8b0cba62f0af373eb61ad15b59a81cf78db4d7ba806e0d0262ffc2bbe526f824f665a8a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99398739817302586b5eeede5e91b53a60a27bfa60435f108a7fcff63f78ed46924f01d6190b734b72a80d99c1f2375f15df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84223537586f033d1054968bdb8392645a89ce64a9d624b1317c5f741948db8932b754f173135dd659dc6d18be0f955b8913;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h394ec5ad2bc9a45bc68feb5709303266db8a35c274938cfaf2fd4da439c53eb074bee1e3ef894f41f6a17ce0a386b74845fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ba9cd2683470afe777620b022fcddf17d03a9c4ded13e315941d5704afd87fdde3b4b561ee7bf5593852ea3256226c9a73;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc6531cf49507d7b90653589175c5d031ab0a3506fc981dcaa7c179dc642413ddefb0f6e7c874da4988cc5c88a002bfb9b131;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h121fe2fe22d0b225dc7e758ecf140ebf1e4dae90ee6c3a1fcf0929f0afd2de6f5a43efe000afe9b148cb5e5bbb977c493704;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbd060bbb3704b850138f34b5c4605bf11574d0d66da229cc6697884417e76775dbc799ec1d6042cabc6f3d056c585888e04;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heda048defd6385ad53848cfa6a2f98e3c3fdf2d182976c0eff992ec34a8b44f238046ac58409f85dfa2ae54a59147a56c60a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59ed8b43d94f6372318cfecca4be5e1727ec348cf411b888ee6e684222f6e12cb871d2d85f32ae5d78abd1c893c8c0045aaa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26356b4c39e6272f0640ae752045038ec762e740f0c2f17c56d1d75121195be377a8eaa9ecfe4c7872f07cb6d94d1e2ed5b2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0986546d371071d9d5102d79a01a56c10ce33a3bb433bce62548d5ed62768f05042efe604635fa376916e05ba8b15d6628a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdde56238ded55ca04d166f217c0e05c41e4626938647c1c1d3e2797ac7ba340ef979ea29ecf2d039ae1faf09ac074d75ff2d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7584e14af082164074637fcf39cd67caa081431fa54d9b7a0a29e1bf8d247632680deb63b94711ef822bd0831491b3c65b6b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb84dc406653cc2bd5e4523567b396d1f9ff8d9eecdb0b435df7b75f879fda7b5bf3241fb6c5a3df4638065b0f17ffd7da8d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6790c4845b79e7496ece8a5869b7181499960947bac9dd11b09b134bdb5187073e4cdf6b16d1c8bc94f408c9ab35ea24e9ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3cef322d58f420cc7f559955106cb56712633f15d5e4900cb14f6664dd8d1eaba9aaf2fead3528e4c4123ceb6bf9627d7435;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35e23ea2a338077e0623279ca185d059299b512a2e558dfbe3cf83bcfe5d2b5ea688f1513db96638ffb97184795701e3d476;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9f5ad27d68e080e30eb31f3f5947804777b89527f907019f2a1837b8b0a443a81778b9b68d3a36e05afc87b107ece58bd69;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb13880d3dfd6de30514ed10a280a2d5fad49f8fd37ed885ffe65ea1d65707e9a8719cf7b1092484a5bed5bb3c8d4ffac4478;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h243a658be74f6376e8a5b82feaae4fc4a28a750ad56189481c538e5338e77e8d15f4385440ecec040882dea858c64f39c74f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b2ee7df7502423a559a233657a107dd015a27374d4460968d89f0522280001b3fefe0947411d867df1f0609a37427422941;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf88747b95b1a0aad6b96af46b1467be56aeb69fb7390063e2cd126a891aa03d64aaa1fd6eebe427811b475c5de5fc1add277;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha102e447631897d0ce6c5a71a78c8e210079ee42d493592658aa401d11bea04f9eb9f5e885ce6546da29fd8e46f735f305ae;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5696110f18406327292ff6f3efcc8cd52428ad5198007375f7935ea04fdb4348bdfaef06ab33e3c998a66b495bc2e3cfe28;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he17784571d7bf897e41e3185f1b32f9667b2a494151b6cc05768b0b628259127c6aa4e30e3ece52684f4f2a07611ec16662b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h386196e6da468b837865407ffd33218d1554a732abfe8b7a57d758d4962fb882e2110042d1e1fd051d6d5bf1ea0eb91f47ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc116ef345c76b96fc86dc5fab88f953b88119866646c24f9b0661987c22656984eab7774a833770d1fc66944cb6f1933af2c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1778ea13984b82a6c3c98318d6cd9974069c9b0dfaf282b756eb5e1ddc860b700266a92145171d4c9d5306504f05e59e4ed5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb2285d8f8d97d3ccc65d78ee94fa3b5787ffc44fccc3c3e960697063741bb004234c3c01d1434e357b5cb28288fc1f642cb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66681732f5e5a0806451dce3f166d7a51cd23a9a32211e9da6259ac2274032aeabef1001e7f9f9d4584c74c1878a67f6d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5457e769500c99c627100ff4f76c88da2ab2e771caaf47ab25c176d3c4284f81b37debc920a0a85733b2bc12a3cc684ab9b3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbc9237f9fb37de417099eb290ecee2cdb5e7a1ece3b416b10e6174c152a1a22c3f24770f601041f7880b36d2d337f0af4e8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6590edf8ccd9494a0c8fe8cf3b94caf65d37f3b0c5c0f6932d531152ad0ff4fd7e2155eb6bc8874317e6de722f3fdbf42231;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf67953b2b5ea2891ebfa2a5768c0a6e358dd5d5bdc1b922143d5d2cd2aa4f6a1fd433ac6ed164ed5a13c54735d37c500d23;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc067615dd087269df50c5aa6b9179d96c4d5f4ff421a703d2a2154aa9ff507c35efc815815c751c59b31fbfd43f44df1b4a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff40133ab6c669e7f4298550f96659855bc6410abd15d7e20d361518836657ba779acc5db6caab382bf9b25ee51e72805233;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd00a6568d2b94d6a1688fa6bb5b3376e414c4f638cdb4fcce46d8d8d3de4e0bb748366fb3ff920af66fc22f172d271866324;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h348a14249400243bb6dd0ddb40aac6ba159eb797cdb8321581a0a6105f682af77777009df8e793fb88f8d1b9d8e22df3a13;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7695ae17d172459063ee8bf5b75a0d555a045c585441f567b3dd6c4d1fdea4545d886824b12bcf8b662bda51ff90273343de;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1fcce233f32491e115676d5ec74d1eaee6b5b1b6f3c50ca0c5077bee275e1f1ec11017711f725b9912323cc8401be6f9aac7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa672998abf0a8ad39c3baf77e47b6a95bf9187e684980e5187566a2c26920834abd6628d4f1527e111ca8c0e6843bc92ae8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he91d9af8eeb260c2e87d1d49976680f79c29dbe321cce958b3e007cdce910e39554a6a4b0cdd8fbdcf379f12631d9195d095;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3ff0282469ee743a2c583ce90f76ae7084529275f3b8f9be126cec6321336d0836a7c12b0ddc492418bdc22ce3c2b0b0fab0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64cdcbf518c88266e7b4678e472a99e2729e10fbbc0debe72b49bd006df6b745afd51c7cb8f73a85875cedce1f43b99a8b33;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f10dfe42947d84cc9c9097e1b9ad53d86ebc1ec87e26d8edfc45c89cb48e285d41e08285cbd142e8e4e7a7dd2b4f254ab8c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb605b62a46c49a03c7001415e4370863fea4b2ccfbbd9f1624e9e87abae551bcb6a02791443ad0a3eb75103737a49ed5aade;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4d5a0ffea2c308dd98ccaf6bbce8bd21aa8db76773ca9ae9152e1881e456d15aa26e5ef649060044e31f10e7109f20da1e9e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4167c1244ae676e50512951963564cacf2ad9b2bc335b734292e758102c25b17171b8e2feee74880a2d6a0ad60abd26542b0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b18ca1cc29acd04fce679acd2c3591ce07123099d99f010d4127be9a68fa243b6838e7b8a9e0a177cebacab146a44bf6e98;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc67146aa480773e542542920c938c8f57e62b6f1095558789d59e70d4b9ec2f65303312bbb665b63525367bedde23a54309c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7954f61e3738fbdd99f18266887c583e851257a490e739cd7be1e3be8aae9a33546ef0213cfa19139e90423ac30a742e793c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb86aa6989a07d9d9e70581e6f7eb33396a7f9e1e60b572072ea74c83e4138e19186d2832d3d2019933a52c9697f913b61966;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hade0560435d1d1b0ef5f7f2760a499c68cb7684c82957a63c005dcb38f175a614f502d2db15e1d6b769f7474391f5fc21774;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9cb7aac62667c9b58a05c01428709c904b0ca7d0904368dec1b6850d7aa5df6e657ddf4eff66261e645cf11df20084ae42f4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83fe5c567cc4b8406ac905ff99b7a09124569d37ec55ca0290d72d75fda86a30327ffad88ae7b23ca7405221b1c773b9d559;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcca84efac75734ca29d7f349449eba10a35cb4ca81437c0ec3b71c8d3b505b8528fa5573beb1d2f76fc41f9846ed268a7716;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e03f34669e2291e885dad850d2aa0356042eda6dfc4b106bf90a6fc9ced2080249aa44bcc50b710e71845601e1180189c2d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6eee69fe31824ef72020d02179cc910bc43f947f10983c02823205a5892836eb6df3f8389ac8815944836942b7df02e1a65f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1101b82b386c47b73743cc0c7bcd953a77ec158f950567624d9a2df72de9c81687d85d6ed4701d69c1b7675705748bbc7819;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95f541786a33e2b43b62717ea73967d71412f41776519266c858d906a8a5b2ded32cdf61a1980beaec8ffbc5ee3e39778fc2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51ec99c95b6e690c25c1cbe682cafa8dd9c2b4bcefa5415cc4cc819fe5d801b1bbffe5cb0bdbdbd24a47ff7fcc7556d4d937;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ead1d06fdf24d0bef8bad7ba769ff215a98783a42dc1ca5e7ae0dfe40f295823f80e0cee487f8ad7cdb31379a560b1f3880;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0663c07644b788694a10116a23c6b4e168a57d3e5b6a8d1965cef98309fbccf822ed6ca6eb828fb903da5e779f5123a669e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h824b608d74f780e68aeda029e02611dda28edab6e7da6e8e8303780c1f3426c38080accf7dddd00ba7b60c50f89c09fbb0c5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80955afad9b46e0d6a748c95745cf3ead7aca607b694f6cbd76e95e8f712a2b1c182ad884fa43646457f4e6d477f08f9c0b1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52764f29be0546316325b32cb4821ef2b9f10d066b4485616a99c544c15f06c0c00b2391208645b233dcaa64939cc1c5ca8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef02b280ee7defc8ff28183bc68b7863b0f4d9af0923b934b07f774d19b180e1d914f6c7f26b6ffa500a89c4c31d2f555f68;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56c0e6ca873e2630bd5a287a1407dfcf87302fde272053b2f57a20e17d928dbdea89206409092067d8871094f712bcc925eb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf68c70bdf7a00bcb1bba737c3511a93cb6c9d55b37be0671e9dcfe9aabc7cc16761652adada4ef0f606000cd7022dfed756b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0b8791c6ff46170f5c109955becb4002358dee8af3a3fb8aedd8caf677d641219a52f44ff6058d141e1eb5b10bae9574465;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he38c4047cff00c4110984bc281babd1d7d4d96db244b5613e13811108cb5b0b6f4c1db5d8c5971ecea2c32dc927fa2ad2edc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc91365e6b56dde186259899fc5f11ef655ad90d86237475c698a2d23a3cb8c30e53dad1178f253a87cd4a4092a6a3a7405bb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c00def19257dfd967088583e21cfc1cf49270eee4a3d3922d71edf4e5c37b0542e799e404c20c539b702057d3198bfbf5f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h924f3a9baa9a935d9bfcb07ce076cf9103f603c67215ce186560f71f1abb7b05ebe0398b93cf69037b02d64ec09b040175ff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d1037ab7d1c82cbf632865119eb9b38b0106f6ffb827dc0f66218bd6a626102bbbf16a0132c22c5416abd0d6e5327e389fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b77dedaecd8fcf8dce8516a0cf6c72b8a0a35867aebd8b4422c1832f2254c4619a66eafe52aef651d9ed757841c689f8524;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4adf00215a4eadd603cf33db9e144e7d698cef706aa2657a140fc40dd9653a7cda64b89c0fd16877e449f857653faf979f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he81127f989373592353a77d10e93e77d16726879e7810e7b4e6bc53104b13d61ede68211eaa3b8b95f38fbb8a859a768080c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2695ddc07e76b3a1d424bf19c0fd7d95771ee83fd23dedf60a52630b08bd86cf0202ad93c8c6341879e2e12e36536f8d2725;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc70b37e135129acb0e8ada7cb31abef7582b231c3ffad28991443773500a793a3bc2c621d574d8009c7a30e11266cfd388fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92ac88b8ee3b31e72c27baeb1061b91f55c837e7cc6deeef04e0908b1d5d64cf0d471d7d2458be41f2b55c9b053a2686185d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f031fa9df069a473d76d50121bc94100008503ceee0b1c72450964c82068eb74065bb2769f9d131ceb6ac0b8062edd8e700;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd13049d2cca3daacb9c034d402275b13faf0fd2a1c6ba58e986696c2d63638cbe9c9d420758afd55e54688b02098ff32bc3a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6564b568907c11d57a472bd206902b30dc0fbc934c7a09b5fa12eb33b6dd54c26ca7d8646e021950924e3b49b1a7379def61;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h324a003123776cc10df98777edfc9dc926548321f20ac2cb4f02b47e2acd84fc8d0ad899b47af47c68eb28139b6e8de5e519;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7be73c472d0ee64a219edbc5d339fd80a01e0362177de3b0df61607b3132aaa7a4094e4d3405542399d857cd4d1ad01d852a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h625cb5e89095026fd4a46ed1df1e4781372f263501c1d9e677dbe83dab5f442af77f4559b7b1d997e4d312ad9e3dff22cf4c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h765675168b4d3f2dadcd52f5664fa0c21e78dfab2a1e417a16599220ec33efb995703cfe2fd55e060d1468dda008c918e447;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ed934e81a30270842deae085a80724f51f0adc619831996e1a00768b8bcdc541cd44478d5677c4215f7eaf6d53886115fa2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h51d514aff0bce54b768d5532e77744211b4c6ec8e1e94352d83e3784acb78196fec20be4cd60b9a3515f8ce626fbc887a02a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h847f30476a2939eec076f2d7d5acbe322654542dab3a32958cf4d18acd3478cc6bbce2cef5760549945c2ad703875575779d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hed7b04669f672d2e06b2bb026a87574a8e0a0e07540623d5fb3362c851b7ba3c6441b2b97b7cd34397f78cf74ccbfd3b98bf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h896a24666256565161fc9683b5a73b013890b9c383af8a75b8852d197d26911e89af996f5c115e04f3819f55d0da0dfb796;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78337f44a0e0059d065da14310ae0c40a8e1fca3b3aadae5f372dec5abe50cc46af8e2d580340ec0058449850870a4f35996;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf94b02b24c7a23f4b2551acbe49282eb2c8ebe0c5766b24b1b9192e4666f31274125b48e577cdb8e7f586d5b2c64455a045;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a4796d26dd406f3dc16ca346a3447b6de3fa7b589455a71a4f10506687bafa0f92dd9027ff88925407b5ab559e00d76d3ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc55ab06acb8f485ffc9dc33367cae04d22344ff4c59f8053313c5b0a0401a7659c50b10c469565cc346fa20262cc70faa71d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73e8824f2b99ec5381938d8ab556933e0b5b5539968335e94cb52f1622e8ce568e1b9655a4e5fa4e34d15675ea761924407c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6259775733d619c219868a49e280ecd3c1ccf8f97c5b08adf20182728f030426b1710c0bfae95bd7feb1cf05c772744c1118;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6137918d6ed6c62c92feebf058e02054fc35239a73fdd22959cad6c802ce9689626bf538eb35263e610b27287552bfff0c1d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h176fb7252f3e1aaf7649025711b606f864c3f04aebb65f1ece0854687f6a411a226f26b69aad47512f3ca628dec583599c16;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc542740ba979318723ace962a0ecb2a114d2a37bcfd5ed45b17094e514f62108dc29ed990a22043c384da59cb9ae4865365c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h91d178d1aacf155bacc68c685010bda6ca65ab3419c178bfa629ee63b8ba7ad27b87d28aae4e16186dd3233c623289dd7762;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef8b078c544ac8be1677dec24abeaf6a8e37977d554b1ed843d317b4458a831e19bb165e112b7a7e43ddbf588cdc98c0f5e5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha96fa04e7ea9e6693206efe198bb12235bbe0d36b970ac231f92eca7f62a1b93eeff97a7aee55014af60f6380f49d0ca6441;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87e8c61f5e79ae772c2e3cca92b90207008479b402a65ca476642b247658e89ff1297f5368d3bda36ad246f86880a2d08fc3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb35b872db7326634125563812220b920e8158cc44fc2086ed5201f10808b896181b1503ffecbe819e20a566129ab1c67aae2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he532c271d644be4bc83bdff39b62a7dfaefb378cff9651795c0d416e2f58a4f7c20f36af75cc55a2f462e25b874721d865b2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d0943fb9590f3566c0f738c7901285c7da17ce81803926be357e69138f08178ec154e54756819aa1bfc8b8043dceef50e6b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0976d1c4a9c2478d6b0c0e6cd401e777a865f587ef67a601684aeb103ed084809e0b73d3e47022b14202eadb17804a95709;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h87698a2e6911f4d8a69df57d25c43ed1f37fa990de86e6ac68ba6de3fa0980e655a7f879e0efe73efcc201e332ff09a345f9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4faf9bee151e829da388de7a996701b543f8c39231097795a99f6db78562dc36dfed792dc10a786cdc69a7becae04dfbf7d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h222ca1386c6c7a24cf75312c9ba14ffaf94fcd0c9ec8525ad6581baae738902f62e2ee18cca37f65c90f4be7306edfcf479d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf850077f2bcf619f08493ad1d38145a65a2542ee566de3b4e2fe1b23ef03beb59c30e7a8f751b2108fe8f3a11ce4abead7a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had3f6d70723e9420e9317a81ae78d983b90fb451d68d4256f78dcbaca271bb7ce4cda84ebabc7793a15dc3b27e48523f4679;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdbf015f3e132bde4d25547191c7a66fb159d55c8f479585bb5e7b5905538f5ceef5901f4f501e64d8ced0334dd8b2e3232d1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha885014c3cfe9cc21a95cd3b6c4d434db0de7d13284f8d78ab5c7a3b7b4ca5e865104022f89a36b5ba49076b7dfaff3d2496;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5d7bccb285441754464b8f5a4755e40760eb7dfd34d6e4deaf398515f51fb8aad3018b3be2e55650c155a3e0289a3473643;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hddf037e12df53be59df65cf306d00ff7b24662cd238c6228b9da87f6b1279e51ad651320bfc23b862f98378dabab7b8cde8b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h450528c2de5b04cbd620c5037e11625237a201594ac39b9805350d1abde0b53ca1dbb702b18389b9a851213e40fe71402d8d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h24552b85a54436a0c327007c43a1a79cc4178f0fc78c15350c4fb25ed276eda5369ce96aa1ff635c2c638f4ddc3a3d9267fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde842466e12394d45feca33c8cf663de3b7482fa1140ac9a7655a35e7f0378357dc908553267c93172cd5e809dd7e18ce819;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a678fc0ba5421dcbc8d8b00aca74869f62f97d8666cdaab2f875a285c07d45d6894f901a071a9c5bd704413a83bba096266;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d95a1ad85b627249f8408b3ae33b5c6192b4a9f560e3648e59708d0f735f867b16e00762711df3c47ed37b778f84e4644c9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd52f6f5f0550e8b58fe42b622b4b3ececdb7e559cebed76514a9a259d5fc7492df7af5dd9fb3a88d46a35992c4e7dc30dd9b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9dc758b7b9da99660192d604176f1942f09c9bf4c44bb0d1c39dcf3c5a5a890b0a6992b2f38f5dbab97505b99ee3b5507226;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7170d2cb28280803094db47a0100d42876d438a37c39074d736b4b002f7fc50f6c2db6c465f70682df16667ee8529ce9c818;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb86b265d5a018663c970240dfa97fb82b998b7f246193f9123b00af1c3c9d39e9dbb36aa8b9322dcd844bbd269e125d9877;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6851fcbdfa4f12a53233f3defda525e6127b8d28b456858461d3a5e7889cc2ce28625e5c54728e914babb7bf7cf81b0a881b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc694932c743255206f0499eb0ba495a47e4088d7d60c5020478c4e6fed7f1d14f75c4e6178408ee55a2103d6840750365d04;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb02a7f6a4549291dbb35a9eb068bb482da9b893328e23447d1a0e4cb99c3339f567759af45205fee48e6466e3526ba88a92;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b529a38b57b5bbb5d052002a91e9a051df7ced91dcf7670dbb6cb9eb382b844edf6ad62aa7d8ef1b7036956484910b2721f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h142163e7a86be5f205f4acbd1b828fb65682a33f64829d2b3dac2b42e13922ff01ab4cf64b812159af216e026221cc495125;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5a635a34410caf6d2bdde10492622659a1fd023ab1b9a7be11ccee917c05d3057dacdc62906705b400a09a5304bcdb4d2c9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e4ad38d7a0fd95c1a8211bdf1f247d7b12de00c7090a6120558c128f5f6e455579c30a66788e88f00dfff04ad412d6ecdb2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h663b8df1a6f20e2aa14c5b719a95fcb5ca8ad6780bce5310a805d3a02a4b41c341d833fbf86dc42f39693608bb371769259;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h296174c0fbc1470ee996fc6fbe4bb53a30a0f66f6286a7d2f5646f5bf2e325a5095e6b101724d1c5827b9298d2a389de43c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h990c1dba857a78bcf09096509b3212a12e181bf10df1c06e8e6fa946c59d3a08ca3919292a4d2a6a37c77c8594d64691c1be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbdec7d8ad0d4a27e221a815d38d91ac8748bde26a40f31e163f203080839b24ab9906b170df227b2a6eb6ef1c561d0452338;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b8a913c8975f23a9c362e245028289491c842556386344bc2e14eb0cc768fccb877257beb8cca2b5836f0026cf8161978f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca5558798cbc576c07a4215127210869c2222a62a16be01d73bf408a39eb2e83d998d92b0be0e0b570aed60203c3dffcb0f6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4700d3da89faed88307838b42c66ab2df38aabbe32e26baa0a6a16bc29a147be7ea4c80f61a29e3f9e6ff077b04a80077d82;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44783e0e6496f2224587bff03f916fa87d86752ba1d6e9b2b25f7abf6269fb033ec161761c29cf194da0eddb8eb0c9f1a975;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb1f42730a0afa2e6e0f039da871d4c7868679d770a17b7e3cdcabd33ab6acdeda9b087bcf21d0d404c77d9d4f066cd035c9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2fc8ae12b1589711c5cef6f4dcb86d4da0ef994d0198acc26e2d4ef2533806fdeef2ab4abe7d23ef963bb8012ac63e3af91c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8627ebd0d4c4e7377861ab7574c3eddd9c59c70bcb72398607e38c664ceb7bda272658e467d25f3bfd2cb539e1e18f53ca3c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86db9b36b7ae0560e97607d0947a9a29fe9c88a918c5375cc4c120a9636fc288ebe22d0defb0865403b976c384e199c73b0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd113920c83bee863166c24339f0f18c1d946c2b642fb3b60a30613c43b29f897c4381fa45757e8e0897f3498fb99251f96e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4ef9103f4a348058c6f9dbd8dbabc0dae4740a0100271318cde98ad0ba398bbf66c52a26422f7c51715ab61fed98824fa0b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha864b28548c3870b36cf27e2edc7691a574ca81ac1e6e1b9fd79ffc9656f6bb7fdd3c0b7edabf047db888a929f91a19a0974;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfc619e52c13096c2c10be12432026d157a67870c8fab20f7bdb4cea1d3214ed820e4da08b75509190f90a6b969e3920b9be5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h596c95df7289529176074e4dc02215f8b90bcd36cd36ec532945a437bf95a8f1b8e28e40f5a88c2586a245c3d79c35587daf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h102f0fdb231c0b55153d2fd96207e4dc011cc71c512a560541592c40917681ee7b94de2958f040478ee6e4c74b7de86e7adb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha66126f458f3b3114184edb5ba242d5c22c7bd00532566908d446c6e32c86cae1ed0a4e26fd6861ca5569fc91ad473ded265;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc76115cced82e28e88f89813ee9e31cbedba2c6f8af14798c4e2981453c7f456f4e995582f2ddddffa58cb92d7ac8365a0ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcabae5a70bc82c038f550947730f5f35feefb67bf37551cccc3b6b47a7b7b7d87eac3763b969a0f79488030e5fe36e83a1df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ce59c535092fa2c84007b201702a50cc67bb5deee20c59f129e7cbced2e0f539bcbae0356431eaf243da210d03efca2083c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0d05455e1f8351568053aed4a918e406dca52272e0dbb6405e113f2d77d3bdd2f182e8e5b81a3f3fe2c8a5f3205db94d36;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfaeac7fb4b116e77db7dee871c9bd00462dcdad9056e7be929e26836d425a1e9dd492d06685706b176b4f432bc0c52b5a53e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha70a0de464cf7b5c4398319f988bcd4b952a6af4d0ff47bd2f7a02875938f39ea0972115eeb9930ff0e6f418b28e2b5a85f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1796e8eb39bbd889a2994237d6e209f82c50b3199f75640084890945c91a9ec96b218bf3b9d4c8342455fa4a1ab9c00c0f4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f8b8df440b6ae80496e69d7440a006b0ba31c23b8f0ad8bdb511f3f282f23a3b9ef4fa8e11e7db680c92e6b4279d052aa51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h23449fb559fe144bead695419eeea125f2cbc5bd0d17dd586044a93a20203978c4a2bf70483a72e894647d367859c619f528;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5e3400e59e448d1d61a18db1141cc0c30f63f442f0396cfa56601c1dec6d69e5201792ca8fef276d5e078e12e8452a878ccf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hceea94f7e67a4bb07666d766789fdc668762f55ad9482a7fdfdfb6eae2d4f69563a9999b039dbf5d794b7b1e340b1bcc3bf1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd11c3aace45d2acd686b892eebb35687c7fc6229a6b6caa58d700a0474efebab733175f34f8bc7e74fe7040b248af61e77ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he58ec74e0456db6a60086ada91efa90ae16b84fca05e2e77a553d0ecfb2410f1f87e3eb3c2b19d4aba85326508b4344867b8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96e8e7ca76eb7a8575f6b51221d8c5b61eea9cba2c8570a34ca560d8c504bb2bc0f43cf80eb708b58ddc207aeea86105855e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbfc22e40a2d30cbfd994b4e5d368195da2d58dc4901f90a37562d362a10ba331153f52d7c7b9c461c2fd9ae60d86e1dd8d77;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf249b32ef13f5b75dcc22405e76ae95b0f7dda7b3023ba516189e3f22ba120a9959b384d2709a4aa5a3963affb3413418dbd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h68e3eee8677cd5bea2355001232a9997196aa8a0f233c3e6256639e022d507d1003f29d67c9d8729575cf9e5fb9600415b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffe4253d827a75290a2ec3cdc8027a5587be08e955680923171f74061609a3d8d60245089809316da5dfa60a64626e2e5160;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7ae37267396e5047acd48d40297034f8f076be44a3a4b86ea349646aa514a65ed0cd265a5120908976e82cd34d696cb5c755;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h902c2fc4a48b88fda9e41100a30a5492011c7dea877ae431b620edead86eaa91abccc351b1fd8d74b0cdc55b758f96b4fa0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f5486467b9efa0b2d0b59d1ef57fa2f757009d1dfed0a2dd2cbe31120893eb73cee240ff5e9862f79e6e19d7b770390a0d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4ac434f958d5a403d5691facff5800a1218a6802fec144e8b766eb7e297c08056337a46e0bfec90f876e03e6196b0e99ffa8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h462bb473cf6983dc9c513a45e8023addd819d394dc740e6c1ca84dfbfc341653aa10749fe4d4fef0f39645b973ad2874f04b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4cbe7515da2248d98be84d2c1d1241c9f4f1ae18806ee5e89e5deb3838131130374763e28e57c8a0949dbb44f42281dd6bf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c5f358258f38fd22f551e660ca03e4344e54cd899b192a65a71ce688b8a52ad5a1dabf0a51b2601737477e7f35f68078a7e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ca59572a37f99a1f394f543ae16237667f0ce44b6a728cbe680f9376743dffed50c3997f07e2e881c57c7e9390e97580cc0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bda7f99278220477dee5d6ef3230c6ab9891f5900d3eb5953c1ff755abec23c9b05fce1b78cacd0da2c1df1f55637c4853a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h15979b4e2a8f6821b7aaf6b5780a00e877c97a1e2dda00f2c683300a03c14198bdee5ca90b80690bb0d4efa00906dbefcecf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h632016098c128a3d920a509ddb2cd6db4e33dc0fd8709cd39af2a13025a8e425b26fdd9cd69a5dd067e3a29b15fb77b9f33c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21486c5e8985af49fe3c6bbe6bfa3b2e3b82ce87009570b76ce0c63439b3fa32e65c4cb60b32b1d50ad4306e3e8930ead4d4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2009efa7e6bdcbf53fdc89683683a3b9a5b602374b0fe5a78473e253aca3642076a76a7ed4fbd745e1324ec069205bda3fd5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7d300c1087e6a3ab0dcd2e3004a310095546a783a2f98dadddd3316ceeec8feb87de499902ca64d4d689e6839420a6460b2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5207069043adb12104f05781eb9ea981a27f80a26c57e4a3cd5202dabf7fbe4d61e8f8179a876fa85e5b5b300bbd645c7930;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha33d9b70111bc4e72a0f1073d7e066c43c9330aec57661a77bb89df0a16b863dec12a5d703734b95472ae1ab61073604cf38;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbf351717c508f60249f6729222d4e2be0c14e34eb36d937095969d241c3d0d707f3968c34bab65842e90e6d52c42dd3bf3ad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h435949a93e313bc609b1649b2a9ab42f5e7996a2a1374d451d0f9dd361fbaa9067e705c8c3fec00ede8a0bc81824c477193d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44ba1f9a0d9fdbd938fe7f7991227f25ce0ad3cb350642e4f5e879bb1201d2b782783cd3f6995285d772c3a0fd06dae42100;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99023994d347181150cd6413ac077b0de6fef0797969766439be0557cb339207973546ec7353e7a64527edc374d7c20a9959;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3952493a03c9d84ea54477799f5e2aced0c5bbe3a7a600c299835fdc4c42c266ea996798b23b56756dbbc1037c136ee96e65;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0bbea21376b0e9b73ac5c2bdda7042dc79202a94324205dfa992343104e731f059ab4410aa6186bfd74dee92cb462a8a929;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55634879b1e06c60e47bbcfaa2769a1cc0d54196e00e6e1cfe652f986b2e6c867cda1b63f7612ce87d4a6519efd42225dbc8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h28bb38256f07a65975fcd6990c36b6c0dceaad1b7195fa61f9b43c331549160fcfdfc0b30a36fd6ac9f586d7a806a935c21e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h22bbe868325df18626a325d55a76af9a34a598ef6053b2e6a7940dd2f23bac4e369d81f020e96bd43019123ac03d1946dc40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca104cd9dcc08a6b88e082257b3cabd4c08bf3fa20e823556fb8f0045f834214d900c316397fd349a242bdb66f36448111bd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h40f7c85ebf059121c16d48e89fe94b40cb2aaad0842079f1937b4b0748a7a3bcf58e428971febe8d30309655016d8dc6017a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ce0e61015ff13e4b4e61de9f47b9965336829f2dd5cc47050be98613f1cdf77a73f58c26e8d747dbb931fce4c4454027dfc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h953144ebc9d8c9c818f1ffc113cebc34a7ed16553ab56f74fc74eaa0306ce3806a9130e088eb81cab0bd6b0a4b7b08640877;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h21eee4237b3f389520bae3b81de4cbd8577ee2984c27c989365c4830330f74234c5c03c99e779fa551c99b33c9eea4facbd1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h753c6b58b03331d240bfc868013af734305d71ed2f31bfced0edd0dacb2c35051c4f9a165f69cabd89c2ad98220f1c65854f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17363bb9b5f0dec5fb372f14863db4c6cf29a1a5115209f4fa1089cbd61109b42e4e1c4ad2a9866ea8c63621399616d0146a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b7ca291cbd686beda14380209dce45ca6d063f9e1ef19c2c7f168bc3da1d65036e25f5158c6d5329495e86b4812093e1007;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heeadd83f46c8a9a211d286c7bc771a232167ac54029e5f4eb771c607e45b94a4624a4f6dc3bb0d18b286ca83029f57c79fb9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had0f0b9f5e1a464b2e07a95ab41e76c399590321f34b4edb518178aea6d6082afad9157ddf22798aa6a38d6792c25777adea;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92c61425a625d9c6048b1191cbc9e073eab5ebddebc7e2d48a8ace63eb3c944eaebc79241f3c19a5efbe033ba2f749d0a638;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h145d99a9dd7065c672f101ad37aff7e66358b545fca43bc448130cc0f4ec8d268c25b6c1c6535b7a2e761ea077b8e46d22da;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8df6bc4e303d85d01ec3aabe8fb3aaaa97ef5c5ebfd0c10b17ec17c05ae771cb8dc9536b4a623a928c62cd9b600e13ae974e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h943be491803ed26bfe0147ae812213815daeaa8ef001dea4c7dea405ee455dfcbdc82005bbe45097504701502795d058de5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36568eca9bab030ce2ee906754f49bb8c666ec7fd5fa1eec11085b3be2ce8eb786ecdf2535b6132c1063a6d44abd33634d6a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf71e164be5dfc31eacdb0fed8cf2a28e1d841ad6fbe528ce0995392669744a4b3b7ae7464c824207dcd7457a3943b4ea18cf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bcc6692e8987e1c1919650b2c73875077dde90e901a49499f6151f9ff74f49b4ba77b9a376603003e5825bad1114569ea39;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6891bb8e425f2ed995b0e38812203332f4593a244614707fdf1cd0c0f7e05805dfdee719346acf0910493174183a48607a69;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c79cfe9944017b028d142c55a640fa084d96b29d06f218fb07c365175662ab81e58e63080f334cf88621b22d314d295d5ee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44c23870f3ea5a0d1d08d24555c89be4f130adce4bb6410e770f38a328a7c1c1dad952c2aa0e7792cc902c4201159971f67f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5ec244f7340cbfef34a3c4dc2a6679652e8c1b651b445bfee297a80d93940990e5d3bc40233ef4fdf15f05dbebd34b7d82be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0ed43f2ecbbaeaa490636dd548d1e8a28463f08b0a878443cabe3ef8cd2a4558df87951e23dc84b634a5ff9510caae8ce7f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h29eaf9c15b23b5dc9ed6910059e176e0ed96ebe857cc01e463040f74966debca8b8c0a4f5ab0ac2d8ba517fe1c4823b68891;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3725009e306538581e66e49870fd2e269fcf5cee9e25d96e99265d10b70e08a7f31e420e3ab04dbf81abfa7b40fe6826cf6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb8b0710bc99668cdb386e8a2aea0ad4d2369195800c227193bc7e68360c2c5f16446c9094c1bead12c520d0aa16c370e2ee6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5787a505192863a8da9fd6d09d1b016dfced03c7602818dddb12a16866d0162a979640fbd238f65f7e900b1e903f665d3c1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcc09f1519c5d31d23cfb198e14c55c7b39e1b45a64a09f2e5ba605fdbd0437ed3300a6a6eb76e2c55b4a52b2aabb988e27c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h127d5aa36d089ce26e8de2d3b7c9548504e29c2ca695d97f025733f0bc68f50640316de85a0d8caeffc0c8623e3ab42a1ad9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97cc051c653e47665a1e2d3266fa1dcbcab66c308a96df2fa7b34d3fd6e109da56be0b93f9081b48e9eedff76a7c548ae956;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97e23763b228c0bb3dfaf2b713503b509dd0a501498ce88b78feae3ff18cfc47b6281701fdcdc08701f7e510f315d82b17f8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb79b0b37f27c97bfbfcb07fd19c3f25974d9ddde0289ade652a0ffc33836a4d969ad3e57b54e0766d4b46ef74936b8668026;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h504d6d88e78c8ace94c8b911f16fa0919d13984df1414ca7862e9819979283b68d327f5298d09f71e3c2e3ee22dff5fbdbd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe1e23b4cfd1dbab719a67a19d554e1c4b5eaa7c949657b67f8d9400180bd755a75778d613bc46460e5dcf8766375970edcb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8cf8160817d24e8e730e841324a922af7ae9b199c180077d09efcb1485418c3603b382a0d1fbfc850265e52675147bcbaa1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88548b287b53fbb40199e271fb3fa27e862a8cd6adc6612681e134d13b84455febe70f40f2714eb9737a7513e99d4ecb137c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h357fed74f24e2e9861eaa0453561f90b1a579bdbef2082c0b8ab3ccb26e14b0816e0cdbf1170af74382e7c1d1165c4371396;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2053a8ad95a043e90bfd256292a580a1a3e7861c22d85bea98285df0ae2d7344caeeba91cf38171354bc760423b08ef4545e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffa4eac6eed9414d381663f1d3ce12e92a965a106fd8177b06487c420417e35487436ef5c8094aca6da3ad9f35a901077f89;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11346584e0feb276195ae2f121625773cfaae13c749f817b461c49730a144406a01fdf14e1ee1a85846de6c04ba976454155;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haeef325cdd640d3d05c357d8fd367a94dc465e116aed9482cebcce47f47f06cc3caeb895a2f577d3e9f28f15621874c7c3b7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h733feac87b8de3a450f503ee6a9fa971019b499d900f17d45083886c2724449d1be5ae8a561386359ce7c284db4d504c669a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdef99a94c71c553220805145cdf47d7578c8670adfa233e99c03149b72ad82046bd34948a0f4df8f55334c3646242327912;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h574c5b9667a477c0c2a42e2d1742c5c9f9a0f6ea1e5dee7c470aae71b6de159cc28c707ccca7f870160125308abc976ead0a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36b1e6f915cb2bbb9d291ae8d77d03ee03e632046674ec4957b6358ac549b894e6c9ec26daeaafc9a550413f63c24044313e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb0cbdc5f70581fd2344849185b057adf9ce6bf44865410f3b90bc6d3d11da4b39f643f8022581f552fdbb79c4f1efc8b616;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadcc5c8e24dfa2ac28a69a62d7489835b399bb79fe02753d9ec7527a5f10f60497c9320a53d4e905a2a5dc17d0a80d494f49;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a006f7e5c9a7d26f8379189fead6c92852e3225e1ed4f84b6e696c241d6c2ef8410fd5aff53f9d6e650e22831cc7a9c0866;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcea27c0e67e75fe9583cbf6d205cb8620075a5c803089ed8b0fce34710d007f46b94e80eb2cc7794d9eb5f8a177c6cfaa49c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd50cea5d7f1acd7360bcf07bdf2cb816bc4361c45e54228c894c9b14fc34413823ce2ad7d0e080fb63b79eeba7cdddae99d3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h544df51b4c3e1c33d96ecd73303b5a588df9d271e5fe16b740a816a9a74ab6e8951a3369dfb9710a98a3e541fb5f04dff5d3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc337bc75011cbb70f5b8b0bb4dffe8f98e6721c6b6cdbb1889020dc98fa6418fa3084d18652541f36925d85734373c0d1292;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f7e24d17741c81df83004b8f80efcd3121776210b7891def6a88eded99b261eec772c188ec963c17ddc73e4571250feb304;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34cba9848a4b60e7b6d6e6c8a7821d0f3224bbec745344cce513892e88a2d5073a74365c3b5a158ac3bb7fd0e4774cd1ad84;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c8e7242232903d01462dbbed4fb4399147f5813a526840236e0adab89d88faa326e932660d587182a64e0cf2edd80133c25;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf32a5d1fbc2ac9945ecc8c71296cc0e8a0d49d348e9daa4add24b944e64e48ef164a78d6605e8a4f47e6d2d814ddf9c5d889;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h85768394955f4bce1d6afe887461b6681ca09013826647f012b5bd69150239d2905f68fd5d8c4d92ba44aa618b096cf2989;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3f5de673e81cd730ae364049f9e47f62d9daf71d52eb43bb17559cb55ad8b0d8978ee7fd7937b86565a55ad275190fae44b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1e6f2fa7e0ebb809e82f32c47ea53c6b7c85a600c2ba24bf6ce636f1f396a53bfdc6ed26dba273f291c4487bba10a5a95fc3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6102911bf2dd18ba08806c52fa847c041a0083ef78c332a84a82af27ec00214fce73588dcc508c54c5ab87b6eaa1e9640517;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0c924d38227cf0386e22daa267935aabfb46d6a7d34160964521722bb6fda425702d14d9ccd5b5e5f478118ff80f65fe7ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcdcedfe57a275c57a5dceb7ac426463e546b5fe187ff5445ef198365dd2f84353eab4a60fb8b26c3ea9072afaa6d4a118d81;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h778d0b2385c3b9dbb269b382a73647edd89bad38408fd68cc2c471ec7b9d12076482452bb5343255f3235f4ea2c4b7373d9d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h193fb69bd3803d80c60a3ba5de1da5d7b4a7ee9fe182600b1eab1a70a0c373b5cbaa223f0172c6d1e327ac05c7950c0df5f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20bd3ac9021f1d99beafdf441420f5387a104c5df24bbe9f62d5d2ddb060aa7238fbeafeb914c806bcabb094324a520803b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fc2b1a9ec383b47c1affec4ece9ccbc883119158fc292b6b0060bdf2771957714f9342e9d1b81ddfecde969012b02ab9ea6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h741ff00222a001d4351aa3ee7382b97bec805b50af2a96cf4e270d3c9b26c785a28e8f95b4dda2585c61c87120b6c2ce3bef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hceda161b29e2983c4c90f8d499222c84a4ad39bf3f6f25162144c87439941c72eb7ff4dcc865ced5453a33c006b72d914e7a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf078e64b8c75c0dfc24e29120dfddf03d87d79bce86c94ab714dd42500f385f45480eef6ec7407fbe4c5e6bb0ee52dd18ad3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h386a0889558a37833e1c2969c39891803c9c052593d0be98ca5b9357885a86594fa942f238b845bc3f974dfbc5bf35fb8045;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h132d76e3c0e4e633c616ad8a4f68fe8a47d48cba90caf0af6338a11144ce1f3c9d818bf37124fd99f6c7942d1a928bc9824c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26797e0f852bfe4f6d872a7cdff895575ebfa5d1f4d432e2e134a3d818c74daf773608a73bbe9ac7f843b08e78be3199f12e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38ec0cfbb3e9107c58c06737760e36e9c9c3cc8dbf231aeb0a6375eff936383463075cdc98f086cad39b93afd24c77caf744;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc9740139d2433767f7211c7a2376ad9b4cdf014b6a36bb647f9fa86ebb4d7da5ade3d37564ae3e8476c094e6af32a056a32;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h631ccd50aad738410a54955c8b5e227259969ccf961115a028f4fee844fd4ff0d4bf1264f7d9b21a570458ec2dc0639c14ab;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h321790551c78aaa6e0a4d452f7c8d348c8f1849f7824b3cf0264f77aa1ad2607a8da052816092b9f5951230fd05a5dba6e6f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e43e0b1bbbcbe0d8a23518452a98a0e3e249b936cedb52d2c45cf0bad04333ac21a4c3cf87b49616d1d91447401646b2660;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef429d55ed5b976b2d055da8c0c096bdab53de08dcfb524634f7ba4aa5ea95d107ed2b2d9ebd5032de04d976aeb3e891431d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6a059a3f314a29a13364b09bccf9c245ffb0f6d7c06cea40d59a4c6eef07878ddd12e032b5818fb4cceaa25e8df891d79efc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2424142345a004ddc1ecb7a129461cf3039e87301ac4335d2650df73e48825e912ddfdbc81ba171550d35ecb4361c7937661;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2ccec9283d4221d6f8b34e8f348c494e0a4b30163295151251d7ec6cf86f806510d4e5572724b9eb5d9ad6c93a2ae4086dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h473a4488506b85f98788a54aa9a8f815d4c8819cb65be725284b48a031c2ef9c97a1372932316d434a10e87369b3d68e2a98;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6dd0105b3f85b7b9ecfdb29a24fac5778ba8b850dfcb0c5396414169844d9a524882d1c32f39211fcefbeb25615fe6115d21;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had4740eca6fdff8d4636af900b9fe3030c33080fc491a8176776fdbc193404033b04fd3f2b1b1db9e2381258bcf4eef5d0df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h236edd04ab81047abe31cdeeee7d0654206ef45e6b96016d58252bf18cdf60233bccff2ab27b314803c8b89fc2d1871d347c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50e6d49276e69c8dafd22b5b154ab0bfb16155c109b99824637eada1a921df7e4c11ad06ca180e8e6f351165c0a9a83ac25e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95900b9f2d7a7b17736e8d31a31fb10b493fd507dd224ca2e444c0a1c5aa69c6c939abcaada1dd3b659e8229ed21d7be0307;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hff8a22aa34f8392ccb560c9bc2638e8752522ec16f11a07c036d1ce64b19d55fe33651f7690e9308c7cbe343a908a6f93a49;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf02d00142e1c4635df6b299002027d65b27fed67feb6a9c54ac56ec241e80d24367430d5cffdc4a4364fc7db29c9e4dc0ede;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf516d23dc4a96ae0fd0fdeb905e463ff0bb9e25aa92cd1db51ca053270ed86a03ebbd6dd651a003daf83c7faade6c0195b1f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hec2621c82390ce03eb4a260f07c883a697df906f76119531f1acf4ba5a3c38178d314ad9823694fdc1939bb2dbca53d00a90;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h576fd790abd49048e69660e0c95cce81b50ab2aa96c5ccabe9eaa8050ec86ce196f3104468354467fc819f6b3b647c4e1476;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha42e8c61435c72a8ae1822418689b402e7bdfd01375b1a5d78e974dec25dbfc297f7db539c34de53f2c4fc251d0b5a916672;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h205fe335eec72fbac547a2093ae82e6b74edf8c2ec01f59fbcef477630b6ac0de4b8934d0654b119245a60a5f5d5a9528aaf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6934eeae0f2fa8742faad2d30338e534de2ed44df0c75a21897bdc6e52fd614d4a74f7c3391d61ebf851cad25be321b2504;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haced88b215c1c1ee2c47f18a7e16db870ce6a0e1b22db3c39dad34a91e643bb5c95a67ffeee45ba857d81be61999dff4fb74;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5755d368251fe590cc68f83388c4bdb9d72960b6d624b87ae213fb54352612625fa694b5f708d93b20e0cf8d4b6365ca42c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h417998b94927126622791d97dc3247e40a1321916a979da172f178727011ee0bcc5165df1fe0f6ae73ac305665b4b9acffe4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86ba5f6002c9a016790606dd51e470c5dcc3e01c31ba56ffad7bf1e039e184c7b61157f65eedf1d3f6e2e6e830058b8231ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9e6c5c2e3be4ccb7341d55d2eb567b3785afd9a6a48285736e785445517422ae855fdea2055090b4a5f662c35cb2200a263;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc59b0c042ef06acc5384311dd1c9499d78eec26837786c1bbe7dd0e5df212433264e54cb55dc1eefdfa1568645ce5849e008;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h761d979bc87349d2bdb7385ade176e13702165f7dc012077821bea5118d8a58bd71d0b4e9fb9c57cb97b8552057a12b8a68c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7cdc6c1673f321fd0955c7444c0d8855d84888bf0053230d7ac98348262ed09c59fc1b19df99b140200d96f05fb1967c5fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfcfc49e516f799e8f883afb70bda63385cc6eea9baf080300655012f4e7e8b573e096fbced9527398f8778d1f3347130b884;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he9760072e5ba70fdbe1c542c4b9ecb27862361f3514424467882900eb4bde4b93ef86160a538db97f9c5eaa7a6306e96f6f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88aea1f0e2435907c6ad4a1c2d4d2dc48001f251c1355aa1d5f4708ab5fd19d20ea8fe7aac0ff329cd6053a5565986fe1c1c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80f97fec520544fb8dea9e98e400fb0f7638505783a48ec4cabc9da30c2d9a177bbfe2c8a6e9310e163e539dfeef992298ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c158f73a462de89be0b98efe816fedafb7a85b37808aa1f4858a77ff4f884ab440e06804c02852f180d37fd32cd4cb922b3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7358ae30de1132ccad08d87128b3ac6a5a95bbee82432c68d8254820f0b3d3b4a42725f6e98cf28e8d1f5eb3f398269ed15c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f38cf49745e85abca9d325608d2ce091c38eaac278df5ad4fc71234a9d4e194735bfd627650e129f7947a0219d1bd85fb9e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6f79fb6940ebb2fca48e43827f5f75791d66be2e66e4989c8f15bf4569f29d6a548f40600fa78341e78b2038f7edd5c15b1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0378d6d04ea0456a5f1427f3a00bfec1e5752e7efa20348d8d6a637cd1b22bbb83feaa1fff75e4b926f211023ccac3d4d4a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7710e1e4ffe76c08c37bb45d3f3f941158b6028ba0ff138b5eb91a9f663c9c7b4db07da492aad863444801a238b1b7cf113;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7c80709f725bf9ac0cd778f8ff23e5400d51f0cc854418200adef4097adf1ad4739454a0bfb420243f8ed7b03c123b649af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6b4d0e37a2f21bddf151432ef881ca6cf18bd5411e9c2b34ca15825d09b8304f2a0d1f58370219084247e0ecc4cf2d33e795;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2099b5223219c15386de2556a9a0853d75bd97ca6c8a449317be40d6ccc1d734452e36741a8b635046f7ef71f05a142672ef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2b63b3b24e78c2b1e8de101b71727ee8db511e68caa1baaaf5ce078f0ad9b1d08f2eb0aa3c24bdf36318b21c85f4aae172e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbbff67f7c4f82faa4f5acadd635eb0f4e21c82eb5460bb2266478ef5ac8d8e02a8cb862e0760729b3d51034be168089aa55a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49902eba94ed9130fb6ba546c4d20511bf7769b3e479932cb46ffa4e88cc387e46ebc3c083da08df0ada13465a6953166a21;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h936fa18676c97b398b0a350ef9792109dbe3ebda17283baf2e3fb1f8086f0793d3d94671f1adf0d227c11be02168f2fd46b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hde2ba4f317e6bf8c35840ac96a7acfe760ec142405511d2928b9f0dbc6fc8caa2889230bc0e75671f42d0bd38f1e2e19e958;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d805bcf89ea4e9c5f339b7730070512d8948b9fd57e25bdb7601bd137f7bb193358e7796b48317135afa3804907a9f3a9dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44095a4f5b96ec8a7bff5a7b216b818d2c26c6c9e49d0dea8554133c93d19dbf84e779b033b889c2a6548cc1616238f30f75;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hadeff0ea0d9817df6593c9780c072cc5e6d3c780209170d2b58853ec154a72f500959d80c02c828c4a1db042717254aae51;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf38d0447b0bda930b5d2fc5bdfd1660ebdb288b5e8166fe9a06416b1606b1eb6363f885d8ba2bab9d2b114430fc1f9d53303;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he38f42578a5c34d57c6b33d4331d982e342bd550ae2a6a7d2796b53ccff64a5ba2c720268a9c54be27ca984519eec050f94e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h44d8a664c4175cedeb65f6e46937616521ab03de8a26eefaa147e964cca7e56a970c805f8fab769780c084bc808123eb3bd1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h64eebf9db90e30f29c24e328e7f0a42df7bf489fc4219cf568ddc94850309df4214092f2d5e21114e11ab538da11e3e97f48;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7d73017e5057ad1f68f0ff109e2747383a380c3727fdcb754605146731a7e0b2dcec4fb2e384d9e0fa67ee68d5d6c4b66f59;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d16b6caf40e52c606af55e3b11486a75bbdc406956d0fb2dbe94e37663f0b59873e3db24c31c338334e628bb01a9e36a170;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h14c45ac8e997b63bc89a22da31c77e0148a4bf8f881463c96b77459eea543b45c2a0d3fe9b6f3ac137dabded5fb4047076cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a993dc67c048117b3edb00450b4e0e3dcd16b6e16c81cc3d641bfcb4e858fb1f9d4bfce02c0df4cf1bf9eff44d41c4f2706;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd1332e5622d30d86f50e55c432611c3eeb0f249e8d5875d635fd2e01531110cde58c62dfe5671ca663250ca4a3714b78e855;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2074d8eb399e06ee7ab93e0e7b3bcee7c8cc99421ce6b14373114668c5fc468d587b60868a83e8403002f1abba76c1df777b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf7d95ea4adf3e610ce78c6d0cf988aa071e49cf92b31de4f00eb9eba8b8b1fd7412c714cb926013d43d25df078ad5a365cd2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d6bf7ed2b0765120e1a31332922881bcadd3e066198f3c34233053d11e71912458f6b57b0bcbe4ec702ff8caaa8907f344a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6ec3f730eb3a0b32630c1e0509996ea5f32851887d99123862b0b2548105192a951271c0bfd550837c05d9005f42ff854a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd909e53bfe866a2477961777be31ecefa00e5772fbeca1117b2a77a6da372e6398d89632074422788cdd3ad538ebe1b750f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h269bacb362a3f267981e05edc5b5da4f3b79f573ed2499e959557150f4e3e416a14e3b0ca39543766d1322115053fde2d1c2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5435f2db358457d0d1e3544204564c44a7febf60c8fe35bda6f556cdf18450fe0c07ede083cd339a467d73d6aef747ad749;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf27b571ffe12ffa2ded91a1c2ccc88fb6bc469833bb4584da67f97b32206816dff2daefca07af0155278276b4e4594f4053e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha697f10ee66836c5f1aaae05d6adaedf740152dac41aaea140381d5b5d59e7097f70177b40cce23b9989fb199bf19991ca2b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d59b1cfcb80223cbcc821593595f63bb5088370a0d2707c5a618d4514eee771660761cd642f3364c9cdcb4dcebec6417176;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h146bb08d0d85f8be9fff94bff3d976fd43a0ef921b3f793c46e6814002e61ab37fba18d9c3937632bfbff074b9a147e3e705;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf15b083bf135b3465ae7c3a690e0b650bf5b1b50d3b5fbe3dccacaf7a54a5b247b97018f4b8cc2be384daef380512fb4038a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3fc7b19b027dec9a9c6fbb6ad416a8e062fbd9ac122c2bd0a3d87a84cd0e3e7357452f509c91168b22f77e378176346344aa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6d97a8c898b3370e6363e69c9aea1f9e0d526bbffa7584451abe5092ba34590a4fe76a9366762553862a19664b7b6d24347a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2ebe054faa8058c73026305c86ed5d70d4975445bf5018350d15d536b578fd2ede26321c5fb4debfac6c8421c87f1896e2db;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f20626b0eaddea5aedd6eee8967c36b0132d5f8b77803e96adb962598b8b4737b4370cfd4f5d0d8b12b284441a6007722a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb181205a2bac4b192ad042e66158cfeac3d03d6f66a6dd8fcf00d8403b2e1e55ae8e7a1818486ffcca9a3cfaeab86d69df7d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2682484edbc2d063f63db6fd89012eab527a992de7ed8ecacf08ee5b3c06be23c59d363019cbd443129501bacf2563b0c7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb852641c18cb164248c05a355fff8463f7ffc5907a6b064cc222a8b007fc02a06875fa3056564cb8f29b6857a22afccf06a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he0017aae0d254227cdb0dd379f164fdd8a183e0da9e2f58701c73f8368ce84b00fffc0508576163dc08c08f4dcb818109684;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b0d89e5dc5aa1fd8da4ebb8e36e57c61db32d6bb99207d10c7804419ad187a50aa0248329f3101ee2c132017fa449de61a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h62ea1b5023fe09e95bb9f80a9c3ee962a7584f5b663f0ac7d2f07804b86572ab52d369e95a84b487760adbeeee68bcd9148a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6fab0d4d04a8c5d19da8b61bb7ade7ed3379d6f15a168d488ab0b6efc062f3d820f97a929bf8e26db3c7589ce514014652d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f6b6ba0f8ac792eb51bdba55abfa9362ca4a8da1a25721df00103707abca7ea11a0156efa734fb05bda5e5042cdacfad194;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdeaed2bfad8297581a79395c33912a47962d476e476a489cff9c981f55d6624a83c73d3eba71206a47800d7adb56fed931ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96e54e57d169600fa4fe6769aa51ced55f17ed28fc4ea1b9f4ff35e571b571e93d63425ef8f2f002b8ff3ace2e4334424170;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0d19c2431e37bd8786693b2472567768e690877a2ef7e9551bafc0d69bbdd7ad99f206804591940d8a192ea7bef12d0a43c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h20262ad9be3831f95f38959530be61843ac1171ce84b4106cc430061577155b324e62f0fcfe92ccf36a34b091a66dbc32e58;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc996f4400d902cd00df8503dd8080abe1fb4ec54c56b9e9c60ed1c93f6377f5a48642ce630b495c0f3099f64bfc178cc44fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a67edf81c1db110355c6b90843c734aca579f93b15d1ff3527f31d64298c43c4cc0b767fffc3f6e2a958d00c7e6a695ef87;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3bdb7bd594f4047199ec6dd230a3942a2dabbd4a5aafa471c0501373d87f5dd31480c2b31306228a019376d4591812264e42;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6ecac84deb934c876eaef9f5ced11b1e2c2ec747739a561eae7b8bab47eab9bc701a0aaef4e7a7ed8090c29e5e2ffb973b5d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f18d91bb87651100d7a2d6e3248cead19c9271fac9e83717ed82ec407e75167cd5a25511af4c0bee03c13f81dce1288084;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h89f8c62cfd9cb0ae18e1b06321b9434c77921c254de5649305db08a05390133535a72db5190be60f3233ae05b38bf5ceabcd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb11feabcd2ebaf28152e18287f2d6418201cea0304c63ab0d6c6b18d6def5501617ea1895db02d9c42c56ef4cdc43c6c581b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbe4339efc045bb77985cbce71ca39fbb6b54c5c4089699a122394f085e44ed532bc32f57b535f9acc88edbf91846f616c50f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84b3c781f6c6b26895e20e5416361a5c72faf1f2129fe111705ea3ce04872f90ae373ff733f559ce5aef90a7726d63a5fadd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfdfd5f1c3225ac6ed0b91674f42ea31578aca24188a43de2509c5daa707c4d27ce1986d209c2ebb35b48472385c31cd98246;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h275357c745e0bab652aa37837ced8c829e01df8b111d9595199c3554c79062906b9e3acd0eda54e7acd110ddd6a20da75d3f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h78abe92f015151265fb0c1f7cdaebdd9c662af194399151f04b9f2429c8e63b3f578f61fe6b220e2bbfd1430074e294c63fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h436d17fee57cb387a6de969e78942c98110c2910f956170373468c66d75caa6c1889b4d0697b3b07b50679285e834e3def09;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5431dde5a3727ae01a7f269156be584d4c1d8902026d971ad3049e54f08ae69f31888d3e1d636a3b8d5758b08dea73e84eed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0d05564d430426533b1dafa8c300db11ffe100ccf57929fc8a16dceb187a95b54b78cf71a64aebf239660137438316cca89;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92e9906a6bf388af9196d7faa0acedc6534b6c1e9b58c2ebb4ddd1bcb366126e45110f1877fc1eeba9bcb51ab3d5451b0843;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f752e4032b0eaaf5fae8f7e16a77f432a05aeba923563b98992d2558926dffff15cac5879812494070fc5117ccecbc03ca4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9459ff5987311f6a2a2939411af2dcf53c558149bdbb5a8f82002a62ce4c794cc6b16f2d3d67dab9abd266b23c259a497a8c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f49ac25cff62238c1be773ceac184f1887322514bdadccd5e0ae2c4e905a23c1e8f9b07c4eb9ab4fc74c1ad00220a4c267d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h969c9baaa46f351bc3bc4aeab9de6eb67fd8cd49b307ba3cf2cb7a142660513be16d04d07ca6f8a23bcbc989a7bf5cd476ff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3eecff795e989f5435da257ae4da6d72e179e8d8002f653308a2d2905c71304c5b91daf4c4ff00aa5cdc376de905508bf146;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h624c8b09822f47ced80da562043b7f549dc67a9011fa8482c99065a6af7817a3c6e971f0365478c481c541cad2c2788b8f4f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h306b6278c690aaefd6dd474bed9a2347ed2757cec9e6272d6060303d2865203f67df0bbd6231f9ed5237089c971b9968eee7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h903f248002eca97af51beb5058d6241afd1e8fcc499bba72759fa243718e4f3d272f50bb1ff0750baef70ac8ff6cbb5fdfb4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce6fefb8719471eefb9b687ff70d7d1d49575f2b650086c142041bd51c575c7b3a048e94a3c64edc4632818cdea495575647;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5d26faec85d554a22d07d2832b9fe0596490f1c1bc9b779cb3fccf1055b72985144b101d4753e0f2f27b71c109b6ed3d0dfc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd70562736d964808ee41117161dbd4d2ebe950b539c02a10e7fa7e7b5579dc184064e650faa51b09b3bb232c7298c5ca0ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25df7bde7ad73b0537d7779bb1ff6646180aa06d9604c087e5302a3e55d79cb1632e07978a5c6b6ceaea9d5fa77ed7a46f23;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h790681fad6e9bb64d63a14a956e85e4aaf15efc5cd3e384324e8c77ee4e4eca24a2bd2489be288cbefea620a82138c041fd8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7716600ca5964d5cf3f5707408d7e4cc638c803b6fcaaf1415641aa4d7f5627a68be21e62a25f2a65557fe8f5d0a7426ec9e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bf5ca973a27099bb023551c20eea0a0f1d1e1ae8eea0c90436dd0535dbfa0b180620c4ea80f797150ec2a692e7839e1c4b2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96c0810d483794020f8122312fb0c411ef3bc3188a95a0320112aed0efed7abc05ce27bf3202950ce6f7e3db021830c92c3c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4a031f4f6e5be7a0480e0a403f208f6823e2049a874d8cd21d82ad4e4fae610480cbbb4d713c0d0d0d1e5617af3f1024ee21;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7df8a5a77baddebf57ae363f3d50671ebf813fdecba9125872ebdcd2c79d08936a5fc4956cfb303897346912f020b323be1b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2facd7cd81e13cd4adbbb7142cb67645b34eaa8e91d5f6dcb16e683af75316344a883b12b76a3ce7c01bbff6edbb6e9a0744;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf59d6137280e5644272df96cdab7c0db6f61f8d41ab717b080fbb2a44bb9c665c3ca0857f659762677387f343c5935abc457;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbf5e049e7da5fd3253c607848c2f3503f9c24acd05a0d35a3e28f2023af4ecebe32934943d1f143cf91733b3ab4cfcb9277;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h48ef1c1b627f3bb14c3d20e2ad6d8ffe9002a75a87e9ff68b02307d013cba0e3d2eec18f88035dd23187df030f4d1d6e268a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18995a12461e4b63061ab8d56e1913d206267dec93112c046f96b1224e74b9a5629cb1d1b8e165964bc7533fc636dee66055;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf7559718cf4ee27ba53c0ae19e72a1b57dd070e9d98a22586beba462ec45cd9e6ff780e260dc76a916a443c3b7bacecf74a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf541e0a91d804a6e9f206eeb4f08885095f967bcd20a195fe43d556519efa059975e039d97feeb2d6cc3bd345a405a106ac5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he59dcf2f3486ca22fb52825d6d36b2caa540be34fc225158660dbe349ba281ea2c61b124a08c920e79ea5679dbb7651d06fe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36ab9fdaa40e62b3281d03c82dc21369009800c3faebaef797f9ead702ba93be705abce928dc39e251ff1097c9b720af5b50;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he1ddf15455d097c52856920c962e9b71543960729ce4147d81c2c205a925e62ee39903cd293b370ba48bcd839c4dfaf59ae1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha63114e001150391ce58987cb6b80e7be7e61a86bf37cd8bfeb66a225cd266f0052e63794e2ea48b008c62fcbb55057fc0a3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2497d128e6f208ea2048a6555ab382819c26735941540d39caa180ffc8c81469568eae0bf1cbac4091abb7d6733cd0a07ca7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb63509b28be72b24ac062f039205b6512909ecc7ccf45c1012528d7165917e66ae696444be374575e5fb12674b1895597d83;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b7dcd9f972de23f334c624e2ccdee8c6f473030d29a91c10148d9b6b2d69f318e64142a6e514e8f02d70e58de3c202333f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7773543d1eafeb764d43a36d77c574d94261d1234410dbaf28ef7d5d94d31c89828710bdb99659ca30fa951566a298df40ad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc250f21f27a4009282a0409572015fcdb2bf7fd5841bf9d47a042e62b50b77711562fde6849d63cd465208f92707b9c48648;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9720f95e8a4b9d7efce71354aa741d2b3d79a4b842ab940c787593bd018286f83d2d0261307df84991abdf7b90c7f004b11;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa11eac5bc14ac6a36058e5fe15d7002923f0cdb7989f455525585743ed8b32190195caaa6360d2515190b407961db850f53;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9014662f9de2b1eb5832af858a049e37e601aaef0ec8f87d69e23eddc7628fea9052fb3302f2fa4bec46b598c5a672ae9b2a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93c5bebf2a3a3bd3ad023c0ea76c031cf7abd1d999e9442cb1f9bc3fee699a14eda8addd984bfbde0679f07dd1e1b379f9ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94c5ef7576f927cf72ac1995ac41d8e3469beab18ed08a0f6d86a682417aab813084f65fb22ee2dc514ae1585dfa0e6222ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f8dda85b517c3c139c5826c3ae78835b5c09541397e75351a56a84023cabd9f9344061d6325e431da163bea05ace084c97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8144f5b74f8d39989f7f41915260b17fe48a85e8980742517af321b7493bca5cc18d19982a01c193a5b880671f2c18908baa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7448234515abbab22c623bdb90cd061e026fc2a633ad116e9a344462a52c723cdd7f6ef90f20eeb1a89d932110d5fc961285;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h83bb4d687bcf215b6d03f3eb370769c9707d485d5c4f381169039f23578fecfbf7697eaf7b685216445ce2de7a24ed9b5613;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd4f336819955ea19dfa94108ff13f42ea8d30580fb1f4b49b1fe202566b025ea1c8bc23eabd33dec5a170044646d0fba8ecf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha7ae7ab23cb5b5da580ae926a7e840b502d11226ef8b552fd008a226035d039ec3fa8f0e34458ae64dca33b44850271363a9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h96355dbee1194ced801158a67f31a968e280bd4c877627e5d5cbcb3fefe22cc8df071903dc7bd4c880abb6ccdcd6c48101be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h276bc53add029cc86c972d68b00d865e9bbe79a883c6e057c299c9b0841f48f0f427f74c93dcc6b0ba4c86f912f8e24ad26;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a053416aeb2ba6dd84a862006acc13c52591916ac5367ce254ac8b41a733bbad78ed90d87cdf2209b0934eac3fc8c8ff81b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haef51a92fd1d31bc66a5399ab64afcdcee1fa293c19a75f2bb27995126a9cf85481a56363b493243de1154103b27e6e2f4bf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7eff6295f69d563c386d84fafad0817b648a1972a67214b684406c4012f4e5ff012bd2f8fa34e50c1a942e3a3216115cc306;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8fb4c75d3e120cb94972ce82e993d5cae2215bca70b963acc2f404a2d6ae245ebe257bf110cc39a7371972c17607081bc25d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h276782cf9b073bf452bf1281b89396fa503d3ccdb2631fca718f2a74626e31edf8ba46abdfae747c5e401e7055e942ff2c9f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h812a9f22470e0d1a11170edd5696dc7b1086552e03b15c7e02992e34d8c8d79fc67df6befc78f6dc1dbccbdd74fcf80923fd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h770b573b47f5c32717d053c74355ca4be8b0cef0085260e3867ec75ce4a8e83dda57f8b783d44ba1b7c8d5653c9517845eff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd20750c97e290a8d4eeca1ee40f1116e61d8e9f46a8d373f0b80061d1f325a1b183b96701a7a67501e867a2048836bd7696;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee8b4216610b62e3bad2d52ab43f4c8f251c810e95f757dfbf6e776bed31f08595993878d6f94f5a28dfa9a62707e80be9e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82e62f57b6af8dc7bf9ff0e0f28b6312ee7fe9eaa605a7ba42df576690289ac6b5fa5380c92191dd06e3ca69c4251f343430;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hea6051a855b8af541d401d6c71f16aee1e8b77cf18717eedec3ddaa75cd8d4ef6ea44d927727555b05482485d0442e84f2c5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h383889e401b30ddd7cbe151893d14b7cfc04b751427845cb3cef94673078024dee660dc63bf03439c35366206a1420c32a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0fec2cbdc08fa865cb5840553886ebecf5ffab5fe820afa0243111de71b67f5891cd0d5260aad325d5731e6e87fa97cd7a1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb088c2e2a4fdee2f565cdce5bf20aef11c59b5081a60a5e9aef2286e6de8216f4ccc6c254c73f9e85b895bb49149f842c70;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e885f5548736888cc5a0e75e6c858bd5db92a90b0008af0d5804b84a7bf02729f466daaa7b9e62c6a4af8c2cb4fff25b86;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1ef1a9631440aacd16ca11e510b8d188f289a705909bf26abe97f9999fdc356caa2acb7e9f67dc40a12d563499836b34032d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h675839ad6323401fa36268971502829038be2872f8ccc3d99b74a2284602abf67c1b7d0476e497c1cda4d536ab049d58c60a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heea10a73390fcb0d9f711908d1ba50a0efeb4dbc30e685c890ee58a5d203e8953625c14ee98dff3049db2f35e8c7a805ce63;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95bb20b8ab27a97b46d316c0cd82b0a3cbac1d6e666b4f9d81b45821bc5aeaa3ee9c46c8e273f7282dbca77576baeee06a4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha745104498a7baadc6ce88fa4f79cb06d84dd28a8f427ffc8d16dd8f23b144595947fc024baabd7fce1f04d99d2aa9d19198;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd27b4e444b6ab98fbfd3141df06e12581a484add88c54ed4712f5ddc6149d480328856ade339fe982f9c7170d723727bbe03;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h84b29ceaeab644abe95d32d169023ac7e03695186745c1b7072b3af52c2594e2878e7c5ccf6dfbfde691c523eca0cd016e6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16b0f0812862b43b7ba3903d7f8abf7de6eb983a84a15dc39c1fd9bd682f29b894aafab504eca433c9daa6fdd6e29e83b41e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1206d6b40f33934bcbf2c4b3a3952cc3b2923d6e12be7869a6b49f3b647d0f75f51eccf1e7d1a6ab5ce15491a6782f2e161;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bf8a5205ed7e3419078568acbc6e59afc4b60ce00d1e96938ba28c9d69118478d705ce6c326f2c552887de9d31b20af12c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc095da53c89c457e7cefeef4688618fc83e1a003c6b5ce880ca7e7028d29d75d1ee85477b4019792e38e76f07992b1f44314;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7e62877322c7840e47159ac8bdb7109cd0a3f6dc7d6072fdce0e925092f2df79855af750f45dca1725c97439a3864174240;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c875187fee56bc9f807414f549a41e08f41d17035248694548be3fa03fdece1a78c81b187831bae8f7706895f89febc42fc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb90522985753ee84dbb6eaa1195d7ef2e6c6ebcbfb0391a5bf833531a3d873a3ce5ef24e2c30667dfde71df3f26d25304a38;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9bfe59e71a8604def65113b543f0e7f4c47f624dc5c5415af952c59c4ecb1318f136e1e36fe212a03c5c248b7c8db960129;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8bbcf6ddb96614313ef49957219e4220610e3396f6417b6e6e38a4c29fe87b421ded941197852177042df4856e85e124ba49;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf821748b1d85eb2b660d531dac0e7cec6e8979f581b198a9917c445e318ce6a1b708157f625a3f308a3cc287ac483012f95a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfa9c73f6d3c9fdf5b4f80039a91fa329008d3c72a93974b7b76dea8c8b8fce88dbc2fad411e4e2a70b0c87cc57680656ed6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2333a0f78ec8d8540b5780c2a028caf24e6efa8eee7596068f75bfb4081cabaa5ccffcfcb1007de921202b2fb7e30302fa63;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2112354271368673885a994626e572a1a5bcc81fb31ea1c083a56ebff538191d92ef403babbd7f414f9b09d32d0eec402a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36f5b61283c785e26a2988c4e098e59d2fd63f568caa10ee45a4db1df91ba5a24da35d81449536d209850b34a8b5db8fbb59;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c66045030f0898c71f5925eff77b2abdb0701972e25bd278e7c647406b56c5278e83641076a89d9b117c61ff6787b198a4c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cc853756d21e85879faef348f274a6a10874fbf89bbd775a5c772ebe465889056364763c67b9f01534f808e98180a035e2d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82abcb253b58fcbf0aa5d5b50d1846cdd566820d59f7792863380ece5bedfd1eecfabd921d10572710088671d54934074f9c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haecc1586414ab40581ca8cc83a412910b8cfc60435ea4a3239de87669327588bcccf878246a2ff3a532209642a3e57f7d700;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe85dfb954188cc20affa44d4cd515b72e1b22e22afd3a6c65ee5c56f8c4e53a3b7e41796805129f1bad9847192610b89a0f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6854a5eb836c38c7836ec0f394fe6acd5215b82933d951e4e1cba524333380c03b888ad4f98e47ae5707d0737df891dcc86e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he6f43d02d1658b3f68c8c92240e122c68b12c9bda1e00e4e9d6ca579737a356b6e14bfb142718146a245bcb36bfa21a465c9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdef603e81bcdca7665344aafcff7242f4e4e3312684568ecbee10905680560dcd75a1e540dd0fc6370b1ee524ded85e5654b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6274ae5598331b48c665f5817e2d64c8b542c727d8a719d5d926b4c14a1d33e288ab6f27e11bdc8d792acddff55a25c0543a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h210d22ba62eebc0f1008302125e601b51d4826906779640779e31a093946fe36373b003b0b91fcb8e3e34546845585222c27;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2d359c68f3f796557c9820491d4130c36c40925c69f05fe9dd52a31240bff4a2f9b5c82182a3a726275d8674d644d5b7016;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7e567f8fe9caad6d9e8adfe1c2c6407a657b6f18392ed58db1ee92fcbe52d528dbe221baa91e73b733448b76b5839ffe018d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c93fe1b50ccee837bec5e26d2dde9806f4770ed9dc6022b9ae0ebd8adcb857642a5b17067b42efd9eaae88eee54c8c314e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2b124f85bf5253deeebb428e5e1bf6ac08526c8908148035807e6e2f3e52c83b1d6ffed7f86f2f933a36c17706d03283332;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcb9d268c6ba84efeebd710c0f73111913a17dd8e1f9978461ee6c2eb4e665128d797f8ca40f2fb091e37e80b314cbcc9e4d7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbae3d2c3258a10b455bc049b7dd41622bd3ee85341ecbc363c1fb39ebae48385cf1d008c15f1181a65a0eb750eea8e15d4a4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8d85512e473874f11bafcd2bae0295500a18a796388e6ec52da1283252113a4d09636f238924c42770fca91289b9951fa9e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4087555dd270a4abf7d84046e6a93b0c70781fed25c56f2fa92171d45d6e99a43825b6eb4da2d23243483c7c2572d33503fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0b14bae9869710e3fe3bd9f5537d9f8b4cdd050d204902610b28ee8b2c5c5b678b05b40e3bf04b3ee7b84cb06224363b1e9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h683b334a2b7912bca40887bfb0ac93bba35e1b1ca4025bc5671e005cfd78fbc6b171fec5a711e307c270f1d30809c529ff97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6f233a242ae0c8b005e23201e220d73bf9914445d2bcd6db297e4524902b68067773c81f6ac759f8ae75eaf148f600f706f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc14eca3a042773c0dee78f668bba22dd33baca59cba98ca7849e3445eaf1b029e4eefca2b2a94002422ae831104463486c27;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h287a197b52fcbcd1fac93df17f50ed9617b35dfd44e760fa0e519c1a6085e9e324104e0b5a35f9d9c25b12a52a5f41dd8d8d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h110f9670ad8e99baa555073003c04d2372dca55da56ca65e9eca6c30f948174b3bd93e92d10122ebda27b7ca72324aceb0a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56160949210d67af31c4467c7df28d890c8cf60fa805b9bddd37edfada327cc26a8aa327bac56987806d05d8ce3d563f898e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h544d1a4e7b3e9c0274a844cd45ac9ca4becb689801be8c9e109d1511ebe7e0045b2ce912276d946929121d013e7419e190b5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53138653542aa8ab62b3cda517edd0b4a7910dfba668167b5775b1634e04696cd8ed3d4856b1f90911a203de193c11abb677;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb0c3022148c1e8ca429e33c6a82956677b6924c4feaf219cfa1abd2a99bf21a19fa8d6440e35214855cc1d2977c40f622d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha9bbe0ab073e3b0b80742bfe03bde92b5974640def13f7d7c107b8e2104c18bf9ed82c5112426305efa57ed058adf2233b1a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8587be9d2a8ef72bced3138a9c60a09c85ab2b5257463ef8dedbd39ac47d96a54cecc576790244f8f426f83aca8dae1e0a1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5117daad440a90a53eea38d9bbfe2d751fb56bddd76cce8bfe6de7e433c08d88d1d1cf27c7d4360fbd285ab70021f6711d7c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7a0c958165339ea72b72d0ce9bce928336352d760428fe88279ed526f3d46e3c79b4f49d47b1387561ad8cdbbf4de73ed4ff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bbb6b11c5924789e2817dd625e7ffe5361b51d81fc3c46774819ce1ecdf068a52c25ab413c811a0a85170f7204b5ec63015;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc339c6b3a77c97a7e90379e2a077fc9b5a72485ad3967dd94bafa4399af296733914666053d06a35766d199e4b8b47a2bc00;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61f3d04d3ba86d4ab8f886965de5bb88318c477370feca6b1bb8a1cdfd2e81db74e5a60933f8b9399bdbfddb24131098216f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h17256793f953e4cf6e3f104860c48e6a8dd45346fce9a07dff4003adc66927ce89056e6d8247b6fde1e0c35c93f39de222e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a6ab0ef89b51417a24f38987e46adb8710336c31ab9c5f426df0e0a738c69c0f2806d75848096af616b8438b134141d6019;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h25d61d35b7fea8f89bd9e796f66672fa467915b2435957bfd0fdf97fbe0759fbed3e5d69db36efc82899240cf5be2a1c3f1a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5f17e96ec9d77177f294558d5cbb22d09bbd07d47abe19abc679201bfbc95fcdc5b5276dee241741e8dce7cfc7be7914019a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf70a399c5a9bb94eb17a90447d8982ca372c0324f0667d3ffbf23d3a23b75e845c447ca64ceb11b4b11307a26ee99dd7c51a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26b73fc1927e68b5ac9df7e65d98a956c45e548137f78a5bff543b818d0684465021982809b3b477a5466aeedd3a72659563;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4dafa75d69c73b47c02243a895f7f1c425c9e3d15ffcbdb6ec1db6ee4818cc66d1894955ed690ba9b0419999ffadfcea5eb7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba55d13a5bcb0b43a06afe9e4fed1445015fa9f77ead1bf659589e0a7d516f9106c446b8003688a64fef0d424791c6d7a058;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9c29bf86a3b2be566a50107768b8abd285e7ef4b8a4b2da8ceadf55b8e5bcb04396453925d0bcfb6f2c73d001859e56ec4c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4dc83ab6b8cdc3ee8be6b423bac2df4f3dc9a440ec0b4cce370883a9976fb3a9b7f3b0ad755d3f3d321f670892d205eee4e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8da69dcfb8b81555a6e4dd5a34a5a8b246acaa7452691feab6aabd64f3e236d1624dc7c21f4d078eee01855fdfefe2c10ac4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7016b9b056f41f5498b33c4b04525c23290ef63899c55267184b953a164ae42ed73d29a5800cdb268612d68da07647ec1183;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee9e97eafeb484cd4ccf3967fe07a99a6b91ace537841488e8c69ccd7f13dd9e187b35f53ddd1a82e1f9b1ddf99425924846;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha45de4207280f0dc559fa5ad86376cb39d34404eeb29b74557904e2c768d62f6bd36f81cfd15d27952c7a9686ed8883d6293;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2cc90a85c108cbec6e89d7a9fe5f27774ca9863303f322da1df93f74dcec6bdc891bf99fdd8489dcc56192ac4b6ea45b0042;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7553d6286970adc105408e2f97ba79b1001460aa95c2fed651e3565bc4368ab58009140ee51acc777077177a757fbb51e29;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h18fd160c7ea834d69855e28764192e0a13b649eb8b7593daeaee1afb20216091e8a3b53b824b19b22675bdee5d13996d111;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2a34c0e2a8c25c6cc78d013cbdec431522ab3d4cbe8e3f9ba5d188fb921c7a69e1f11c83c68f61332a29cb994a6f12118d2b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b880a6d204ca9dec3ac82966991b586cc663f1216b9dfa11566d8eca21d609843fb5d521260cfb362e01ff9d1ce204b5245;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h86c08ee9467652494296631e60e0848027e0ab5edfa08b03c7a8d6766449bd8918596a68f81eee310c3683b323a1b395190;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h274364ef10b315293a17cd0288a53cb6d65bccbb033ea379e9fa10dd72d721a9b4b138aa837e2bd7301d504564fa3a4c6a5c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcd2b92d21d3010c9e1c8728bda0565d057b8ae8238e47e4343c985ee008fdbeede73b9e3753a297065ee7e74db29365077fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbbe3b7b7dfd3b5efd120d4afad47a76ba35974a336404fb675acb99189cb5c76e535fd95ec67055f245569932a9343b0cb3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h311d4c4ed17b83649226f3e65c50e59425ea742eaf02c705f666e5695ffa26a730de65b60fd68ad4ccea2637e7140e12da54;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd482290fb979bae912c9eafabbba6daf4bf22660775e226297a13142c8ac8d0b2606713c866dba3e1eb1733e271af3e8bcee;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h69e5ce758b24abfe6a815ece732b12000f59decacb69ea59332ebfbed34668f6a71b18ea5b954fc90460ee5234a8ee68b50b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h35f8024b5c80e49c61d666eac30ce69a25d99bb4ca5657ad11e7cc56940b54042df220bad1f85710fd1ea2ac0fb04abe9792;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h88d9bc12cb30dd7f9d4a93dcccd17eda2dcdd5207aed8c45c4527c6593aa283daa8c46ee4199cdc43e83a1e8bffcb2fab3ef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3e18a7f6e4e20a2d68ba5db8ec7f2b1f9e070c3e0500bcfec104cb3dade72ee7879f56777603b6d93d1fa6418faf07b6e700;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdfda64e8ad714968d49637c176f726154e007dce66999c091d545d5cbbca23c2059fbefc7164280b9ac9d92934885bcf57e1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hce30b6aba83f5201250e102f886518382e3369bb9495b793a7e9db64ca98fbfeb6fc7958296a47cc1b1c471747c0ca3f5c8f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b4f1b7cadccb68172f4773a76cb3044466c9322aaaa25e9a79d99559f14e919c4c03bce36c5de3294f79c85cbf986dfe206;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb2b9d3cf55215bcb74b5afdab47dc5fd9220fa41f15627630e5e43e44d7472c552710b32a7de674a9f1d3a207bcd5443784;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9da7329ac0542f6a1bc9a21041b938dd9d3fbf64b5b9b5e867f52953d5bba701f81e6ea80a4e7f8cc89ce8f92a305f4578dd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2265550e668ee7ee6705a3a8af98834034f20219b84dc3bd4f9421a40d07d6caeb89508fed6c24757903da2b0838b1692ef0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc219b4bb797412c21077709556006b4699e78ea6ede9e371906720f6968726adcb16b4f23c2033c827aa274301ad66e8f4f0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb4039c5d07febfd67fe1ab1403b71e33d9816f6450e21092deedcc2b6e32e12a406217389d132f6edb2cc12a8b5a9802a7a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdd02461706f9afa5ca39744b276daf60b5f266ed5f1b170285e6ed3bd9e4e0cc3f8f80e8265ed4976656e92e8a1f79096106;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7f1ab6323872ea81160ef3d74986bd6a18e4bd222521ae6fd803a135706ddd552a06ae9218109ca7aca633e07a958ebd44e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h94eae091654803fa59cdce98dda4ece7c2cdb9ecc6dfbad259828612a8e77da85cf4d9fa772298bfdff28d6fc7d40b73e327;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h6c9fe9d0660ee90aa71810a9c23d8fa84920d0b0b561bb73a15d6c20e8e0f790edc6356f971433be4eb5cb40886994d4a3e2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e6078e1d11709f77043cbd93d11e5d74a1de367d5d125e99a97f72af0b196a1a5e5b3c04f4239bf2b16d2af69ad7ed2f802;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha77d99b92d2e6769d651769cf80ffa2e31a6f410c22f26798920f22f47e8bf4a430fcf114be9895cc10fc9744414122fc6ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4493b095273fe96fb206ae4cc7ce46ecdc93adb66d5ba1df21f998e6cb26f091f75af31ee89fab12c2a8f55ee40afab38a5b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9f0cfe20df725d67698a37da7190b30f05c63fb1ee09a2d80e77597fd66ceda633c7156e2dc4b86f8ca6d55a5548f024d547;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h217f87053f655466bb8b3fe6f71829195e199ced98dd562c8b6b27039f2683ee69106c9fa53b9f20afba2c2c9c42c3c4379;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h31c7720c98b2426172f34b39db66db17e0295e219d7cb843f2187ed03b6174ca1d48099dac78a5d3ab9d4326c1ab77cc80ac;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e34c6c1ba350f942aa1c75239214fd54020ce560cdd9bf86620067324020bb7136770eba407a8d98910a961de90c049d396;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb317b85fe2c0c460db7f2d64f0d2cad9ddfeb8303d9534e1f4b3b44e959e0b5277b243eb072b5b8fd72ba2ac9180f4f7d30f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8df7c8852e20dbf2b6fddbb377c1fb8b6800792cdd5dc3c9c21633a4b4a2f2a29b7164af728f171dd02fbf501fe556fb9ca3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc3f7fc812d14e7cbf00aacb146eafcd054318bc0317589dcbe20b452ef6e0c20a835e7be4929598d3d6497c96b4a177170f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb7a89aac25fccdedcdb545365954686dcc9707d7eaa49dac5939c1cb641d16267ceea3887ad96c517b98f1027c7193a5513;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he507e115164d771aa96912f5cde4907f9f4c6ecfe58fb166e748807a8597c295351306a1a31715e1ff4791d4f82d97cae2b9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4fd29360aa6b71c1a6ab1409e477d8a6ccb9bbfc779f28763fa2382ed057aed0dff1564d75640f29cf9eb3aa661fcb6de4d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66bf2f5504715a1f225e66d99ba962cd3d51a2057dba6cc35451263dbb1997439cbd3fab7d3a008c266141a6af8cbaee6629;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8f5a655eb82ca1a6f8a87cd97ef677b3230c2503445b2b2f85d0f73a00f735f8a0d99c0feeabcf5318ffd134cdb6821bd431;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf8f59ae5f82d6bf236bcf5155da75018e8036d166bd39e7ad786552220bb04ba3d74321c0b9fdb09d93a3f1b8ef23f9dfb5c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1247bb889c6841b0e5b69e9e433f7ec9d7e39dc989529c90f4568fbfc88cb21192491c9736353b9fce242313c88bb0f97ee3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b922579043fbfb37edec09ce577f7265b2f96af6ba6ee339d15cc60de5153c6045d9e0ebf4f7864953b2150473644c37173;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9eca77d84dbd2a0438bb22492846af7a776c8dd662decb9c74b76646b288d93460a0ceda7d88947cc75a6e0fc91ef478b2a2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h283cb0c24f6c43e11997ef59aa3cbbc2452659c14ebe9ea221c5ad749b1210f3a03f2791883a1b43cfadc1e4984a94626a53;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7fe4131d0076eb51703cef5295c9e568795c8973b1fbea1b4ee28b7d223b4c278b9562594027c396617b3995f49a5f6e85d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h360a80bcb20a8cda74dcd4c05c698fa1a321dfef60ee1af6b7ffb0cb3f1ce9527587df12ba5e9ba693532d3ce098d0ecb98a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha754494f2cdece38f62d2458032e4f3022ff823e5784a1397320bb4e251768dfa9ff94a7e6256aa8b54583d8b05ebb4d74ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc06b990ec78d0d3ce9ab3c5d59ae0f6c999538c1c8911dc3789b8acd5a24209ca5c0f7f583e29a3388375cab29fa123904bf;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd3aea7c1525c261e657436c1048c63acc06d1139157b608edce9283a6924cd6a6f7b10b69832d1debaab63af2b25524cb863;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f91e8ada2551d69e09a6cd95f7f240257088df00d3af91f2b8253a2f0010b15b196a10f537417f5ce5dbf08da4eef37fd3c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9aeabad5f832f8a0ca4a0981035800e2c2a57e30783d983138459455942a4550ee18b5f1d8a459cffcafa6f296585130d023;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb80a4c4ce4eae449e97126d0b6cda09b90bbae6cc3e709bae3e7aa339ece00a2f1e434565cc2510814d77fa40ad75b4692a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7c30b148b00a991fc03e5571f66c790a3ed9e20399dad250f4a9629c2d1fc4ef77b8e7944a1ac0a94904d4d5a0254946644;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h58860700e46addda4fb9342052af963c92ebf19bcf23445d18cb64e8211d21399e58d4b840a2ed969081863ec14357a95d15;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7a7b44dfd9f5c1a3ff2ebbeded781b6cfc5de3ed98cf8fab3618eee2b35ae954e8b07dbe9ce4dd14bb101149a5c709ab5c8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfe329635e5b8a0cb9770d5c0f0fbb593012402f6be1d7de6b94d5ed605f938df238ffd4a38df5689dd223e381e5a27b81946;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4f9b4ceaa638393511bb5fc538d46850fb10ecbb959f79daea35484d015ef20e1fa76792f318db9a8e45ba688d963017a5b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3a89b644ae62bcd6fbdf61bd240debf09aaff2430347e8f1627045c9cd242961cda52d06544c75c0de20f3fdc6fd9767de7c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b160ae0fb1202db89a334c37e9c2ee3fde4f71982489250a4e989f734815361db2417950c66d85557aa8c1a3af367088a4d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h53596279e4ce351f21721ca4348dde54cb550e26c9b97c15eb69feb6c6c0bfb69c534ffecb1842a4e27b934b8aad0313d7e8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h66600249e56bf1bdfd47147135f37caaf6b678c62fff6a05550e89a5a584f87fba377a9df5cf23e90c93b37988932dbc0b5d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e7a98b77f9a2f9cbfe7c82ea3472ecc083a03fd510b330adaa3466a22feb54b9a3eeea65dae62112ff32da3da48e474f6d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf4ce54bb3fc22d2baf7d4fedd372c1db3b0e9576b4fdcdce166e32e4b5492430d3353c339d82e53ebdd9400d97ae8e82a736;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha1b4217ab136faafa6cf14104360fc60ee94a5ae68a455b5e0cc48edf04fdb7f004bddb1459c72c88311723d67093a942e24;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h178955d80d847186c09c58e15755172b602940345530daacab63e299a0cef97c3eecd0b0a1ac8a070ecc52a8d1eb0dd7878b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heee3b354897b82725dd7787d6bd1da2b12352073f641143ea475011890472351114a008b97a817168ed20cca6984a58df486;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82898c9c3751620264c5694403e0ab8f64e61490792b2971c4431a907f5a2b4ed9dad5a4a88c19badad5e6fd999e64c2b4a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfee67a8db99c7b02a3e910861b3a8d039de96c760e353efb92d84ac1480c7e7b6aba68717ce4d2023d18f0e5265dacd73fa;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc614929d23ba161411c8720bd98f8887493b1b6266b957ae226fd93d873e72db974d9736c50f967263a310c5d38cca8b18a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9d23c42738f1078fb4798ade02b11b725c0268fdc8ab9e9f31be88a7be58838b46a2b765ec834e4eec69d3b8317063c0530;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2387a7b891de8cdb98d4d6bdbc760625c97c1e0a12887e98600c286923c77d97d63833b318686de6860abd2ddc66b9ded6ce;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc13cc427a1aa2fb6cc6273d36d81ee6dba417a5ac8e8b79ecf8f6cb6bb29c19baa891105a0eb96cccc0b48d05f7dacd11db;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12365583a27e6ef0f2bd7c17037415fea2257ff74b30e56dc2eca777b753724e981a7acf74d039f8b605030d0773f308c445;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9ff8d2e96a035716e3ffaea92f87d6b7f595263f5b55021251296adec167e670ff22c5bcfa6f85b4f145910126e60c9a3634;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf6f2e690b6009090d1c53be8f761a375e94cbff8daec3781c217f67a49d8a6d208f1f18733638553b10965fef066bbdbed14;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3708ab9ed8071e8f764559b4112b03ccef7ff215b31814a2810fedfc1e00f5dee57e06c7410089d210d246bf49290edd895;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee57c4c600598feee8e1b42b3fce7c9d34d04329e38217b40a6caec3fa0d447ac141a0d9d98234fba39ed407690b0d5c4887;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he30175e48c4337209224ebf237228f86028d2b3b19ac419b59e223abd07659a2cd11e689997928534d859d89f6e78e9e9f8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc316b4c6fcc62db0a351191b1fa93c4379a342713aacf1cc18ac1815d348dd51a7b8c0bd3f090bda39734136ddc71ee661ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1d11fceccb94eecff4c9b2a0e4c16e8fdd132f285d810210f06669aca9c167189fe99cac2edf0872c80fb6e1c25a620d0823;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc504ca0e77dc98ebe7987126614b003166fa8b5a4f53a849fb058ea65345e9be69ea0126019dc54a9e64677425b4363acc74;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h365b0b1be55bbb0d1876e3cdd2216a28d8f48264bbc6021ea8b1f59fa05c4a0114a3901c68674b1cc46260e47627c034cfbc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52b9a9ec22c556d2c51ec1191b83b4677a840f5538374704958e4075e8d3338ed7e9df0d9d636ef64baf4af89ae4d2382aec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h529f0b94f4a1fee67e4379a3bca238dafb4b2e0d36105d3a0882a22a652409943aebcdc36ae40bb97c2701dadf511a51d2db;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'heaf64958d3741c98b3974ee153e2716fb6b620274861662766bb00db1dd59a579a304228c764ab67ec96c8c5830a4c73c14e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf09b03cbae2d1cf6eae57bfdfb78b4ba775625babca94e5897854da32a9d32d2d89abef3792517bee7f2f03ebbb7f870c2b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2755f76c05f7c5f5b4244ad8d89e6acaa7231542207af5bdb4a96dfe76a12d8ddcc6a17232ff785c5637641cc9655c3e715f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haa0e812f8c4d0d62a7e69e5b72b0476c33f84ae74bfe223dbb068f4b44d4c994034fdaf32142a572c5b54fe6962b5a92b8a0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had1b734f3753915684f155396ed7072c12d5afcd6933f3682618206ea956b31783c54803a85f6f2b9bd5bb47766466725200;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1bd8928259305f4b5a7603de86f8a140b7c91787143877ebffd26391fe7da07b2a249ec29831770f9f1ec3966c817631666b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5088519c7387cd3f6eedb797ffd89ab090e541c8ab65e350db569445c0536a6d51828223e856453e9f6b46c1a72774a52d37;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34b9f938eff7029f2f92ab417c261d35391c029659c00e5ac81ec51cd0ccc2cb797323d5d19b2d57e26b42fbf0f7a51beaf4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0ecaf6f558f8f8f1eb011c1ebdb1132fb8c2bb167018db05244daf8bf34f7aa99bb986625836f3b1ff3036ee9aa78f4a7b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbb8530f664d01e70b208b3831eac5f465eff49285f20aef4282511e58e84e975749882926913b4e4467cfca17507a8759803;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc339324d5567bbb75045dc225a586e07edfa315a6500825304d00493e123a3a59854acee9c3e91c40fe74f6fcae2270c5160;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h32c15e4d61ab4de8418ebe52450f549318e19186d870b2fb00ebc4a5ee7df80358728f4cb90be1da18a8b2f397fa6ff271b7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a04f016958663f200393d6c1d991f0b6988531276e3d98ca47564114af7c3d24a3fe7fde0c2691a13a7e6ce9c511efee917;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h26a2ddff05ed3be46be2ca8fd7f0f83e31a3c311daf11686740f29dca684fcb226886713090922adc1728c1e440012bc22d8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4076a513208c74332c0328c671e75bbe24887bcb9423b9a70b9a4b96f889b38cb4b892684c24e0e34bc63c2620c6313ad30a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbec5f301ccf3c5aa37fb452e0aa457c45825741e4056d57437381801c305f8ce49327db9ab0268096e7e00d694ec1139a57f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ccfec70f3efae364e466e73f1f2a2949e8c5ef0d0eabfb2f4b2e822c020bf3bb50e46d978f86dbb60d890c9cb21b82f8aa9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfb75f46e6452009838de8df24dd8a1932ce5d09d0df952815d4c6f01ca10ee36fbed82ecf5c8e81088f6efaef822a8678c11;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb09164b4a33775fd4240ecaa0a5c8b1551b6687bdd1df9268d2b611d4692c892ef56340e5ad45624005f9c1790682111e06;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99c830827178677a6f4b8a5a95d3c53a22e0f7f252fc6655363558b89cc734d965843cc939b9c6aecaf047ab55b3204ab343;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8c395a6d6a8a6627c85d634ad557cb343e48bfeb43529337d15a3880018baf139e7580e99dd66a86fa0c2419a6930036313;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h97dee22e3e3c63a039bbf40dd2b4f5d8f1c5c91a2575e55d902acf84ac57f9103fc2649186efd3d278c724e824850d806fd8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3d8a4f2212d5248490f26973e18d8d0ca5cb2b2e5270ddf362922f75832bf5cc239818edf435aaade5ddc5a198d07e34a3d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcfe588930a8469fceaa06af6963e71f7f17bdf8151165b5dd3f2caa4a3fc5ba53e417a998fa88371774c9aab8e6fcdd212b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h34fda9d67577d4def4b8b91a0c3077367d116ebff3c9d3e378ef514cae96fa2a951fadfc64e8024d903cfd296f3f40e6a867;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2cb82165bdf30f59c594320db91f8a3610b8b07ab3322279337300f97a8a034f7159c2f352daca3b307d28e49e0758b07731;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7be6b4a58d47922d42dd38702787008b6a7fc4d8e5e2a160bcc29ebe35d09210acbb03ee314fdce80b4e23dac1835de87817;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h485de3ea478f9561affbe8d8ab02d080129542cd775425be6fa49441e873dd8eb0c7758f456f87a2d7051dedcb3f07691596;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h633f9b6fc258b63ec00369024bedbf3eab39b0db2acd1e342ac1d6da3c8c979e8513bd33f6499006b59fc1b3b9e686f3a71;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he28b3beee13ece1a2617d76ac5dbf1c37c2038a79d01052c6672a5f29b45a36972c82bf02c7c88d6630fc5114cde3fdd569e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h138521912ee22c52b56d616bb8dca8b312c53d9644b273d7d6833973e0728283e60227bae76d1fff061d50448c591a76caa8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdddbdeba68c1459c0cfa18c48f3b024ac6bacb1ef98c386fc4f5781bb62cca68b8743be2eaa4161224a0fc6985d380fcd4dc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha91e334e6bf982133660a45973ae3dc1a4aa60902c242a3caba0e441f95f60eca55150e8b2a7170fffa515f3be6c870d602d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45ecdd178651b3863d6166f937343e9f040f7852558aa016ce21ea1ad6ea9d5e789f435bf48ca12075246d546d08ce335eb8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h52e75c0b058b1afb33cd248e050eb75f5297ede14025a4f8a9e06ff8d85e13e79082042327976c876c1c076299695ecc1899;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h13e873667895da91d84feac4af2a47842b64750fb1139800f09fb7384ad371525a464994a0a809d7f5b8a4182810f1068fb8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h659cbc5dcce0c40692395e57b5430c67630fd76152f4baa16f16f6cbed86f87bae7588fab0c840e18c947bdfcdb5e2052c31;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b0feb4ce481d9f6118ea71c7a4e191bdd65ed90e41cdc6a32211e04a962b852dd447b347964d03410a5295b237982f1ec42;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9e8f4c031ad416e7db05efaa9d2e3e10f57ca3633ef4551554044612222fbc8ac7c95baafeccfb6a8773a2a15ebc6a1c40ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdb917397398259af08ff092a919a941183c5581eb87f369867b647bb01249288106004376ca22830b255e8a230f51da7ed8b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd9f09723db9bb565589f738573cc26520b40105fcc875899467b6c3f77015674c517e6a10166cd48686d9df339548b0a83af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a8da12a6ca680b6448330fd0d6b94082b5769f486c4ce210e2dadc1dffe14fce14cd142c104db9f83892b64a85df263b978;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e96dfb6310db8dd29dd99e8d5db08393a0d738cf64753a11547dee6b73367920318fd0907767f24bb5f867be837ae1892df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcfac340eac906f6b2cfd4c5ca10638267c0d31cdd86cf85312ad14f70639f33150f323b0d347cd4b0af2aa6c77977ec7d36c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8690983f87a8b2380bfff4b8bb5150e2a5e38eb1f3ecf1a1b23eb0fb99f2e569167ff74907c6b901f73fbeb26118bac5740a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha751a1ad33d52dcee06fe1e2c5bd401e8df0b2c7175ebbc051eed7c5de261c96058cbad34f34466b7cbda71bda6b47431b4b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hdc09a1cd49db448584494a6209bdc9f8f627af7eefc45acdf98e35a28b439c83ba78ff2e34a5d84a302cabde8c4c01903ba8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha6e747df93ebd5e7ca6be04143348d02fa5236e9fddb620366f64e97a71f52753970b632bb57c2deb3559b47ace4684887e6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd0720e06d3f26cc47ad895e6a4c2f987fe53f89d699729a47e079447e80c39d19d7ca22f4c98734768b047532c2c3943420e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65a5894749646eca4cbc8c3d206a8af6b1f64d52d05ef87f13f5aa08efff65854f4e666b73f9ca8f2fe649a2c026ed5ea70a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c870cae42057de0d0db291f1ba839c439c7739ea54f24bb083a56cef21da60a2ebe2fc9a16c7bbfc75386a958fb2405fc66;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he8c7371444cd10d6b4a08056070afb612509fe7c1c6b3947c47d07159c2120b1bfe7df2f353223c48ea9b5dd09ecc0aeb035;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc315b532ecd72ccadb5d3f8c6cae7cfa601f3e64e5962bfd9d908bcc98e52d46e5124a35a933c5c54bd779a5e9a217cdff3c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h65b8846d99a687c17f5071d5a51f83e4b5cc1f71db1fcfd3b46b66aa87966cb3fcc3b4d2a1799936ced570ec6fa15d6419c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2935fce4f77a9abb4476003ea51932432b98b28538282fbfc3a1c3b6309a4ae842f28be247ed859f6c56f2593a3dfaa18c13;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h885e3a7351a91f0083e634a0ae43641aefc5071b5a3f73612f4069dbd762bd5ac13f1bb7e64ec0aceea59f2cf54605f0efda;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h70c605bea27cca05d11c03064486786b71c472eb3a84a3753a5fea75e851c482845c6da64f6a9d38ba8a6edc172c68f7bed1;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h521ac23296dd2a7d65a992ebd24202ecc37cfa01b6378e8b286cab2f52633aba8f728fafc577911ca3ab778c863da3cfab97;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hcf06d2d28caca0dd2fbce36a57831d6fcbb01cf6a721fab6602970df04aa04021f69bc28d18d91fd145a90d60e2a83bc39a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a159b54133f102c64bdd1c928d945db3909bcc5071daaa67aac0d628bafda94271702d5034f501394adf8330648af59e34b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc1c936db8cdb3c27535e08a92cbf9b36cee52320871c3fd0fcfd9920b02646d65947ea105c99cdcc90fbd84c58374da067e4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h12e45cfb526ae725e7d8f3fc107c884c7f833e7a21686014e07a188a2998e3a83a43393405f10dc93a0576cf92544b18d3d5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf9e896edd1945574e15814ddf10ce14e5d2a138f9bac4a9ee5a7aa30e57d6e1b6062a1587294614a48fbeeeee6650ccbe753;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hba9152d9c38971e4b2c4d7379684aead574cbd9aecc71040f7f1dd3abf293cc42452d01657fb0d8cede0af251c9c6c14a63;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbc0ab7cad2f1edaac83ed6d316ff9dae11c3fb92744f220b426744c37daad04f911d263308821c228efb11bc8a23c756f165;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha982992472a3e5a5ac95f5a75ea9a740196170fcbb023cf4cb223e197027b604db1cbd739473039c50b7758db3a23a9b65c0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d252719c4b4630468f769c4ebfa0ac73276ea82e0021968d261957e037c1b5ff4d1ea0560e00dbfeff26f5c609dffaea7df;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1f08cccf143c23a9d8bcc8050218ca190240d3c52c847040474b92a80a26f16cb91dfe07d761ba6e3c8026c4bb79dd80ef8b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf06486037dfb809194d806427d2e58400b3afd7b6b743ab173dbd082f8a37dff80e986aa5fbc502b5427580c6cac7e16a4ba;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h56263cf5c8f76381607cf2353ad98c8b0e4bdd0ffaafa126533d56a808abff2728361d87e53f821fb07ba8509083cfe3d60a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57b21d84e9c01fcde50424c7e942eaf4c1a29dcc23c995ab392b42ccaeed4cfcd353dcfa695a611bd001c42405b5d7474bbe;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc4695f3cd856fb2d706cddedbf4d83e612ad8e55db72676b3425f941084255efbb95f4f410a9a27833b2b2fb6cdeb4f3d792;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1a235a24bc0ef470472fe13bd18853741b03eb7200addfefdb15cd8fcb1b1901ded10ed2b59ae780973ed4c2eac8c14c77f7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf0f06120a226c9eccdee062ee4a45c2fd62d10d7461ac6605de014e4cc7b3e8b992b2346919a524e8258675a1274ee9bcacb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2977b7f9157112db04d00df145d302d2a02bf2620f201fdf597254382f3bc9d29b87715b41fdaa92cace2eadacb084363318;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h82b17bc5ab24f751aa89da651b1d0e52e278f9a96a800977b6289c972b5ba3fa9ef4eede8e9c69615e855279221b3f692b8f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf2053b802021a37c2cf3a87780834d846a399d33ac33a426ef2d21d5192995ff1ce178be730ca88e62f39c7602f72ff7245d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he7347fdfc320a9a033622f43c587fa65b0fcb617f555dada729386811b434b6ed9f715191b8d3a0fd0129f556ab3fb6937bd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb29d2736ae8612ede3929a9b2f0b9ac27821bf69835f42a2e86317690abda05697f559b18f787a4e77feb14195f975b30f20;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h91b6c181841c74e3bb7d4c5bce097e67d97714d4bd178e839a850f79e976146b555e3149e80212c5e5eddeac489e14d9bb0d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h240ff4e7933b48dd0ef80b9dd5687e81c3f03243a99a6223fef435ce7949a1871b4ec7cd651dd1fb8d7e0b11901a1cc54c52;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95060862874ebb154b8b20413f1fa7705ffcb7344285482ec180146af0c28f73d3b67d39abfc3376953a35822b8aac9dd197;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfee51956213a98423afcade4507f4854d62885bf35fc0addeb5b9395b04d26f255e4ab6ad24defc71c1d544d5b43797d4675;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h38d9fee1124ebc1ddef879ca55958136568279c047de6e7789cf038871131ee034d88377e83cebfe741a8bc85286b9fc89d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5896f2315466be01a74015cfbb7c99933e8cadf1adc9216949ab2cfe0d20fc8f5e17727aade8e0ef83e9fd5b57dd7367770a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd11d85d4703ba8c65fd959d1a3ca20ff80375fb9485ab01fc697fc3227ed35114bdc5bf9c6e71d39743262a5522e0f0c3cf6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd23e6193001af8050e9afeba37dd16bfc83cf7a8a6e75169c52da3437755660bedf09b19d7fe49aba82a7c00848315ecbd64;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4c9e5a7b6e3a8c8fb0cc84c4a6d629a33b13ca539cedbc6b5d181d5207b8fdf87d9f743c98be217674333d5fb5fbd979f8cc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h202c95d7283307cd6e54a4d9eeb1c6a3905675c41d0d25f831bad3f7679a5330342ec54d692529d8897a9845d2b5010605fb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8224d62e5882d7bdcc52465e68bb4f86065a01e57b3ad11d71736420c2125ec5d523c392d53d3307e27344ae6278c5bc9fe0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h346926f15708aafbae446c0b3d686eadbfa8f5be33aa271111b6468938d0305e64582391781aca1ff3850d865ce0e72d47cd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hffdd25133d7a586eccc43f6ea7c2593f815c80b89c216f695bd3b10f8b8d6d481023553e14d1bef2f54ef8935fb8310825f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h36949f2a4a2c70a1b54afc8532e302aa0a23f503b7010cff9fe123a55b1453266d6a9e5c8a2c0065be70c07b98b00f7b4494;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef504328340b04427eb38301148ab7aa16da99b71ae21666107e8e394f0641e598b84f88c6826939f238a8eaae4d3af15a02;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1865413f7dc015afb9c7e81f553367d91649912fa83c11a496931f80c1670075cc993f799b75174dcb6801f2e57dc47d2aed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h61cd1915464d5007141bdfc71beb45b034872e4631c1faf0d56094b669ae9bab9b85b0fa91de57ff38a1a7ec89f46742ccef;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h67854003cbea7fd370fb189932230f0e470417a6769282a41545aa3d566e3e46f80c0e77cb1c2116be38e206076cb0fb3fbb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he329ceded2e93148765347d0f76c164ea4146cede669082d400df549ce4f67602f8afa0d23a0495ba7e4f8b16d3095d1c446;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h410e10513b6f07d09691a8519a3bb63ab768a41ba81f03149fc5a4fc5bf25e2a738c7f9f89dab1d617f07cd73d4c1f48214e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h268aa0ac497ce8b02ad7f8ba05a8d274ffa9a9ede4cda7d23f0433d76c4322533f39a9a23290e48de901f9b86853872fd844;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h494779eb54e50870f2c6d933ae9e182bdb5aa10d62e42285f97973d8dbf70a440cdd6ef7b3d100726c9a4ba388aa1447f4e7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7b4e9fdf7d0e6fafa7c6f7623bc1c0e96baee45bdaca87a62c0e18c17d667cb526e4a75cf4d5f0d25b14c70562d9f1056802;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb3f848da42ccdf8e65a6d9f68221327909a097d2652862b9ba3ff114f88504a334aaff1221359ad77cdc5db8a2076061a411;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h98484a82c27a7e6efe5f0c96f27ca253d3c7e50d2f1dc0ad0c05051ffe16e1b924299d6dadf10bea4fcf4d7eab1caf309205;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb44838aca872c1122a15452976976ee4896b73157edffbbfb1780343066e5296bce2b1ee1f4813378ba4e34191b43a99dde8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he007da8e12a69a36b541054e0d8947c5877a4ae7e59a236a285cc5a0910e0b59a17f511891cd3e25567f31164c81fcb2075f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha18f7921edd40c549e9db0cd432f4b3c58076d88c7a9d7e3d5b626ae71fa9c39709bc979af51a13fdb72375ab87f137d0000;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3d71bc8edd37315f7904abff229986e95468c470ad62922e1373e4173ec4f23bd758e6b2f590ca53d3324bf1082872707f2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h506e63f8ceb6f6a80406c648aafdf2597d2604edd5bb2545dd4efe7fcc6eaa23289d8a5bf3636be896aa0bbca9e1dff12b33;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h843197fda4178176caef9e443ebe8c58c548e3446ee30b52dedbed26eef986fbba3e4c9cfd0f19bacc3b7f60a0f22bed98ed;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5c918e0920967126a7f09085754206d3080a703f5b79edb4e51c1ae8d59c82b506df0c1bde0098781f25fd2cdc386aa6ab40;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h883ff6ea5ffbb6591a98f76697d8c219aa6d1d78f977c3768790a96609d86eec56ff03bb939ad0336453a9e6dad7ad704c15;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1c07c245caaf6db2ea403dab8c93e3daeaaf36795e2d37d687d3e0fb7b376819d25e20baedf2ef3f78a5bed07f93bf16dc2a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1b096d4d73a7191e8decbb1499a0de8d139f3af5ba7a651d28c3c7503f50639baa76069d2e5ad1b1c2d781b2cd5e9f3e2af;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h112cd07a01ff24f24756cdcdf40670f1c9f9e324268a04ed9acb010d5fe14436358d79c461a857aa69c913ec3d5c1e83404;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h77ae5c7c8dd17251223f5b529fb41562297bc62db38e1ca09c63dba006853e3fff531e001b4e51f5b6a718ebccab39b038dd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbefba7a8ed96e22fe0baae06bbfb2ef935eae590fa696af0edc1bbc4e91c4bfcbadc242eefb145cfc85bba8091a1a45a7f16;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5a8f45b6d9b486c7e917588a29923ebe61bf3f309bf73105ea02d35825a1236bf6556b32f722e83a765e8e600f2a943d37a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h863b04613cfe605ad87b50574141f803fac59bef013e8485005c99f7603e218ebe25bbf12f73f1896f1cb5844537108658e4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2f3f143d3fac1ea190d2562ebf974b9e74e990d54a85a157247e42c6acd16526a7f5e0c3618aadd1fdd11f25f111676ce518;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd5cd6bd61eaba64dda373c6f7c8b54fc510a70d961eccdfebd010b0903398d18d209a9b8c8f22f69bd9a6aad0a6227036664;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hca554ce081f74212c7f0aff0af572d5fabd9f8f2c4258640a1001d21fd49cb146eb2fae30583953067e39b16937004356050;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h926ba0038e4c23bae35e51eaa6706b0b60120092701adebb1419722433dc368bab31fea9bc3fab009763b013d8869f084d03;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5348dc7d1577a57e60d4ddbc7595edcf1ce42b28e5f92bc3aecb2e71f18b0dd2deec1aa4a5f2828c7fa3a1e090914dba4c9a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf5ed389f18ace21c5f6bd02a75382016427090603685a6bd4524d4734efc7a9064c2ad37616ea19f114058bc4841afc6afd2;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h578268015bd38b44f9c4136c07cf3e5fe7dcb1465af878b57fee3d2058459cd8aa5d17163e799b8c20ba34c58de72505c2db;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9d9a29f199389a25b624cb31648bc1db6f6eba13d6f57c66c89575e354bb7ed5aba707996f67ba73cb2eec007f9dff667dd3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb2ee9718264c4e2ce4b0bb6c8cecdca81301f591ded8676d4ef41782c3fd01b035e20c732dfbfa0f11d96aa69ffb9555c54d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h50cac81da09bd3410d06a6154bf33b60bc125427292e41cbbaf5bbc158ec406de2a0a3dd480ee497f59a3ef9b4786598965b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c89f6b515720d4ff149bb84600c72f8bf2f10167d6897438ecd3c2940009bea52558b56a0727f480cb1382e1816a4f395a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4e8736365ed3e529ce7e1eb22ab76c7bbdd9942f4a0efa5ed4b4520aa382f4494457883e68cd956565c49c9f008c91862f36;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb540e555cff6fd4e50fa7e4ec652ed4decfeceabc3fc17696b51a1ec6aff411e41cf3fa12c93d690e981746ffdc6b727db72;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf65e99725432825e6a17154666ab0074ec714f2b81eb3a38e1d2af67625fb528b7f0cc483e24a92d06eb557f14dca3aa1e1e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf1875ef1e190b68d5057187e0c357add85520e8cde1934daf6fc1b9b496e954987d1eff85026cb90bcd3a10060dbd0b92bdb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb79f3c30e6414aa33e0c9defa0946f5613120557e7dfdbc38446339473d3dc54f89aecb0c2526c4e372a205994d49aaffa59;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha5c2aed8035fb4a3c8f75211aec279daf534b54934173571c6d24d3595e25614b3040292c5dcd37d0d11acdc4dbb9ee2a4b4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb90749c3f94b7ac5451efa8e581df92dbb9d2b11b3d48d023fc3c3b8ee3b365d5058c725069aaf712b2797264bd4282ce149;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7c43d79efe731afcfd2d493f7068a24533525cc4b76e07218d5503540b31258fc65388fb950e910e91e58fcf39eb19031753;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h428287d19d163230ea2df3bdbe753cb070e5bf299924a2d412635722b4652fafd9f940a8fddc53f3d34bc9bc8e2e0f7586e6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7945ce8da1b45215423fecc43557857abdbf931a608eb1170d257ac343dd1a446c4a95fca5de5a345fe65c53fbdb495302c3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h49eaf0615bda5cffec6a7a0e614e12fcb97b06bf4c0fc20b57604361951ca0688f7b862cce98cbc1200c46dd529d4dc49d7c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he22c82399698cb4daead60dabcc0d1f7633ba7b12250d9d7a239e97a2a17801ebd96c145d349b302c5aec12978b23d59a2b7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfbf2494e89b7dbd9338fe8e7c70c439c76d29a7d719b410a74f78c92957b567d7f344e3aa7b7ead05aec6d6fc5c86f883625;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h196a5daf6fe2cf3559a6fdbb32803b4ff7bac421f8c40298ed707039dfc2dbc8cff6bed347bf304bdae383d9a5b6ca64ba9c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2e40237398873787c336264da0bb1c010d671badded7ae147690200b93621fc2623d27a33ebfde7829faff4c50097c8e367b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h301c06e2497bb22838f2168fd59f4a8e43faf1c66d8881e368c4568fa96671d64743df8f4c95587baeb0975e9012110f34d6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc8f4a8221763604491a31778696b9365882241d343b62b99bc3ae6dfe44b82d815c607d9f17cbaa12840965d3339a82154a6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h343a8da6cacacf3146b21f0c50e082166f33d34b6b6cd801b3442c62571321be86c0e02e3f4b41bc1151110dce6d39014dec;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hc58e766c7579eb0eb4aca1e5a18a89d62d76e821850b61878603b63c0b6f7356dac3960c01941c8e95206d86ba6b483ef664;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h400d44f2a50316ebe4e4fa44218f80fd054d10dff0823ad9c76687f25cc5a6d585eea0bc3f7473e413b246ac9b3136bb58be;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h92553af71242d33b368206572c923d29bbba6c679bb9d6112608d6c93b66f26b94290fc028ca4eba6413ce4c1e6acaa3169d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2c0bb56de0df9ec2db2967d85b8d5f7a63273c62fd27e89dec618bc38aec5a5795b7071cedbbcf3342cf1a05b6a3da5f1dc3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha07da74acab6d458e56cd856141bf24c9a57c35293a037fe60665aa00d7b163ecc3c1ae9137b1e8980528720bc1a4ec504f3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hfca977883129a140bc222d1fb1abf01842d4c8750471fb674f730d901a341024563926cda85cb3c3226f13961cbba1c10b1c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h55664b47ea2f93f16794b658c2cde1a32376547fb6248422865f27013afcc614afd963b685a158e195f04c94268a95f10044;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h283a7e08a4a61ab586563e4e9b77e9084b4cb8ce4b65a6e394023e0bbf7063c4c0dc0d03c1a132434b3ada3a277debd60630;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h95c16056cc0c8a542ee2b191e0ccfcf6956e4cbd6c640ee9cac7ccc78bd6c2eba33afa2a6d1aa32b23dfb53e172f933b2e6e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8ad4f7a8ee7d86db8b9b42250d1b4d48ea0e6301e0a70c9671aa164eb6584e86a9e20f4fd6cb72ba4133e6ecdcf6b0cf67b6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h80d19382bc37ba6b9c297725614e585f3a308faccc0b791fc9d57da3767d02880f91f0f6fb42282b5bd2ec29234eaf2cb199;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8651d7cc45733b3457c74dd72550c3033ed9479cd6053d8f858b37ba04351d35a3781c21878baf2f7fce085199366717f838;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h199120cdb3679495e822ae081e6e1009c1ef1808fc4684e8f62fa52216e729430f7cda9fe1e52671cac5c62c838467d0e5ff;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he41f6ff0e2820681a5ddfc7d109912c678274d6037c8f85f171ed573fa56c4a269594948399ab38940be2f63249d0804af5a;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h7dfd568863f3baf4f7d5265efea17757490e629595b7f69f042942d033ab6c82761dca95608fcb1006436c6552521bfc1cfd;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3165b51ead1a282791b31d54254b0048cca4f7d41df9cf92c519d9600a3e6e8a903bba319cf917a74b736736880aaf9c3623;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf825e9129874f7b73295bfd853bfdb0c033692e108ab89762d7fccd678f492df8f35f87c66ac5126f421846ca0a0d86ab830;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3047d8d99b69b07bf38ab6339a0b6e16db060e6a5bd8d50272212d9444b991cc11905246e67d76ae66c22bff621e97629322;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hee9f66ccb41971bb1383c1709330a84c96e6edd93bddd9d1fb5e25e087e0b55050f610b2768a37d7838cf137700458dce070;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h16ecd4da97d599e8c2ed8c6f0aa546329446827059803160cf986fb1b4aaaf4f86533ddb61b893ac7152c05fe8984c79e05e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hab9e50fdd9f4c04972c828b9b5a2977753ada180e3803fb796d1c86f3daa8e89b174ae3c184b461ad31320da589615a18510;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha3eb94e51959499ac75c3e138f34992e37b31f9200a920ba3e559770fd6e47f051345c0cc8010c133b394d01f9d4ced1d83e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h746bb2c3ad99cff6f42e90b90a6a49dd59add0a9a419d75f3fa73d46b7b8ca1151c0301f06265f96447bec83e372b96d3bcb;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf6252b9998c8e8e42bb16f161585c91f629c5acec5ee59d0fd1994ab020747def35d596fa59bafad6aa81dbc9a6e8b760a8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6a9fc192cec4afd96b3cb4b7be5ed45879740c7332a0564da97f5f99781967d760cb5729173bdbc6e81d96c362637fa1d50;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h798db40204aff388b50c4f2a5714693ca1e9807e7c6099ccf9246d6bdf3e113bcbf0bc2b3bc1f91ffd86c0e0ac91bbd386a7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha0b63017541c0aa1926fcfeb50ac78a8ee85068831011479039b51a18cd8dacb14398137760d8b8894533d5de3228c174e32;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha398d3d145715cbfde21d0aeecfcf761ae5fec0710cb081c9e94f0eb17a61da76df2716cafb5f35e42e2a11a41270532914f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha93bce2cdf8f7762a8c72aed2d8477a38ec62cd99f3342bd96c264686fce08103f3c7a83bd8c095b7735511fc1261f0eb2c4;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf007058cc73b7c7e61730980ef5ed6b084637b3dcda9c2dd9488f6098f637fe6ae7b496840fecedb4932fc48ee247b0b896f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hef668d5149364d079511ce6aee2c92e119e76d6a5913b93890d4c5227e594845205889c6508eca93aac590f9153a3a795917;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9203aaebfc4fff0381b8a33db599e6f491ca0866db09ee025091ee82e2a5f28e0671b6d69e07cc491ea3febec2af51ff14e0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h1cc04dc3fe5375ee95ddc43ad7f71d3233c3eead2d80ed9f76d9002d2c96092f54ac66e7030a9a76318253994ecfd0480f3e;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha2d67787e1557ccea774289c6487fc4f5e0d2b0eca4aa23bb44131ba1d02a35b4df3803c191e0e07a3e57a308c4990e22f87;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd6f563cf61821a796a5d3d4df94e597fc42b8d92e05eea3a14f75d751e05858530c6a1f807453735c984720ad43574d7d533;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h560b4f8b0c3c1aec78733ef0c050f584afbfcfb8b0a4cf6366ad9be9c4d7b3957c06edec97f1042731320cf341439129fc12;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4b11c2528f80c2741c487825309ed7e2413a1a47ddd85e7826118e88b4c5754e48b1bd8a373ea2f3c5b320e06894a31b9bb5;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hb5a2c28629eb13db1c927d93438b4bcc562df5c8cdae496a73648efe50c131caaa8a55916fc2303c4fb42763f0e92eb8e42b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h557ab172b6380c2048ac49869bb8598c4b5c0a09a561e9be9c24297906827e54e089b776ad6237e2de030bec84339a3d2587;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hd2519c82b0a8f83955adb92048584e9e8a71a18092b2d2b8f4439629365cd419ad4db9a4c0a89bf7a0578842aabd8936b764;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h59659537f833b468424ba504554b6fea58b60c5a75a896c015b9fb01f0b52954d0ae5d5a0f027f18f1709f7b283cb5c1e787;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4cceac9262ed5ca4c6672b21584e14a1ae20a9755af897b9ca998d51517f0f7a8408eedd4d683fccd59113e45a80e16ae5b7;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hebd4fbdf46805dd61f2378f87c7120bc1b625b530cafa5f126aa6967f53a766c047b37f6f6603a245e804f49283ab84242d0;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hf24a6ba7d76a74b4486abeb286d7c0c63ccb84cf661b6c99bb7366b9bfc7897b32b4ceb02ab2c59062b9340e5a9b17b92949;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8d0b4f5955ce98e9a7d783f6fede1d6ccf0e10941e81e386dd4706380ddf90719fe9640a0e7e142766d0db3e1cb5b51fe7e3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h4583719d49d8b02341a91b9e18463ab977cf1973c75e8aeeafe742cf4a13c63bc9024274573dfc7473c45ba9f4abb5d34819;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h93394ec778f3a2922d9f619026bed7e2135a3145663fc97817218dd59c588d31546e2da67e77265637e6ec60946712c3eb2f;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h9b32c96e0dcdf0d50a3c000935f148c2c1d9b57ee4393ca187577a615ba3eaa2708854796ef34b0a1d83662e3bc984343c56;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he85715eaeed07d260318de4c37fbfa80464c0958f082057854639336447234efb9b74df75ae1713d6107a1a40a57bb453a95;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h737262ce13d561c37b24b8a3cdaeb08dc2d7270e451ef68d2a90ef6b0c56c03e5f9700b4aa50955a645c0c64e5c98c9c8ca;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8cde5f79c21be6dbc213868b06ad07e020d9e9384b26da70af0b44474f8f2ed823e02ef45639574e777b1e54b4cfd45e55b9;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h834c606cdbeca41974472ec451288d5e085ce6151b7fd53e2aa9259c7f17e3c8f1e8a4f6324bd5ec90f6fe76cb8b0efa142c;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h5076d2aacd63d10235a6ffe46f3bceced0c05958e99a39a5742bc7a47c08b356643b4eb06c9985e7a73b2374facfa5dd8f83;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hada0f3b6fb9af9d712ba88aae94aeb57b49e0936ebea9b9462555746800537bb00134dbd2283f3b4c33b21103a4af8556350;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h99d5611667f6cd8f0ebf7a36f35f02d94cad812f210922fd913286af47cd92c2dde9052db7328200b0f06b29eb6fdcb2dbad;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'ha60d08ccc02334cad96b7c7e61949060cd490c1f36b5879a1a0c1cb976e24151c0df6b06a0eebfde4eb9f436e7cd3c1f5054;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he05476d7dfd15c4667c307e37b2f6c93955b916cf249c2b493769e9347b00fc26b9336b3061e840365868a735b69b0ee708b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2b33814ffa03647f42f6ce9d36f7ba41bc014f0ee1f6d53a3fb4b270f7f5a85e9da86087b18d64b63b5dd11fbbb3a48d0f0b;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h786c76b6e03ce103a03713b0be1b732829973819da546559bb4e5e6c9fe26ede7e9ff603bf6ef7709b90f587d9b2d8fd1be8;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'he59b11cf80023458301ae9d567ae8d22c25f7e3f34ea82d38ddc0ae2e0b080fa8e2ad06c0c53b492010ed22891c7fe2d863d;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'haf8b9fe74c00babb3127fa0a33787486471c0c6e344e7ed0421dcbf29807e7cdc17b067fb1e80991ab26f03d3f4773851359;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h73f74cf06cbf16bf583bb62452001a0d390dc60f09857e33b0656f407c2ad0fc4e69894fa99706a0ecd8b2479abba938e925;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h11ebc59414f86f2a9e2d07db8b5afb2b8a7059ec9b07296b7b908151cc62373ba6b0642e925ae703e60ec3f32263789aea20;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h8e329d0aab7e14bfef46a74624d2d082dfcf63ec505fea7f05850ae07c319b9bfee18d62f114b6343fdbceeac803904abeb3;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h675223dd2f2297e75928afe2d3c5b14c2337720c1c768c2ae1f4693e70e22b9278472d5d098e5fdf6413c7ea9dfa238c9efc;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h3f5027b63662a32a04c157fed4b1a47d667d9edee0447fa247e4f42818e432bc9426c8c85d9f90e3058dc1d43e604e760b89;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h57c710100ff4fbd4dffae0dda6b788ae045373f872e45907079fa2f150ec11f1771a2fbbb0cbdfd5ddadee0abfce8a9f5284;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'had86416ad3f036debe429bc272cdf66145110c292cf491ae5532394ca77a000a380ea8bb93c46fd713b33891f72dc32d3435;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h45bacdea93c9a94cc9dec1b4d5130564e6ccc89efe8cd5c198694395ac7bfcc1d4bee8d7c91f8c364d6e9409a81c3e9902c6;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'hbbcd3342322ecec8a143d1612ecb27de99ea25bbcbe49f4550373e72d404b88180cd2a205af8cd55e6d30d90ad359a319468;
        #1
        {src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 400'h2131034c53c2a8bb994b48027dd21ebf677e70538f97795759e65aeb9f4c5fcaffd76753403945529d9ed5e8ad4ca7390222;
        #1
        $finish();
    end
endmodule
