module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [26:0] src28;
    reg [25:0] src29;
    reg [24:0] src30;
    reg [23:0] src31;
    reg [22:0] src32;
    reg [21:0] src33;
    reg [20:0] src34;
    reg [19:0] src35;
    reg [18:0] src36;
    reg [17:0] src37;
    reg [16:0] src38;
    reg [15:0] src39;
    reg [14:0] src40;
    reg [13:0] src41;
    reg [12:0] src42;
    reg [11:0] src43;
    reg [10:0] src44;
    reg [9:0] src45;
    reg [8:0] src46;
    reg [7:0] src47;
    reg [6:0] src48;
    reg [5:0] src49;
    reg [4:0] src50;
    reg [3:0] src51;
    reg [2:0] src52;
    reg [1:0] src53;
    reg [0:0] src54;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [55:0] srcsum;
    wire [55:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3])<<51) + ((src52[0] + src52[1] + src52[2])<<52) + ((src53[0] + src53[1])<<53) + ((src54[0])<<54);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddef6ae9a8cae43a4e83d06e8ea83aced7443b47375a43a10d9dde30db3ace2de7e9bfdff95a5bab68dcf9d1648471bf1140140938a3a3d34e86a717f46d38d42ec233c1827eba47573bf0ed594f34aee54e0e5161e10686e0e7fab0c176e8333766;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd6cdb35e8a4c4122db3ac3b8102374915927435e5c96c0840b30c22591b068821e1781bc1bb6ed265968303747e6b48d6307bc8702291d31ac9084ddcb255fbf573d4c75c9a8cbe3e6c7199e797d99e80cc9f77b86b264b423c921a9f180edb1897;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92b8f3b0c7065a358d2861c2eae73cc32d56159c31ecd2ce005e74ef04cd811f1e38cb43cdb1bea4fcf39adaa57aa1a7a8c14ed59388b83d59f3e082ba01be9adf6d4d5072c57f1abb70b615cbd56aa144933a294989d907b402c68a9f06802567c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac20f499596564cece2fb634eaa01b2b8b9e41630c2b10ae8b3b8d3ef48f68843be62ce7215bb137e433abc19edd312358e1cd887289310bc836f7d7aa02842e2b1ce97e63b6f7935ad2068b62019b63710a8559c7859a90b2c2862ae5a3566085f5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf3d8cc4179f250567bea093182cd7a570d670b5c1bf8622a3a9ab30f59d8820a92b53b71adfefdd3afc95f607a4c817314a4ab1f94a1add84802bbbce95cd4823c412a3673690d16776af0683bba54daca2b8ea4e95b3d00d339d015cd7b7ccbf2e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had48b2215a2aca633c1802d625974fd1a07b824c8db1a941ad90cd4c2975443e5e72ed7f48092f22633b02bbde65552a7a3e5f79d03c5fcd4f5dd271c221689ccadae469e0be0e8da24a2ef5da5c730a34fbf534bfe91cdd55f8ff52034c8ad04504;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5c2dacc4da4ea3df2d396c79f79bb2ab2e3651e4cb80ab9b9c639c4539ece874b4f76b24b20b9163a61c3a0c37159ceabc6f35d665bdd7f987ddff56eea0c84fce136ee2f8b6d7acd39c88bf62c9ade567b8ef8d018daeb45f810e4b3525ab1ab79;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dceb74ec9e42db6f26bfc5c54a76be1e8776686c039c85e5e85febf4605667d9142fbbb77f560ba3a700bc984e3ebb4103f15d180799c87c9b68c21f4532198b3a1312f390de198c5e4395cc2f267bf97a304a32cc749d6117b148952fd83dccf60;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a2f0fb9fba801adeb100bb8f46b2775a6be1559292b02d94064da6bd8c3af0dbdb5e3d8a195300c4f02e805fd2ead017504ae50c62eae8a3e671267c11026a7bfde4db4611665e7c8424f0ad916b38d133fae5b94b4270328b0a92cd0a1aef55f0d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he651ee1d3edc26ac4634a7670cfb7f517d019c8783c3663cd7a7d06b27ae0d19a9d476ff467be40d25efa3b4af7d7a673db9cb9d36c17d953e44351649885602a8919a0671e41085ba9476c2af9c4151f55a1e507ff97687a15e614b5efaf6f20c71;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d9209e83e6b2775a7db7ad15b3ad515f4ab99352a3b2b3f431a40fb9ab773d9fb2861f7b03f21a8476e00bc6dfc57eadd0a42ac0d8d958035f77d573ebc42d0bc237a8a5c78f946966fedd4fb5d04b57373b510a0dc1045f4b61189dd0e009b57a7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c4d8fbf76d5dde932284a6d627fcc5cbc335a49ca042207fcf489800e69f8bee600d5ad799017745da9079c4fa60733033551e33f0122b4e89decbaa547bccf975964dffa6e82a1d77c4f3c0e03bce871091315ad0901fb5423929046fb0c9cbe3b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdca89a959b0e12891fcdb3058cd2c9acaaf3b96307ede8b954c54fbac248053da1b3364d38213b73f51cd7cd00468b504f907bbac7be40aadb331071001b35d882796331b36c2e9a5a2cdbe23ec8975531315afef241c9fa32de87f8cd71af9b3d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h350fbf941ada0370877c5d80892b574b538e5e25e0ce2d4579efee1c0be3bb52e4171484bb44425b061b0154b608ecc5a3459506de11c2b7e303c21602990b5807b9443f1f0e151e82a7d2122418a788c1c972c7f87d5959a3dc01e10b3e511c77d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4b77f14e895ff6fc9b5888b18734666c28bd463b1f8804d113471784ba401ace4521e76ac96febe42ba175b89630dfed64f1226bbf6a50fc4fa59c7a13e240427ae6fba3bfab2e6ea77a340d8ecfd16863fe856f4614688233db9878914b52a9116;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a957a3b03f5512e721de7884ab875798dae2472d62dba8e4cc1806711f670cb677238fe254062ab8f4ae9502fa7874a2b740facdcf24b6dd84e2d52883a27cd08e8ba6de74219544e53809b1c760c9b6f16d21d73efa8c695ad999a68e15ff31502;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h440de51756ac273591d910b8018895c53abccd74f22b5c3051df78f7c4ab7865acf35fe35080529589d7b84e122d66009a467530aa1223144e7e71096a0bff900ec0340213f9e270c22087fc346fe4cad779576dc60673644bfc572e46c69fcd7cab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2c86f062eaf8febf3072e4e920c3892af0cab3e7da1ac75b0762c9d81e2c08308a3f8ef877d3d7929feeb7df82abd19fd1fa6bfa60da99003eb017386790d63f71a0936d6f463353b18e864a6bed3ffd6376c481c2ecd830eb1623b72b2994b276c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd014db666225812cbf774309de66c3191247ef0a2c2a4fd7fb12e33283fe4f5695dbdedeeddfd73e4d406bf1efb3afdc08538826a06c06910e881b44a72635f7713c178462a5783a0ba2b43869b3140ad8dd52f14de991827d76c7eac7cd1a15676;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74629f708e2523865e957d926f5152e537b9a95b309c277a2a8924fd35dc963e92b443b0148fa05b7a613411951a28eeacf225c8320b3b3233be21290c0f3d400ea69d9b7d79d7e33be8be041cd0cfaa8bf180a5ed196ec3663b6beee97f7eb319b2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f120a94277b61429956b8a613a63050626d11a3dcb9eb5f84784836a2e0e60cf7fef1ff037de0fbcbedd2da198de1b28e2b84c95cd81f287cd7331675009a9a6563a190d735b736b130023bba3b151dfa6d61e9c90609e82b6303f5f1940eec9995;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0e01a4aaddfed8caec00b018d6863be91375861437113f59885f7c810bcd41b61dbf3c5b2700a5fe6aebb4aafa565293e284d899b57e40b9b1ab22bb286ae1f3a51e51703844fa568f05f4c3913f54c91a6b31b04d2d773c9935a7e91f296f900a7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3438d9791d997a6da7f82d1cb9a1468f17c392e00c1f2e98f5f77b592ffda47bb0f0e74ac64d5c40c3d511a26fd0cf3975c6d92fb0632df8e90ae744faa676791f9397fa0d33be04e701e36caa8e094e093837a46b124c5b65941ac916f911333f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h661b443e25aadeb8c43c29da04feafd2fcd62b7e4a897c859294e58d0964a16b4be8c320742d63d187cb15f1dcc1edf384ca82797b7e4a4aa0e5ba563261c5801a61340e76b0660ce8610ce14a884c277587e5f792005d85e5b36d0ebdb7ca1e5f9d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h559fdc95211bab27b005d6e0cd122b72d1ce7fffffaa11ff557ad77a036700732b21a21db86ec090f78f9c12062dcc122beefa55e295cfd41941f9a0fdaabf6506be7453cdcac0e5bffd606c4140c093059a7ea0456b7945e73799aaac0a258afd65;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2bcabc2444f8564addbea6a01764c7708c137e212e17f009fcedb5030cc05ccaf6d21a081dfd8a0ed1139bf634e31a854c862ada6413c4a7efd08368e33e7f58ff337ad4d3749c901cbbb7227958162277329d58a9d92f41476e46a8ecce10003297;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc81b7e61c5873104ddf554276187205b7c7dc95437beec523996b76d76a7bdf7313d29fcb40c3782d27efb617fa414d55dde8248669b4ce2c1252a2aedab334c4128b7ecb82ff0f979fb92349b985e421e7f8901c4f4bcd6979342bd953c4e33e4d7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha06ecab2c98e85894c181f5f421fc9a6eb5fbb99ce3a54277e2e91381369817de1bb27d6598e03e0b9bb52648b9bd0a5263e43bd7c7232d1984876837848a55acaf623d4571b867d892e65c8087fda7da4a33c0563818aecf9844bf3c0da6887cad2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd837654bf4dbb296ed099a9e6ee97963aa2685c38523502c7aa20ae13fcc486187f70dd6445d22f91c4b218e274ebfc6e597d36d58c1ff4adc7511e5c94c0eaeea9f0ac17d55c1fe8de270ea544f06bfb96e4f5c7edc75e673da621b50b3435dcbf5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ba2bfba1303915b5f844090819c4b39552a852216e1d09ff3d2ea8e97d133513fbdd23fcb2874415a69104908fdfc0bd17cf00dcb55d6bb171f457f4608c1245e7bc6c48fba1fa085362f52df57fea8f0d8b7a2483e90976eb98831ede882f9bd90;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9462de1b99571ce616e741c634bb6210f1d8e03e6b2729cd054d9f581984d7ca15928f7a921794435a71259a868bd47d17e1e991d1bcc36d53087e43dcc63196f60f71d43c1d7bc03ef552c8541083ba3932dde7dc5788f6705d097b1711830f01dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc83391d048ac4072d7754d101803f66bd805b69b96a5c1b4c34bdead78eaffde015ea810fb62baff0dc7d9b54c46be9401d2cd5e87e6d9c7e8b4e8883f5e77835b73e1915e3c09e9d9139dd8272032f4927d0bb1db300d024dd3f69fba8eabc1466c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h295084e180d0a12883ee8d399df74d8566661d0265c729cc5d74c98316ad63fecf020be9646d1916fbb4b29f374a05507b9e6b775361e65ec1c8051d0ab94490dedf3c0c7af64abb4fe3e0a051ec85b2d833f8a9a5717f814699bbb5873d799f018;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb221d24defe210725f7e4c9a4fadcaec4d95438a874fd1c455f44bc62b5393fd3d63e485349e6110ca442a4415772e9d3f9d8c4103adea498e79ff2bdcf50b6f09187a31f8b6be02a3d3aec2568ccf93f4474e2e5e45725a4edaa521e6dd92f192a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7dd1a20ae643b973a317af4611aca96ca382d13ea48782c4ad0380c9642524ee97094e73e1a83e3ba0917cd2fa7dc9ee895186aae37c54a6178088596660a7b63889af777367bf2484a3d162aa20ffcbdf7c55d77eec426f1b5eb823fbdab77edb20;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he913148dd00c914bef772e9434b09ac1d77f3055617459b421cdf4ffaa34932907d8845dab49e57f3535611200aa8e5b95dc618753f0294cf20c1ea90d141f6812748f48917a4c7da116afa0c6f16ce8d2ae8cb05469abdacf1566e8a533a8d039b8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32b4d09cb7c053c10016e99edb69971afeb286779581f57bc30bb4a2b180ee27927f5100da9b385c7697adac1fb2ff5b2465536f789979295b8a3f453c850e5b7b5d1367fc90604e716d7809fec4727dc8886f760bc1c86c71585687005c79cf871b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ffe6b5eb6d4c277fdfc54528f00e6a0d0c5f5b6ce3b4d049b12a37dde7c5f1d61447a9632ce4aff4aceaf6a94d7002e936859e10699d3cd751941a01e81c57702e743a70f6417e557296202e25385da6fa1cf27bb3259c43b36aa1c57c94549546f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd250e281eeba4d320543d87f8645307f6e7ae14f4ce01ebe06e41efa3d4d1c1dadb383a7ae21941331ba692cdc449595f9f380993d5e96aba2862f9ab1bc722ced83cf41f98a79228bfc324abfc51b320dc45f16e41e3d0b512c99b1fdd5978b21dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57353c29dd0b37c15319b024875f24faff56f42ef14200b90a4568dde4f191ebe658c8282b54ac6f797ab2b703aa1438b48744e318ff48a26314d45c08d097e87a5e5c294c044f4bb8f0cfcf07d1865166a2c84a2a2c03a51caf64dc903afa7d98dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87b781fc9b55dfba412b42cc185e1ee594fa75c9afbc6bdcbc2653750709c901b377f50a2c1261be0b2c363411b0e935b70c1ceceda9155af14e1fb9c1b5f31c73cc45bce95ba75f41bb2e062d3dc0dcfe32372dc33783a579153c6eb2ba69dd91ce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13d84073f1d17f3e1df06388a150c6e3aabe81f1a59118154495f4ccf4e35999252bff76ec79c9f2e65f154fcc36f5915c2e1a6e1a335a2b13849cdf5c9fda39d91ab0ed469ee6dd982b9f087a258d635af61d06f358964c494fbaccafe74674f49c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6da85bba9ec5f19fb93b724ea82900c86bcedc57d6a83308b16258667b13b94b6dde5d4e6fb942327760cbb494aceadb67ca05c95e62a2b20d541276fa450f32e4b87aada7e1ec1b9d7275410f3e8d3a2396b6620e37f9f46216ee1d4c4caac7c305;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4436f602c95bfc6f838e970f86b1fe3da2c72f9c6a309d6ba3797b24dcdcba0cc0b9b532361667b83765a7db53ab565e806d6cef13fa33ca574efa9433d44c969dca400c4c41845e1caab453fb8b67b687e50d403bf7ec102e60629098903e435b3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb74ab5f5c2c7e9bfcd7c8970f1b6322fc6dfd43220b7eae5a883a6d36f3c6c7647bf15461c1a5244e0540bf536fb8c71143480b65d68c22dda0d69abc1d602e0e86c5d78c04ac73fe95d89b9a7e5f7acd840eea14945b5f62ad12e9a64aa4f5d25af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3764e733e5de3a85504c01367903aa2e5f1c41c57e5bb592b23beffebb1f6a5c678da3de5682e514c1071e3a3acdc947af6957a84769bb8b1d1aacb545e418a75bf65257d3db232de9bce6853451bfaf2e4d3ec1225b14bb2e8643470f7c47b8609;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50d962e19c1ebc912d462e0a0c818d57c73414ef4a179f0eac9f0bd8a583834587417e13f5ca815f9733417f8bcd93fa863e22717578bf7f12b51098a79addc0e7d5ccdf8cc34b0df47e971425ae1b4a8532bff38a2144a8d983b44571f08214ee2d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77bbc3bb37a20ac2c06fe3c89dfed2ebfc2bc04ea6d5376e38400f0279bc2976c97a3c3a08573a8d6f58b8736f5a800a6cfa11b8598c143074e54b3fe3d260e0a9b04bae4993e26fed62d606e9b3290b24c097e321ad6fd65950411046684e581f34;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c76c482bba23ec578a003a659a43550995648442211af13bb719f3ecc01d7fdc31bb337ed157e5e645e0f5a7109aef8d5593f20cf1a56e03d6e6a57c41ded540e1517e61f940172deeb938663707aceafc5837dcd2b9481a7f7e8e72d6f34cac507;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h930e7713f2f75d65f460637cadae0839eda2b25ed83940b2c836a2d80c4fadde73e33d120949280549bb6775fe491056ce9a4cdd78632c2989ccf292fd379a9b9437f7dd98d1a3bd78a83664c264254d326a8849713b6e2918c72f469296f2394316;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21ee2b77a9a2fa009b6c8dfd2d8354d77578c1a4a66dc114c7376d531df298bf481060d9d5d8fde5b983eb9ef3c52c5460167df0fc0f8e0f711028681a9a444d295319617c60cec1d4232b99915c079a15dae4448ef0e10647007a101b2891bad8ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd98098855bb41f1612aaae7ff51e08add41f5c2dea630b4871fa261fbba903d849c1bea80bbdae4d9f9c3ed52c82f96c670b1ca7d701e83c2023bf9b058b8acebab8476c408a8d8ff89dc2b7bfae326b44591001cc1a9bd103cbcd3c57f5fa997648;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79c97a296bfd4bfae7811a702119d064143ed99bb0755946c0e0e4a47c33da98e847567fbf7fdcc401e30d949cdb65fdddd23b554be026f3117e28ec0109c28b357996666cc20041cb760102e12a29a17f8f53dfc2f6b74b90c8673bde965828f152;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec2764bd2b3d1decf5fd8e06ae544587d9ca7f91dcde4e9b3bb45421c62aaa4bce40b88005d097de696466d8e04244216fa416328d5276de8aa645d6c2db113c13dccefd867ce11de211a59ecb70319929b1fc7d53a2c0ae145c75cf17bd48163234;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cf0104ed4c2fc7a42731e41c2df3e32cf0e01e607565e1f466feb2de84c64b2f384990c1b9e6f44e158f114939610ab247fab45ab880068a0dc18c97c8e718cf71443bf782e6ba56b182a256d60a3c142fb2bfe77b95fcb03d23b5b78d86961d41c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1e9e2620ca75bc732c6937946444fb7809e980a2838a1c37af7fe8b851785c82d409c78005542d44b287958976e3f338a296e10496f73b47536f52625a15ffdf5b4b60844e6acca02e42a3ed57a673a4d4b662d8f55304d4529eaaaee4eee7f60e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb3dbaaa6743bcf111ed6dac2979af2ba849473d78226e8930af572df99100fc449ff47f0689bc6badcc00417e6ad098d66b7f2d59ae626ade6a960599acac7f881fdbfb40826ffeb2e215acdad4078b73e2bdb1578174ef2c7daa537062b4cd68cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h713dbf48633407ec2dab593afabb02a238f454791cdf167195ded7bb82090ecd79c059c7959ffbe048adecce64d5e5cb018d92446278f654af21ab8820ffd80e22318b3ebf4723392d9760d4c9d6f3aaf3944e89260effb50245e2d225461aaaa014;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d2116c6362f58fcbaf522ba8580bf3f4ddd69d1d823957ce4eee17555b08e577fd2e01942b69c678a2d1ddc2685727235e625f29418549b04687825e428ce483d07b5cc4fba9d7196a80a6b95e4e5ffd5c1865ba95d5f980dc2f0f13b82b60118b2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5c32fac76ad8294eb95b793f4cf0f06aea96f139f1b72faaffee25c5df2b72f92ae973ce07b34b7e66b653ccb2c0d2baa18dbb56792232049b516add5fc67367e00733caf47586b62c62a1684d436abe1b69f73c101f5e0952e90f6f25a30e729ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37c0f25a25e5e0e8a469060ae983f6bc21a827212b9f1cd4815aeb7d525862ca3cc333ee7d61371c2224a83351d253b57567e8a047a8c9ea04e3a7d4e776b0ad084993cbca9c6cead8713a90eb98626487e84fabe1417791d6a6f693773de167fbfc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h618aba6f5e7d646ee1a872f4090db759d125ddd421a8632083c5b4b7f081748f2d91d0224eeb28037c03f1b8a47966fff9e805ac7910884d819240d7492d7da5500d6413b21dbeb9533e11391fa637e9aefb2104313c72099029d28cc552353ceaed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h967631885a802b7f6985b548a745dfcb5b2556d19e9dd35efd7d508141dec72fe15e8de11f4515467511febd9f623d3be5e9e6c46600a8fe74ad1364e8d85d18b65d3e586d72e31fd724b82ea5bd497aed7dff48fd8cd567e6ab0dc831329716182f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h496e5873651170bbbb205371468149d364ec847fe4824a4d7c3f51e3deb23f40eea041ddfa685dbea9681ebff5bfc5d66576828a1374206bee7a510dc03f54633d1753e4e28c77695d70cb95fa57a7ff00d579bd83e2137e24cc6db46042f4542b24;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbdece7f566523c451921f210145ed89035975a56b26e8f3edb6c12b3143954571d8589f2e481099981e17e9f7115196ffb6b1f9d63d39922535ee84fa3182c89f1874f57adc76f5f7248849482b5869108fc5edb3a1ef94b02881138cbf2619cd53c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc79554a83e20748e53d154e7255c18cc8723b0fbc37291a939c8e1407b4ab2bcb11d2c3d16dccb74f12e7d9a5adf22fc11cfd649d94e68d500086f6c3a6f8efe895c58a0ba0dbecd66efd5c142ff9cca504305e263d495c605e732561605a6d89a86;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h365c510a40a9ea11b3d47c35a3fba3605ea98051e027359fbdc27dbdfd86edc936f8e6e89c24a899ca185ba02a3cfcab09361de6e3e4780824abc4206259c72c6b4c5f0fa801a0e416ff6bc860575c6a70ca8ad7f706e43a2fe696d3515e7aaf0958;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h278c749ac06e4d7169871c1bc0eaa76a4284845a4715b78d8aa73e7a24d8609cd7b40cf568fdf56f212fe1d597fb76702d46b0427e38445fd0e33832fd8997d545f246483ec8b7e785ecee653db937a904d310939f5aa979bdd64e93080f861a608f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e30589e67008cc773f8cab06dcc2512f1eb0ddd15e89fd63aa2d23c23be0b3f637208ecfa95b4b5b12907370b7d528211d5d77b5d3fcfc1463f52d7f1386fa0cb8c01267c5f1014da8b5e761111bd115c785f3de945b654a9fcb987c4be77263a0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24f2419738f2bb0e79f99032430c7ebaa56c91b729cdfa5cb8dd155de8ba6423c6672f5bf5e3a423e2aa81093cb1a1026ae89c4f919c7b950580e849361fcb9707caf99d8d22c064935a9578a140f538b83d3940b9caac86b5f58f97885618e02827;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd80aa8888c4e8e48e619c80ec24d560c8d4d4c831eb200c5710357ac271ad729669f1c48b6c8da008573e516e98252cf8e08b139160a180687c3088f95b7a81d68cabb66717ef9e08fefee5932d03690cfbe56777cfb5a9b174817c8bcb27a2c2fd9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57077574a368066d5f98ab25b8047dce9bb9f501868e5f7cfcb3d45e8028caafd9612e525c639ab97360858c60c55400edd50ddff6c492673730037e2b457a8f586a393ffd80fba6c7078dd7cf556dd766c0d8957c249ce41d84b3f0af7a4cfea579;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5580a2b791976769206e716b717351fe88dfd6c463045a5787a9f68c2ff8e3c2ba4af8fa6b184ba7a690857f8c0d81aeec21d8850bd781346affa4ac16f966fdfceb05e6e721308baa1083b3401854993579f0f27bcb7dd473bafd952aeafc9d2a67;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc87b839175924f48b95a3a3ecdbca218206222dd77b1db91d6b4a3af3289e5745fdeca18288bd5812bc293592ab3d1246fc548cc29d9ecf85e35dd3a46d422216ad8e9d55bd4eab7b9255d8d62aa70e49ad4aee60f8c7381bb58f067c682f217a8a7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h692e79045e196d18eebdf984f57971a8aa442411516b1e317b48489e948f42d1020a7cb301e94508bee03a37de154831f400c51efc6c624e0466b8c1feed786a63d92a770d8a08576662764da27b834cc47fe15fbbbfe928d64d5ea3cbfa26f1c368;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf45887b3ddd4e982cc5378050392cc5b20c7b208b1a968b83713922c24b2d6bff4c5878dab206028c546e2c454f20e29b92b2df9cf45a86e2f0ede477ac0be2841df695a8894e174f6b27d0987c52b4df1f74317e0b532fb7685145032e6c4cc2db;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee5531fb3efacd1121f74f66b524914e27ecbdc6cbacf0e0b2f8f8692786652d7b4d52a4def845a04b98eaa0a327750ecb612cac1681f4af22b633f27c511398e1c01d0138c0620e30527ade3f075fdbb09b299a92c5adfe55fc48ec71cf2e223989;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5027aa0bc2d16fc57442b16302737437a58f016204282f904961f2aa8d04d5c6eee951ab406a749852740256699878d2298bd90e51043adf007c456cead662dd413457a5ac8c3255e22b6cf83bce292f055d8691d5a81da703df3eb7a7a892e009e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7063ee0b6bb240aec47f7ea4e45340b511b3ab67596ec52dffa5909715fa317917eca727014346a2c02c5472674faec224ddc1ea98e10abe2572417b67a4dccbd659afbf4115de2bacb1654aece64e3eac0bae8caf88b27295d2dade5b61078f701a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5ad7b454b2e4e02cacf62f514a4b449349f3ae98823d3e2f6073fe9e266fb7867e8f55c91a4ec3675bb4c5bda1ca3c119b14f3713976d03077d276cf10fb828a5f8eb07d48a3d460e4455d0bb017bc1d897ed27c06da0947f911bd675945238a775;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9916e3d6798efa803b8c5b2d41c991f8286b7ff9dcda7db00d495a57ce5626f38ec813bf2c9f8e852dd7d3172245009cf38bcf8e6a98cd6b460e017446e478742808a86dfc42431adc084f166696c5a04ce091b17ad0ecc38825f028a1a63a378b3e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a1f77a579f9e2cd9fdcfa0a07034fce2a51e46961620724679cb698e765d303c414ae805ccb05cc07bdec92bfd291f206983c290153f06a1cecc8bf01be91675a4a6c0f9534d4093aa0c7ccd3cb9858571ad6b18d59cfb327988f618e30148b8b99;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd67d42a8570f404747cbac9ecf2a88e656d736416e33479014b882ab7c12cbdf29989e5ef42afe24ff7d76d6d1e9718c82519be3f25c56e2912136250c189322bf7ecdcb3baf2419819083a4269e478b155ca4c540374d5000504790d116b5e5af9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd13ed4971151dd1e583fbd1c3c422119270bb4a6e45e1afb10963900505827d3a69a684b4632e0535b954b42ad120ab3d74cf297172442e53aaf204fdc1ed32158e228d74a1524065052013085e281bdbc2199f274514388e28f0d2287bf46754e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94a17513068ff38e348325ac2029a7c337233fdd1666722661a503454216c2b7b0f1d17da63c83cdcf15ba8772f66c1f41e295f04c9f37e9e57370df717ffc9d2d70d858c759ce9047440e1609f23251bf7509652cc6b5331634ad423b3547d9b337;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9f1c63f45e54bb8695cdbdb53d7ba04fd9c8f82aa0b986e0cc3ba1d66586da84c64b2fe7fb894503303cc649973d2dc5e84331c59c694eb0d6b430f559d47484c5d21bdd37b4e6cf562fafe93e31827620e592576972358612a95b1e69b85fc8bcf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8592907bd5bb8a71a6db8eff04be6719a394dacf90d2226dd06eac428ebaa7cc7f001163d78e96e2b697af2cc51adbd4282ae703487a0b6abd4b08e113a373acf03de406805db96c967a70ea92534f62c9647c79042a8b7a778dd69ef280854aee44;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1aac6b2f4e751da8f2b51706a6499cace29ca195f64c7a65168837d2b3496f94179892a2888e145574405571fe67557493f58a114ecd1a79c430db23c202e00de142443d9242939926989342c1b82a4ab7f35c7c967dbe36ffbdce4596de39d186c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3ded08cea03c3d16b489c22309c97c274fb05484638481e6402aedbeebc5a4597f026ace74b302cec2578234c687efba6744558b9557ab791f2b0fe441f46943062ef415158c3a00479a4766ba62ffe8f1d4622c02ade249a1a2081b7d074da6c72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcea24e3194175eefa94a9b0500f6b4f7b54b902c373d970d2f8cfb06b482de21f9f31d2b40737ca4c97210c851a74c4d94ea05d47f4a47c78357974bc174ffc8c610e8b7370fec11141640b22147bfc7733f3af5866f3d8ebc3e5380036d932abf49;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfbbb9afde4a3fe407aef35173401e4c7a755f866b0f68f6b37c6fc50376ebf6fc1e5c3b4f3a69b42f1ce441716d635bba278d65b8108df81e0a4d1457dcd92f0d32761a8ff3e5ee8bd491ae2798b6d5117c19acd70c101cfe7f00ad7f80ed7c1b9d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeec69beb6313fa2c2513a9b8173673c9c01dcd13d557cd95d0b09aae95c3f4d2078f399c42e6c5e69cd4b4dd2b21fad7607c435f2452dd337d5de202ef6d72d503c868644eadd49b5855970761ff4e66a985f18985cb7e457776e2add4e8c665a98;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ac6694723d6e9b1d1e5b498c5dde1e05a232fb19a784c5f50d2f32371ac47125d2308195848a7b2cacbafb4fbbdaee93162640de3e8c0d2366b91bebe88c09980b8ffb741b0b9e2b9fd504e197e638d6a45453eaa751e0e1b1930ca0f638452fdad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20eeb3b17daa5c9bebeb7269c052361e3bc5ae2bbaf086abb0c5f4effec2abeba41cb10a4ba512e8d77e47baadd4387b9d70473d37334a5ed6420222ad41eb011a2f55bfb4bfd72b395c38e96f66d0e4675a68f3986a710be451bdf259895b329c67;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h395160d1ca1acd5f28ede81b631909fdf4f0f8ef4d12c643a4f0b2b9dad1a71c432f82943711aeb3f27dff3f399c940b271090e45f70b78ac0467b88cae6b40b6f53545ff6ba251cbffa1249823f4fc37dbf3f913735e12f62679bece9aedb6d6a02;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17faee8026e6d357e13c70360f44c913b0bced84d6835cfba2887689274bc40c1c4115b1a95b6c2930f09defb1ce4b8cdc5c1c7183e08482260ec6be42a0a2ae90202e22a8a6c83774b65677e2274ada8e409f13b6e3ff2186f39b4c8c5c18c0091f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he917e723ff3cb89544f523f5cf2452e1814d945c00eb40e83d78fe466c1d9a581885f76fe1a3689d20f4b04ccfe1035df2a9b13a1a6b83d2ee0f097884ed4dcf63e90ef52dea1778093017a91c4b67fe9c121e4064408932f0e004809adf5784cc67;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7e28904662bc5972169b7a04b252712e661fbf5a16d9aa800e06b1c09c5c52ee5fa4cece7ed3e4259f7cf5c911acfa71176062fbf104642b3551bd83aafa3fc39e7c770f98633d729bc2183a065bd4fc104bdb95e67976c817152841cb7a143a34e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6eb4ac721c03d3dd3863fc04fe716b139a33b682605c8b35006097ff9c37ada23db2b5355c520619bb64c7b805d773e588ca9f0142f451332f31971667e073b0183ec2a48a1459e839162e8c737f9cdb6312e7bc0e6e054a277a287a7f89595f7c71;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b7db6f6e6bcdbf43faa70da4ff22cec73c8348db461b9f40c2e7345355c7828cda728b5344d484d4aa8d19e76ba57f74e225d6c1095fb0a1c387b8889ea299a83d055d86fa2e91bf54906b7ac48caca23e496d66fb42afd09fd992f90fd3b587d88;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a9b980d14c724dca914ea8c0b87fa982a593bad560adea05ba08eedbbac8b63b243211debfe65f59733718a9a4881730703f17131e968602dd718248f4e6d3dfb098f6bacfd83021588486e2d98dd96c1b06c424cfe2cd5c429264e019e6865fef8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha87d30f92650c0b1b42e5c62a7c4ae385327518563e8898e9095c9ef3017b4ca85c360374bd9e0b32ede1ae4264702689988215fef6114668ccc86101063968969192735f57871611ae968775e36608197b8366c42692d391646f3d3fa436ecd2919;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4bc2e0e0daf2444264d068c8874c1b99fcad2932a841ef14c339e534cfb82360ef74e644faafeeb810915e40732b5a32b586911665b07b3b767eb9dbc4237395e78bd7ca61e60d418ea1fb0a9a5093badf6b68ac7df7edd27fdbdff972b5311a7e75;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c5aa46db512d71eb65e2c393e8e0ed8bd738f395b420614cbbaa9de59521a9878d268bd7da35349ebedf1bc072e0acb763a098048ebdca9eac36a6f1da98a3fc316b61e152d4d706a53cb5d5338d558a008b4b068a8ea427d8d0fd6bdb7524ba544;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ff17f78b34c9b318c6adc7451aecae92e9ff0b524021be1d9e832156c6e2c713945f528f7722d1e0262be5bfb3e7737a7ea4a7ca9123eb75bcbcc44807cb5f2aa566a8761499bae410bd86d36b3e9063d20517a2cafa471f3731123ba74894210b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79691b45764aad16a4379f057da475a70bf6744842f32f50b27cfec844ada3f4ce52bacf9d1b04de4166122198793604118981c1e4ad944bd08ce892307686604180e40d889846e14e55f9de143bb4ef6f1b8853477f6808268cfdd3872772079fdc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h654a4dac9cac7e1729c81f4d46d7f67d442beed92a71efd3f628f396720601c467c39cb624810d71f13ecbd387331a1a0ed454755c610eb376eb67b7390f7f7ca850defddac39895a70d9b964bc9a76fbc2d60b58a69028b15d011ef7d52474b0e26;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e850dd2784446cb56d92b9f170fd955a0ab77c8acf3fbf1d8b3f1423a51ed9ea5058a0837732940c9d1e7fc00854f375d18bac27c6f03e7f216f3680b1cc49cb4e59c5cac68a8f83d4e2db77bb0b5647e279ac02d5db9645746854ec746b50e3d64;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf475083a31f08476b6a9ce7c61c84f45091eb215a63c7ff1e8c0ddd38a7ceb36604e2f69cf2e9bf8ca794513ac58af9efda51bdafc7a31f932543b619fde7471fe721e2ae5e078819fbf866dfdbb1efc80164c64b86a95fd623b912011e01c4db326;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85b6dc0e34d838e92aa537a4a104f1ad7c43e71f66eae55b67b2d859bd83674f7f8ab81c43e6bbe38edd95215ad46b34521f73681feb9958810d2c27379d13cdf551dea1d84d19f6a194499836b01b1a6d0d7beae94d5702db63ae7f0ce90d95a95b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2be154f86102997aef5716dcd03c04fcdf6ad6dce205a076e6876e4fa64ac276c79745d0ddf808df8d57c26e0f9dd42129eb997f3f5ede6ee855a720672de3612d229cdf807506edca5734a370544cef80282c2c2405e0221de74a17af9eaa9e3668;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h998e684f0ec8b6360176df3aa5ef674a98bff7ead34b7151d5f5bee25f40e50fa44bfe796f20b5d9e2748e86d0926be960832d3ea1c892cd7525ea274123f0b2b73926a4e2bec357573e45176560f2a1acd00cda382c4f66e21557773e19236c5003;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5dc0722565da25952d18f5d649a317a28463ee132f720678e6360e4c1dc02333a588af6aa22548247dbaf35a7d4d45204e422558647bcdeabf74de0ecaa39891798c7d610f0c5f9d654bb90a0cc302d4cb235e8ac5e2ea13284515a2e7bce9687477;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1a9c8368c96c90ab926525164891f814dc1b15ffe51ea24e2bcfc6bf2ab3ae6617c5f28e55d9b103f6e676a864b395c871667b4c1e7b7b8091f66ed29ffce5305874c099d2f88c7d4bbf29cc85cd1813798bbeb210a5a46b66c273934d0c8deb8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h486b790d96d2b8df383518ce647d4f2675138291595d568a0e1399351b55c37762a0c92ef9a4c8c676617cee2ef43258359a7ae46e9f11d8930c2a0473e2aa62bbd5ca40fa1bab30cd3ee34b1e9e7507b0ee8248039cce88f651df906ac39fe85ef4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h802dc6aca190bee7e2e240f0d419ebee1d42f974b4bddb1353b9f0f44f3483d4c11f959aa5d3ed4361fc7afb732a94a8a4cbb3a66ffb15b8856ad13dc138e7480c537a04ebc139fafcddfdae1b219701890eb0d2b8586244c0f8df00e75719268ac7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b3a26242a7da28b6150d442a68a7e47aee1a4ad084145269bfe970214073c04234e2118c7f7950346fd57a402f2bd5ca866d30a04fd03d66d8f7b3b3e436e91e321a176691b134e7508c4037100e96781311fa2732dcc3a05fcde30af6025addfd9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42538b089684c71ba995262c91cae6401cb965e86a4704824d392d90791fa3a1f6e975bb118ad8cb21008271441219d8e8c8d309e41d6ecb4c1378ac652d7f297ccc8e6b4028f579891c3d98fb75ec187396675971d76f36f62c9308d05360461707;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39d61d759c710ca6fb8577eac957475a35eb6a52dc44171f47ce7a1b7ba6cda609d8bf08405c53db090847591d7cf6f24234ec1251cc51468dda883bdd1b09b1021ce0ac4508037d0896593c54d570512e780dd46973f590a981bf6574cd6f255dcb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27663f7361a1751d5eaa83fcb45c0ad30e722b1669d5658645175533c70cb7bdd37ddb815ed86d8ce6c8fa7212efab4a33ce5ea882b245b0455752448b8f00408fa6b2b5b4e345cd55f3ca963873dd46210d3acc8db5060179338acf0599ac6d3cbc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbaed57168052e80e9c9eae97e9aee524538a05e36fe88b68607c4328007bf6994943d632cf86942e337d5ab8190bfc641f3b4c1d26c6f11624e2a192c2d973cf3f24ecde936ecbc6071f7db41ed9a03340e292043600f5afeca08946c948bd542b4a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb708fa0acd9d33e6f65466141b5ad91a75caeda633eb01d8ee455be4c70ab6193a22728cd4274d9f6db0d50e8f9e78779abcc4c5be0be2477c16d38ffe2c1327c4d985f8ad78535a5a1f053dfb095afdcb034a226a38bc4a18f39a9e33ed99cc28ed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54708f31e407923cc2a7ea8610f448c784dde82d6b258117e8e0dc6214e1693339f41e91b279cc292c6576b6d73cc1261a7eef21a90b46f3886384cd992c266ed11e74e44341833428c8b1388254c51aab2b02595765d25cf1bc8137316b39f7dd28;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc51da232068d0747cb517a831b8c7d62a1b095252d001ea833b8cf6dd4101cfebf8414f07d56af0f51e3f5c05d797d1a6e3ac69ab88285ff0f6bfe0ce6a00dd185d19aacc5b1a7cbf15033748e04bcbc9647558d5fab80f13a232e9da34bf217745b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacfc470c4aafdc1382881e9cc0019363c2a88bccb71cde10c790631ef8a05647f119cae21985e593d679c9e8ffc583e9d2665646fdc9e74c85bd47119b5fe51424c385a373170f6a0bf8aececffa9f6ba0e6a8ba07f48bfa9053a905a33244518030;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74a19d96704e2c3900cce2271805ee58f3d482dfc9ee3b3c26ab32aff3f12a98a4d416f1a256a4cfffbcdf3701b37c55c12eed15302641d99dc4c59cc3daf129a5ebe4fc7a813da040283652be56c12fe5316d21d2d9bc615c6b556fe6c989ae649d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he089578e025f53897709bf403b297336544eb9ef73a4f9e14ad664c62a4f2477816d5be4c50290a4805169f09351607a1570815d55818880efecedf3f5c3eb6a41d2f7ca69b0b03958ca7706d0750421d633540cedb92d2d7a41673a1f206a0acd03;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f6460c5928b9731c27e1d5d130dd1c19ab23401479c906861ae8d79df1a7499a21e158a49aa9a3c0b89afa3a162b4f9bedf3786f7b48f8bdb30c974a9b06c942477a55e9ae46e632f13f5cb73aa982c1a5880353691793a116f136276f51cca37b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a195843bf2eb84d566cac3dc08280703188b94e2f0fa9dded2c92004cdedefa1f3bd2c1b9ef4f7a1c62e0a4b88a08f22a88db1ca25135fdfeb06fb6cc8bdc42108b68dc6fd4c1563f756736aeba0410041673b057b5f180e83e0441eb7d53f7f543;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c3f3bb16b31eb4ef7c2f84f799da68cb10302d634f7a93062145f66afc9bd960455776ad88a9002d12893d4f2d3672ddea20a7a19d6353af0c541e67186e8b03bb28bae4674488c1c35b8a2224a8a070210a4bef06d3f47dfc109e5a75b55cfabcb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h273980eda336179d1a4605a47c7b963f23d266885e6a81c4ef8c4327385ee922777c74c7e4c40c4739bb3e7ed0357c48a87f15fd3f21393e9191015f3b6a5053487b7c00ae916781836c672d5dc610ddc408403ddfedde5d2687a85412e7a0abdd5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c538f3f5f9e64389e514ce403d4ed7c11695acd2ff6f51c6d5a1fe59007d29cc854d3e123207e901b2a42524d44c956c2be698c3bd5183dacb6cbe5633206c690d3135e7859eb75b50af030c172f2e9aa48cc4244d128f48fdcf4e1eb82fb5f3ace;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf95c7dee503e1ea09261c1128befe490df17ea1ce118a7bf8b204f6be166a8c6992bc381ecdbd2534887586b00e0a6e89e02c476a124ecccecc0583f59a78bb4b12ac91b2121a83a5451d14ab5a682bf9ab5fb028147b33e3f363207ef499e410012;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39fd13e65577365d7fb5d7868798bcfb937125dc41437200c67350867869b7f51a1a91a63c3f3f400ff12559126e7dba1ad6ece4581ef4062241c1049c034ae884b544b08addc3bc58ff86d459d0b009dd1e2a2466207bc18b38d07502d72d8b8b8d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd524bdb1052bba37baab7caf9c1e78ddff1d026c4ab59463f846f0fd21f7bc4f5eab7fc5f551ec24888d7e5a889e3b20e4525c34b5146df169d0882820d2fcb0b7666a7be72d0a59eb95d79bd8f13f7b07ca18731ccbe0a713e7a56feabf37a90f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d70b663669d5909de7192ae787420c066c2bd7d1c40e468105010b12de4656c57bdc0ebbe2f467cdddaf9d9975c8d436fd0f1ebdc2764d10c4d1db3184e61127595bdfb30f5abe0e289250b52afa4115b6c8d3db9da2ef47337c9db8a075382ff78;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ef81dfab44e8e04cb940c1679658cb8ef6e5ffb3a58db5cbfbc92b93eeba16e294206928be4554370aca30f156d60a25d150a9c6610914d6bdaa1865b2a4cf72ad59e13b2b4864ef4ca5881e811a149373aa7c8885e18c67a649390f3665cc1f320;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b2c5bae8f177381a7ae14ba63903428d1be3c3aa2dd879abe5c2da22c67bdc8b83183dbc3e20b0faa9a0debea2e7ef6275961d41ee728101c143e7f5535e988efe2b7a2f327e2f6dde521945d97e75fc58243a7d9b6af1931ddf3e7cc946f928f13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h762833a9acdf506437408590c74a7fb81ea8c28bfbc3272b9c3f248971a5b448e7bb6c9f10a3297d4841033d351debf8c95bc55e1d34b6d810137b528d37e95fe83f8839e123c950f57e84af302e9c77e16b586bfb5cd3e87207d8aa228d7c4fd38c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h971d76a36424f74b74a3ee13e2fdee1e1c6c8ceb2052ffc4456d8b89d780304baa9606ffc323f95afc46580ab82ac4c10a807b1c3a8c2e9d0902b22ebf364d8b07304d5646584f4093d2109653854ad748c7acac4f24a72e6aeefd308ed8e85f3b16;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f18db529503ef76aed6621b024ce5ea1379b09447b858692031064475df854d9248118320940c552074b9c826e161b8f805927d72602c9f70ed1bbe3a91d79f70281de54ce11ad37bbae885451410c7ddb3391060b0e9b7f501b4b3e5aa0991c2c8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h919f5cef52691597673d5bb6af4c5459c35c563856a3bda7d1ebc251808db6ed570da8e5fd1bd5aa34a3a6f71adac25055707eae470ff711d555b95c2c2cc56fb5eb71bbbe058cf6d330b3e790896a344eb63c612746da95174ef607649109d8f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e4ba1c691cc915e0ec77d919d420dcaf25ff761f56a8459d111bc6e0d8521bcee818473e7a3eff4df227fd5ff747f680a2f19f054035aa97f5751028f3e234e4510dad0b4596c7ab7afbfaa065d94bf86936554ddc99b7e57ce542f0f7ccbd86f2d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7d48ecb94df34d608c5f04276fdf4e8906dab3de6ac28b67558cf623f2c032a53a9028369de4ca70a42beef528795c7bbd9e9f0da50735874af7fef4df68721e4f03deb19f6791bcfef859630f471349fb8b9a987082c7689aa4eb1215280ba869;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h642134f2f089fb9585068cc631d2c02e824e37be166b0bd27ac0a21c1654b924a87c606852d65483e52a34491e5a39178ecbf6a03200a0176f5e740e8d6086345773851a64bee37fd54cd6bb9ea48567ef4d3f919f8fef4f9be6e56e3022d204ed86;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72f04a817caa36edb53a4b84aa155ecf08467cae8dd5a0877a55d5a9c200b9a0f766526180c0c485430cf3d3e23072a002a528d2aee58ade521cf1369c7c891299b5584559a63c8f66cd1a1d12c81b92741e64cb00420099afa282f215bf1333374;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4d238d037bf1b76660308b06e684fb12e75f14fe2ac601ea04285844c3f479d7af3b24884a0bed25f6430120f3ca02cc0d2bb6c0c3f51a839bbabcf8441243756f532fd8ee5e4c8887e14610052b0480aba7de416dec9bf3fff3477d5e188e95e54;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5051ecf3822c6ec987812632667e73f0437544e474ea4dfab5292a293c1d2bcba5923cb8337eedf7c4294abdd10e37fa00c2e21b0987e9075f19631c373110ff0e2d32ca4910cfa08e052d687f99d40720a8c67272c210ae94b3757958e3ed2146bc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58095095c1b8edbfc5377e11ee5a7f2df7aaf0fc3c3b374dccf6c4481b5679a0c6db03605b1e8102b84645e23975f17d953ce114483d3bc5722004270dc3a621b251cd58d52cae320c11a0ccc8d8a5bb80048478e42353a0cf5cc6ca40bbbb426e4d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2d4432df94d2f2dbc2a4efbca8623bf0676b7d1e6ad9f21f1a44564d4ae53d17e3f2e795343dbc0687bcd5078954704772a90b44ca72d25ff21f448abb3b39d86f54a1b1f0369489de460070979ab9f9129a5d2916ba39494adc5112ba430141c75;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h303189b8a90dd3e90170f9793efcde696f9ef2fefb1564a720ff5716baeb1b09efcaf7ffaac3596f048b5cb72bfb6ae3551a4e8161c12fd162c9a03090b7d2b5872cdfff09d307597bc98caf85358b0a332a944dffc63872eca77beceb00c0059a29;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71ae5c7131fe6bfb2c1c1f477c26900a8c0db4c1419b9f9bc9e538124605c837b3d6bb6e6948a5e55e7093b817d5293b5fc82c92f4c71dec8a81b5c600743a2a8e18de9f50f0f00f04231bcb0ba9b1967d82a067f59c5b41fb3b6f479df14a358caa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5e6c330062f4d3eaa0bfb4f32307007a546d3dc2be51e7c27015ebf61db4e0d86abb6e52959c72617abaca852b6b5e934fc080dc617b1e8b56641238e844085869ad1bf44619517cbab0991654ce464201c3f1f3d303f5c7060e3ee54e4e0ad6a4c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba36b2002fe301c01a5076000e368bf5886aa89b56e6a986ad202d248459c1eba5feab628f74b94d62c025ba3961412a26e67e2ab7587ff2814fa57a38c62f5662960a4889e8a08d88248046203aa1358d7d2e1f81916a6ed949ce94cfe15e2c11d4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a9a808ee178e8bc5cf0250ed481d9f1fae8cde789c1fe4fac15060256bb1d505255325686a923c153d132eeb88d794bd2c29e17a11255e8aa324c1902d0e855959a4956f62089ba15ad40529eef1eff49c351bef3ffd4f7c419029ecf04cff80def;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6811b414f9eddf549d309363e61da2c094bc115e0d6204333b2b7e593fd1d5b67b94ffb6fa5bca2e10f3808b01bfc9119d1e08d49e6953eb0ca41c2d5180c068467f5037d7f1763bcb99eb92aa962e18e96ff2cb3b358dbeefd2b1cd5467c5c3065c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecfd6d6105ad26f79f353a827a5ba5f0e09ba440429ee8cbe59c03f860b1b4fd979795b7d18c87d61042a45b8d4fc2e73a0842532a25a3980bd0b15ae7e4365e6f13df0b1b798bd0b12de7cf661832ca596dee29d84bef6abc5a84e139833b0661be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd81a028b8708316f4df0680193228d50e0aa771e8e04c269d8b0dd32d1b2adbf4154cf1959109e7b501dca97751da4516ed9d1aa29515a988da744349aac59ea239d4b32398f251f948d86084da71d964448bdbea0800ffcdfe4353c42b91a1af8bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52bd9894e1032a8c7a93d8a692a1b8212a9cab6f166b8f35d1b855b71f0774a49bab09f1b99252837227af7d1933879df5a2948fab06c1b6743e5fabac274339ba947c3b8149468ae34f5c3dd983a65ae4b30b324ec339922668d03119afd4d0467b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6fc6b68ec967cb8ba8e07ee0e80e2cba3bdc1ccfb3e5815c148a5f2e67645372b00cd736256acf273fa3f1afb8e0603f11b572ad7fe077bd285c32d1b9364fdc2318d38d241cf37616f7273f6bea8040fdc0c58c18c295bd19e54eaa8609446db64;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c56918eb05585d1500e42dfd526b141bdf9fc02d9f2972baae6ad84896fadfbd70cc6038aa7c07e047be30fd3775109c2fffc99200550ca366dcb9431d569fc8313a303fb01751d3727f8bd2a50a0a836da91b582107a02a1acaf9f0bb8e0e9bb1c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93713548b8b2c108bbc7163470aa0bed53f3319019898845f2b29e6751612c8e63be9aacaa768d21cafd7413e37de4255ae3cbd6551583ce1647d84a0464218965fdb0a77805dbb22ff11c779fb96c4fb70ce171d523ef2f76e8836ffc3738fbf0db;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95ca10e28b5e757fced1eb0a91ec2e522d6e5fe77508398e7df02a6612ad8dfa8df306080fead780d5e606756f5f993180dfa901eee61e6378602e57fc3e06fa94636c9e443cbcce85ecdca2a8bfc80aebdbb86b798dab06d28a64f662c561ba3a7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he908928808ef2db4ee0b2ca7291e4937b0c08afe52a6fca26084df01a9e4830bed52a94622c7b657904f7ba7fdf6a1329e28aca816f1ee16bef9b1186de392d3169f7d49de5046e265eaa64a002bbaece0a38c826464e30bc0b64ae24a9e6fdcdc99;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86fd175785fea7f2cacc9ac36e75bcff2794505725703d4a983e583e7a42d698a76875b7725dcb665ae6a3e41264cd6b5012261bdd31cf21cdf294d398fe133bc693958d050aaa44fbfafdea47f004c4a301e31a999af650e9581d66e5c93a59a1af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2699b3848ae1cc2c675e446a9168d2fc21c1d5cfb20ae40e20eac7a3ee1db13f1a269750856f3cdec9751e7bcb7e98cd9d8b69f31ecc9551f759e4cef6d5cdb8558080ea52a11f25fcb0ab7500b5976ce73379f69579ba2b40862e753b3d1ebd51f6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90499c9996e25d58a05587d7c152a888576ac3002cf941db49ccd86e89c3f4ac1b4f4ed18a369c2a23c1d0abe5d626800010907ce1c1a3abd89ed82601284c9f8f12af59683ade9e9ab35d059a6212d38b6ffad7f57b735458f4783bc152a78d19d8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf78625bd71f9dd9029bc3cc2b96814ebde64778954c419dbcbbeb110ffe784a4fdc5ce91a8da14918819869a2f03e8b2c92aed3b530a6f428fe98cc8587559765e997784ceee26f1a9fe5913feaf2537c603664bafbbe84dfc1ed59f3c61ed57a94f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb71d713e7a7dc52128986c6d5cdcda4ecb0ca42a8384651382d0fe3a884e0b648fed6d7c64947672e0fb8d55fb086c55a193e55c631a4f0783b05602edd7035d4b0847f0c232ab4bb01c2401742da4636305a8da59e7a1b422825bea86b4dac583f0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h616b0afeaa7f70b4e2f0ae1e54a0a21f7d58d0ebcd3fa5e9c99468fa5d5e0f048ed8b5010e36ac3cef8f334a39b9f9f7a4613110db33881fc32f6448b404a84d5346f9cf5568812862c01d5543869241ddbf3802c84c742c6b87a2c411fc4dbe9bdb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bd7f8ceb1780247bd3a7c7ce0875b517500c8b96194e150e3b61d27052f06699201c55cb93fc2e15dca600192ee4df60344ba4b1df6cf8af32a40db8bb43a4c50dbdbc7613bf8185840b3e4f5e64e0efa8907a1a243cd61b8f41d7ebc9872446d1a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ac81a21c71e05a9f5a83a0904ffa9416b21c3918bce7ae681801fb037dd32a7f3e6e52f1a123b7213b778f8834a1a03b6ce4add3925f6bcbf001fa410d459e0f90e7bb3129cbfec2353f4f0eb1dd651f8e5f8ce5fe461346f0ce5bef3a848a62178;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafeb9a3daf79ad07e8074e07d249b78f9e291fb63ca006f813fb8e26db8ab6e2bfcce3a909b7410cf5bf98c31f877d62746ab7394719357a4f701d68826515dc763f637120ba3981151ac72bba5eed33b71a50d996f999f779d82ebd4b61da1bdab4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a395d9e19e1093a590d9fbb49f1235a59158719e385acb3a10c02138c4c99a3de9827bbfdb44561cf20724263596a159dcd99e67d80169dad23b9f2dc6836fb13135b991bbedbf45b7a58089148ea9595751596b525228dccd829fbfb163f452521;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95a33015b5614ae68f00055e52d7ec13ac246c49d8fa00934fafa5c081174f3f6522262c8828e14ba8264cfcbb90c70470eca1f3510747f72a1eb9da81f04351c7de01a320d9b64f76c8d5e0e2dc4bbc62ce7c856a73eaefe639b8bf667e1e67a224;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91407c83b30b8735fb16693c80ed0ede9a1b3d46d97967b3b625d1cd0a22d3810cddd66802dee3f01eb474591b6a78d910f79eba51e930e00cce31507e9269c85effa01f5d434e62eb8cb3cbcafa7976e22cee4db423a67ccfdabd7b529b6256e27;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79880fd3ec5cebd76c332bb5885042fa0212bc7333e82da210fd0c538802fbd2ef2372fe41a4e56ab2a2e86c7bd007ad403b641aae58789cc4be848da5932703199a2411560e24b2d94d2bb2a10deeea1c7c306fd321979f9ec6eada72ce92894ce2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9aacf406c6a9748522e423b2ce36a97e9326d4afd65348b22b8d8854481564cc7e48b8a90928c87c98799a610211b9c309121981d4f10c10c0c4260b98f6cd5f36a849ffb16cdaaf6f8f1f475c378865066f2e3e30f7f1bc91bb9b91efb32c2e8512;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he98a7be3120815755722465a0dafd0fe9fda7cb8fed00eb7e3989951bad2f1e1b1336387399f16594a4f5660f24cd88855423584b8ebd92625fd26328445715689a3140af4fd3ead2ff8f2fb9df370d9fc76f1803622abffd3617c0b4ddc958383ce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8da1f0cfea331407602cc1df63e8837d31988690e83d70568dc285b1ffc6e51c4f7f9346a371859483bedc10332c6ba9f0efa6d9618660b4c2145c144c6d7743115c5d44bf1ade89f412cdba64df396e32be61c8f196072463b61598ac3c7b57ca5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd24ab77779501edf76c186e108a166cc609814a106b588b3256bd784ce8547cd42136a7f349b568893c087806d5fb64131eaf467710e1c4eba711dbcf1c734c80bd825c43215f942da0a880ba1b6edd25b9428bcde77b43dd68508acaa5a7aa46b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h528950ed2e27a0610e6e4179ee868543acd073fc596ce05f2d2a8d516e5b56175e45ad36f235194a1fc65b96fd8f78ba2e8e6ed663f2d36400df712a56bbb66078d4549ac6cfbade3655a76c2d84f9caa7f06cd88f4830e385346cf15bfec31e315e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha14f1bc2619b3e0268ef689338cddb115c79db3d40d187dc2b54ee8376745945247cc494a345fe167c2de77c3475571cc53226d7ccf5d389bfa6306ba43bfc7b30a172218262fb9cb45ef9cc088e6238a11504f65847b2abac62939bf9484cb278d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c471f93ec6ed6aff37de45b4d73533c611961cf24104a313b7dab5af8151342564d101ac591939e146185d29496bcdeea048189c420ec5e817817d46694816b824a5dbff837fd62fe7e8aa564702d1d8e85f65792d3870d8599862589c3243989bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd61b23ad74a56bc7500245f5d69f2d3397818397e6cd7f03d58e5273f74d9a9d1786290f01e24a046f7ef28cf7e417c53f591638a5b55a825906a666fff8a6190ec68615f8b952391f30330f644b403fa20c6eca4495621e69763e776bb9de0709ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h615d49e2e6a86716b5d85627d014b971265af0815fab8e120b86231fb601b93374258d3baf36acedeb500461b8b4c3b9d9d844b73928564dd6039e708d1396da2b4ca38d2d1a1b653c5f7d74b84f7ba17091257cdd31e7ccedc3e683ba6b37d747e5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8be22421e1f031f36a1b6f630eb151c2f966eb4ad261cffd30035ee7c24ad805c41a8c40fc24a2176098b646425766a2de772ced151c33e306fe7cdddb907f43a25d2f147e77255e779a1321ea092fe744ee60c92b47073be5894f999f4a0d85bbab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39e983e7d614f5f97b90b3c535b8da900cab1cb394d470e61d127c437f6a4172724850b44f11ba8f29a3700d6f3d0c87ba519c5e202f62dd0058f1c0f6b711ab05b62231044c8b067fdc187ffe513b12d3fdb23f00850f558212922bff73d0e18322;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9990868c598955aaa7ce7dcb53a935f1618471738f753373b644b432a62894645e0a7085a0c36e2bece26ba5c474a918588d5f299445eef5e89128de9a3c540ae610b9bc70b094abed659256e5b4e1fcbfeb1eb9af4a45b5b95a62d2da8135accb6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47e2a1aacc651e1c0581894f8b4afff4614c1f571311d261090b0e89d0356a6d6f7707e8f0372dd852f2c3365dc92998b66c3f5bdf5dfa4d706398181036f78887cf2603a2e5d349b1aa051a7b5e468b11f3b0bbe9ec1ac40df701aa05a25378547c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6778ac69447bf842cb441aa7f34412129c90e50569405d9cdb09106a2306e8b78320bf5410f1a5c3e07f3d98cc6de5dff1485f2b10b5424a204a071100b20f8a26248c0e213a1f57b95d8f3435bac37be8e6c821a4c797a24ae97cc9525a6cc8b4e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc215235d4e44764863f290519c29b106c0af435f53f0c7f7a357e933712fc38ce2368e58e8cdae7ea11f2e44f123d24c8e2c6509432e7dae15678c937c76b840206b3aee34d2f3248edd6da17940afff57bd7a46b6c9ed668c0f959121b13553836;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5f58970745cfa61c8406d0a43f342a31faf872eb41f34ba9d27d6f9544effccb4470aa43c6b08ae777f34a63a6077c74265749408d4ddc2dcea124d8f6c61d7a85e97333a0bb0d06d1a34a02fa99ff634bcd41e47be8d2012cc61ff0441bbdc58f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f727dbf5a9d368803877744933d5aafc395fce7aac6790c9548605059cdde26513d4311cdebafe04f640a67ae774d00a1cdfae0b80253e6033103fd55105eae79a13b3fd8ea6a411c853e624edc09390ef0e06bff1594a091058161fb08f43adfa1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc90863f7891c752509992ce05e4805dd5bae1ecd2c70acc7e13f7a689c8db94d75fb709cefa8c31376cd63a479748702f1563789857eb90c90bf892f5c8895afcd75a26147fb4321ef2311bffbf324613e2d81aaaf3164ea88e47e45d25fae74801e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7617e3e0518cc0958e03071edab503514ff2ef39fbea5d7b154c9a36804aef5a52be2482262cc89b25b7e9470faff9d0cd85a8a9ea4edcb1452901331c2ac47bb0772e349680705eecd4c60def5e8f9d95b7a72f94756dacf81fc985cd3e6871660f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cbd7c6c944aa1d1b2810c142f9be8e8d22de071af13ba944ddbb1fc0340e08aa70733ffc6f18f71eac2d6e3f2423f2529111601d3749a82a13807161f1c01cc78dd952c63a5fd5900e8708eb27446c0f86c70011d9ea56426bb18205c2150e5cc99;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff05d4a22baf6b33a7fa4a042b295e5763fd4ad092bf2895f575abdba435935a4a58033685137cc39a3efd8755c810f4917bed1c9d6bbb77c11227be5ad7762a7b7d8fcdf6f4cfabc04154c01e328d1ef13c527124517f4d1ddf693a41c0ce92a309;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0987403d9cfe06a1e3d568c0d5e8ff8f1ad0f2049849a65823e7bf20249286a6e51867d73199bacbfc09fd71e49ed74b4ac2968199e00f31867fd9785677d9d44befce87f3776b853bd7f7ba685d49f67b0a4c940205f1df478f6e292aa9dccffb9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h245b050bf6a5c0131d69bf7369986305a896459f203cae073cc7303d7278e18e2946ae01fbfd4933816e1db14241fc0cb60c1f069c8cc5b96fe34554a7d6e44d22c304943bd2dc25580decee97b316ef893b4efeeffc36edbe9b313219ec407830bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ae45c3c53f9b4e407ed763b40de1d6b5ca2b4e129c8f99c9467619679fcb48c0365331843822069b163900d14c5f31bb95cc63c5e557d7b5063815f597ec16eb5cd3514062a6bb1c3a4bcfee7c1a5f8a67e8ca85eb65671bf5f00a6229f607c68ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8132e39246af07e880cebbb6d2aee94e509fc30f4e73eedc0d06cd6c110788cba681e8ccb87c12b167c966b68e148072c68d89ff12078d658642b5dcba9accd79ff3975ff769459ee6c1b9fa39a5ed9c0f9d5d854171dd8cfe6345a37d502d00ab5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1728ebd890ec86404b7f9273611c34bb833101750362c4451724ef9442b8558ca39837f76513329f7bf8db6c1931e3df4c49064ab559cff9079d086dab6bc645b5953a5f4ee9ebf0e79655627fbaab0e7fe3f98c2d0a3d243e5a4f5ff34881ca54c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd9b27976f3f8905ca752ff3e3be13e894cba9d6af6c0c3d0a4614420ababf6f36ea8bdca2122d4114099cb6030b893b95bbe4e23f7165e1cc02c84a4716c28c7284353423f41efe3d9d56207468b05a804a4191e51b97f555eba1b8c235e80389f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h382066a9397fe857df55cec7d85b0b34d39e1e611954defec213f5bae9a8cf77bcab83c37f911e787225fe52d4ae976bac09bb14eac99306cbbcc5724d22287f048750229d2fc3ef3b545698251917f1b4ea38792f763cb6e198721cfb5de818f53d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3fbd9af3f2bb63a0662bd5c665ae02293bac7177a565bb32f4933a7533ff702ae360f175fe92afc2f9fa11aa6ac13f8cdd7017ac8e8fdf4e632ceb729bc7b11b8ceb290f636bb968ae3889df08328bc439b7cb9ddfce765316faeae24efe0e04a77;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83d342af5e3e92eaebf2b81f7d5c3b2fa7f5b6a8934905890965aa3c89376e59adb4134f8a127b2ff1eabba7cac690eb2665420c30225220d5bd5151a5cc7baeb7aeda486d497f351eb463637c18a724d55954056776715c0f3e73d419f928e34b0b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc535dbdf9c04febfa18fc14ab22cf5d397f726100d9899482b0c7702e9e6243f6a7ff114a08830044a6d0a4691a42423debe22c0d352e35f368dc5fe07dcf22eabf23cfed0d99007df573c1ade68be66ceaf622ad679b1323ddc9a2f90be302aafce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0bde273e9e9d2f6295eb199fd341ce632b1011479d64abd2aa78591b04948099ecadd4cf9ef17e786563f369e58f04b2a4dbc6e3a696752578ec7a2ebf5f6c0daa634527552d5725439afd4b281277eeb424202c9f167dbf3eb3223bbb4aa6f39ad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd1cc4d9bad4c907596f7e4b3736fe5dd3cf4646da1a72a48f8ff20b8e2ceefc8a48679b27d49cb885b8507b181173fd8baeb73453b065c948449fb5b7a5c19d78ff310b941f4e8a2b0c3c180edb5c2cab6d30db5ef0c10c4c022b7f6e94f3429c87;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heda54c9a17e33983fa8845b5826a8ba2c6fc3e02ca436463b6ad04fae89bb8c7adf7b90473e9984aae445a340151ed516b04e6b3f85773984c491e610d88c6c019645105283ec65820ec690d8576a61f16a327be037464af6575446c3b43cd8cf8e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3205a1e7b852007a1afed1109eed4b784eeb76bbbcad701e2960da8c43b1a7e2c0894d814aa0039983693080b60006f0380d080c7732a436144a9989c84ec8d9995caad8923d3673b58cb3be542d485005d3c7325118b272dc11b4f257e0244344;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90057d5dec7292765693680e7a5d1f26824e69fb112fabe82d9f49d34fd956a18adc07a361e642ec3a84b81f07c29eb01b4fe84d603da9b440d6254124b89da39083121ea017e2252bc91d251315fcb6ba93de54a4e1c10aa4c5be5f1048d617acfb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h895ed01d93cec05c9f62e24a76cf59d08da9063c2276be4701da68cf6e08be8daf5d08ee1552c7792f60530e4dd17a8a1e618db7867189047d64fc39dbefe6b92f789bb13777fb20c8f551f8dc81a7abd074da042b565b7dd946bde1c459f75b7633;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1eed27ea10aa12ab43725b4746982b170a0b7634f137b2e119482bca009078bbbb1d3ed99852de3539404a2b68d6a108d9900b618ef9a5d56d5a900e768bdfa2a7dae287aff170ead5fae81b7715525283c491d96e6ce855288bd3ec552025349eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0dd905e621d75bab8633498487fa813f667e38c9e4ea5888794fc1fe5806527e642096d99e2ab0a7f42b8a6311241dcb9d2ea3d7f923567c114621e0a6ad9ffa5236f3de20d250c9bcb308cb54560f922650587a5d6e76378513f802f07e43ab500;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd896fc15aaf08e5f8639b28450b30c2733c8518f41ea5a4ec5b1b122debe8773ae20ed8afa32096338632b6887d42c81fe4bd8ec154dc80b3106ea38860e058fcab01899aeb667d2b9a84906f818a81b97345b4eab6c8983e156fa4970abcb7cf138;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd221a961a9c65c35c3ae051157a2130bdec18249310da48ad09689d3b9d98c970bbf91a2618a9261bd247e3ebbaace4ab325ad5c33693d29b891b884a04ba55937beb94757ad31d8bce5663e7cc7aa6c5651b895e52b5e501248dbe86c2616c920bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2cfd641e5cab434a352fb70b437914e2e7ee40a16565695db919068b3a6ab2e03be4ea1e854dab5619d31aadde3b1c8ed9f9d080c84b625eeed93bed5bce82b1ff2d11280be63b8faacdecea209a587c427e5b57a124b5afd9d2d158dba87d557d2b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h959420b3267170934613da86b5e86d2f8be94a50506acb8add5c2ced8daab981d91fde70721e2db605174d26f594593f62210b600ea598b5fccb88a236a5b79399657a4626ee7d1845b2e8626388dde2f644e7df8f72298f5629b477c52e95999009;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf5eac50196bcae4b6f8a723266128f9c64a808732676156629eaab27766d7165864bb1513aa6564c795bf65b2f14c7fe0590c27bbbcc64927a795a2e0cfac4c986f8d8ddaeb45fab55d67682f5ce80e36352fa309e91fee45b64871ee32324319f5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61cbc30b6120f7aeee1e1e8509a0a3f359e35f35fab472ed33d10546452db2839beb21fb9cc8044cc5e980d203974eba22913dea6d62b33e6bb5f19946677ea9a32f7d8ebaa4ff525d06521ba1d57884c5425bba0e39104e945ac74364f9590b46ed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa62ff25d32c2541c4a5451e21a3a8957ef268005cd984dc1b4b8d119cf08d26b3175208e3a1c3bb470ce80ea03794731cc8ad96552c385bdf620cce812e9cfb293c57c89d2cd4eb04a78a870698633764f56ad1c9edf055f39a98f4e360b709b2b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2be1505c4a4536239bf4a9100247ce99cb8133a4b16af3039b880fde5a9aa485ae8e133ea5100617ea24dfcc68bffd84a0aace9a2dcf418a2c08b20b30504828d9971500130120eb4a8a6dd6863a1bd8b5e22b42ae5bc3d2cde2a6a0225cd0df2469;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94270b57ec4c9fbcc679bd7f4d9b6ff2fcf4c3fb03183dbd48aed8c5a408453559cd974371667d72a68d16889a0580b21725c991340573e72b6cd3bafa69e2391a8a6674bb4e6fb7bb7c9db27f2b39da90db2e05ba5a18067190d490842ba10ef65;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6ed9f49867f9750b129aca77b44aa6338c306c1a44776e6b54ed7f3b02e586a20c11f2453e4d8ba4f6c29f5621ba9f399ba6fab871125f88e8132bf024abcc294638611d25d15a718b381c68b97a25b29d385b983719fd5c440bfc311aa5dd8d8dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha287b9373b338b66a2dba097c91fab42985d834a00157e32dfd23ee125261470b2faefd06e02bbd65572cd85f02a2b0e35349b2b0b9542ca8995ef2dffd8ca83e97c6ef3a7281c1120a419a62a9d303daef66e06a08cd0302ea41f9dc57861b422bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd81c31bbd713f8d119b5be832e1e73921bbaf83874e843808e3cec15c113d4d38fc31eb51a8dc0619c060c954c516bf7369d4573560ea6b9c751f9e541576c21903f0d223a317a6d757c7b17a56045658e0ed01d3ad625de9ea71047154db25986bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf705e3718211fda7d05b9ce3540a1814f5bbd2aac3e24f8df311ffccc9fd40088dc2109e5bed92a06ebee575d18795dc129705c847efa7c1ece5455af6969d3bd53c81782616dc75b753f30adb33d0d3e4ba5feaeefd0e7749a2e047fdcc36c16506;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h745e9707e76d3bdbf0f55e17bc7a8682242fcb07cc93ababe71c9e33dd57204038086b86aafc3e53a914235a1781355a194cdcf66aa97d423ada6597cdbee000ba7806f571d2d42fba5d5f61236d8e17ea5b4f5c082388f70e90cafe790fecca50ad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf10c610bab3a35fe769093836caac256422160f8b6015e0f9d0950bce8dd79ff22235ab21228dba7ba9d6e0057673c61f1c2ee49056c39cd1fb83cbdbade07fba94e1d553b1e313d94ea7b2aeb9bf53f0cafa6474e57d6499e8809aea7b4bb215eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6aed063f3729e1ac9c86afb6850b61726fd24a0d17225b044d89346bdf143f8c606a5a8582fa59e40af8d8abad26a30cb7855c8219f885858a3b7d67487c1fbf4d09170be8bc56bd61c6b52dc45e8860094544bc661da72a43ccfe7a5f82a61b5205;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91444d1a93eeba07d42f26982e9e615ca9b9e90829f6b289f9279c14c4d43073923a67bc1cee2f18d6c6bb9cc1a2b7be939cf3c68859f473f588348a1fc3f7d8b1ad771ce884fa69d127254a2273781f375f34c7c958a4e019e25b7e5c846d65325;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd624e0ffa0f30d15b8923db3b64e3aa94fb5e46fa07f91560821a5b6e632fe819ce465bfb9aa7a88f66828e8c13852f87e649db8d41defb852c1633f2c690005f2db3c237beccef8e03d35aa9824f9e53e5f45a4b26245a066cb548c341b15d1c955;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f443c4d279226c8849ace12048c98764eb2675e6edfee4d72ba641833a057377fa610dea238de9724a5ab0abac85f1aa8050cd2b385948d3e147d80f2e12fe881b140699a0e8aed4f54b2816e6501b196ed21a73b86f1b710ec65f3b515ef7cd8bd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb49c6b8026f998fdfbd0a72d831d7e98a6c819fc0613f03c4e2600430bf990aad67d8e977084af4ad7e602fa2e8ea64943c0b0f508c1d59f844a4f65d01231e21cbb769327c928b3c8b24988e16f2fa6ac231337d3fa4959c68d254df536607b32a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f1a80ca2f438ddac8e73698d04eb4857fa5d0349a3e793bf43c7eed1f154097e5d4ab9d20a475af62817bd876de248d80fd9ff05d6f86b76eb5ba0d2f8e3761631c057b26ede27c0a927c3c28c4f921df1d6f95281d133105ffe4eef39981737542;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ef5f586cca5f94d8071a7798ac1bee1b8762e1730e1e3be24009a8bb14bade9c38e55776c85188631543443387bd2124b93ad088ab79514eb3c7d6a64da00f7b34d2770f8dca45aaeb19880218dbee750dd23c442dc014bab26d8c6efd00da81d67;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54c607b33ea047fe1b85c12e7ceabaf9b1a93dc211176f10a47c8dd14e3346be810bf9f92ecb7f112a10f58088fe0383730ebf7dbcf814ff4518edbe860f167dbb8c747ae5327b257d8f1ba8db2c7766bc00567c53d82222222909ecda83ace188ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h446439d9651ac7786d7a7ec2a6a6a3538425b5db8b71237ad6daf1ea6deda8bbb03e8d8c4b4b3190d69007da1c69661ff67d0273328aad865f133d6c4771d771e8d06f7752c02acf7a587feb478348d44036c564aee52eb057386d3de48d24813ba6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e6854e39d268d226adb8b5337e0d3fafe9eab9a536ff63b3ebd2b597217828a850c25facc01afbc4eb3a9251d7bdcd9386efbf20d9144943550a9197a8abe819733a7ae9ffb3d72e81ccd34793b288b8e51af7d35a71df90bafee4c6f6382c91981;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3e4befd08515f2d9883e98b01b0b64fc109a2e3d5a327aa70fd104c3bc42738d24fe2d4b6f7da625f8c9d4d4dbcbeb0d01b12fa424d02992b197a675a3f0e3ef9cc596679bfa4fe16f36fe561b73fc3e307a8e5ff882872dddbdb65cf4c886b8240;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95d75f63e0e0c75d20efa9738a81f19eb10bee919397e3955f3fe0953c7aac58c2fcef16fed784eeb51e42227978e1701151129ac4c121c0cfc90c35babfe67e39da338dcca805e1d9627afcb88ade85a87fcf6cf13ed3217dd47d21ffaa5c0e50d6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb95e0685982c63871117e6f443791d08a5a7a401add0267e5a8cc6c16ae4d81f46b6a7585cf03a0e1342e9cc16850e3f30993255751d3c5a0e482961ebde4ea3ff228cd555094c11dea347ecc6036edf97a478d5c9b310a2ae2ea5acee686673a33;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4c14f057f170a81d784fb9ed36e957528fae7d81ab3d14aac6b44527aa6830f5c0206520a75e480bb8d6d6c5af14c57fee0fd7c27169e51456fd5d40234976b22c1a07181a31f92233b1e6ed9e9e9fcd999fb35da1f1011f637c9e550ad6e8bd372;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22d7c09f872a5c5c1ecd759fa9dc08a2f250c1e66bb85904a2c2bdea50bb088e136f70304f3c938ef786e245473245a935f4222d5cd5f50799103ab72ce5012c848e4d948b7c3b5062eceab5dc0627a57a7a6b05eccc061c42aafe7ab84501504255;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b13e4bc188cae20921f6518903cd840ace24985beb8e8b8f89e8be5216dd2e3b2158402005c7730abc6410a926172978cc871c61871097d6e22302779558600a9561e0a50ef5052b4acd900f801e541919ab5ad518b699f547b91ea55dbbe9bf2a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde9e1798d39ab4f8f219318e9db6d890c7fbecec8f777e63308a06ed5a33fd884ea5a2d598d00481ddea5499b1228936f35eee7e7dfa5ee582597657beb7c5b2c9598709f4879d757fdf1d426308451eae20c604ce610b25d9587182fa640830cc24;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h258238a87bc04029d24f40d50636f9ab0806a7297cbed1e0f3021c8bcac713a41623485a408f75b25e6f7d58a706eb2530f96d8daa3a1869bee83fa10bb0ef0bd0f80da32bdfb3d25156c42fc44395e7cc367ff6b37f7bc47a60555d3c634a590831;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha55679fb34363f2b649c20be5d5c3a0cf5c811907aa7903c912739f5ba093e2bfe68a300e672333793a978d6c5418fd887a2a2e0aaf52389494517fa5a3387896759dda29c890decc7d9e7f374027f13af89861f24cc68d2ffb2ad99b9c3ea4f9386;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h589331ee46137f6cdd698679862c08b4e126e306abe0909c4109854e2c3d77d60bd90872c413e456ed6265fa08ac758b36b420824d888a9b5da028bf416b41a1db4d27c24eed7df84fd81f1cb354f99befb74fad31198cbbe23ae5167d816e0b9ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h486069c2c1d4926584b08bdc591240636a2434eaedc69f9a85f0bbbd502ffb5c9498a0ce20eeb249b02b965ff7349b2f6e9b7cf0416da87a3c13945b58e4fe7486661a7f52edd43c5937e62615fe6d230cb0b122cb582e1843b660b81276ebff115a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1e000318e6b36a1d52710c26be488be03b71618e4de93cbf7891f7d490dc751857869851b69cd88f9da6dc75e0a204f01f137034c64976734d2eed7fa761717267c7f37f5fcc3995b3540d41b8f3caa190ab4c634512276794e0ecb67444b82b548;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13e2906568e941bf1952fa7f49a7abfc32e72e4efc23b48add0ed93721bc8b60c6ede3803dbc4bfad58ce2a1f84c9692fce476f3553746367d7a79257f9a4e0d58a7a6930b370ce2d4d01acc6ac1ce3278391cc91f84e19d8c07e48bf5f3cdbc35d0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8de6ab1bcf6ed281be25b6ff940b7180e28ec324e8324d7eb9a4285bdabe07bcd97f81f79508ab22237c120b421e2e561b71eec513acaf47486135c6cea03d4aa62e17ab1e1232250c73e296496ccefc8d8c273fd2fb4874b3eb406c5e3db7f42e0f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h940b5d773f01c46c4ff38ca711bbff926ca6c20b67a908c0a0238cd6cfca70031a1ce0af82678de94af1c22ba668c5e0552afdec897b4d6eb829426a6918ab46e45cbb0b31977a1e138cbecc79fdf1c744c3dc59d907e9231bbf850e3df29acb9263;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4bcfb225083d5792541eb991b8d53cd6c47a02555992ec1ba6f34c232e5789db4151ec0df0704f26c16ff0d74e15c4dbe46b12cbd0a2de8ec81168ce4c77050d67deeb54278ec9554c81589f35a21e59b847f8ffde7bc48ecad45a84867c7d8cdc32;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec2be369f962f5d93ed3637f64e700590a7a61ea0ff5bd328cc5a928a9a6706ca7bfb148966fe9ae0e9481af840736cc94cb2f787b71f1e8bb5509ed36cf38b2962b5e8cda55d8532bddefe08167b6476b0dcc7ccacbe4dc225edebc2b1a9e4b73d3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h694da387da76fd5903a2fed6b77b420d80f2a0db6b3703c7a0c4809e0e470e9313cfbe894e5fba70b057bf5ae3372b8e45150af3dd0410e073648f6490bbf17cd9d0a10f8da7dd63894fd686b3efb0909baf6245bfc5c3b419f754ecd8198784b38;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6afee33b3b4cd922fbb50b9c3dd4293b0350848055ef12aef6a2c8ef1f76cfc1f006d48a474a9eae21c26028d856bb980204f18b6f01a23ab8761c480b8e228e0805adc16a4533417bebe463c6dad7de2bff3642ff466cf02062df30e4d811c04c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h347f5c82711ca8120c9093192012f100e960e97931b50a9707d32141b73a97de00f8a3b00d273ea2fd8d2e9596cce4ed07ea78c12cf3df33c8068d1430b38f823f85efc81a64223756cc48ddc60b691eacfc80c9e042f27f4c004a0c11cd3c331a51;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39855082479d6d4ec1b85f6766938d50aafa39da7e82d0f1cb6d6d424d972f94315881e05ec3e715ae69ca1255a011a42770ee3bdc74cb2ee2ba70412d40905c64edda6cd4bf1cd7d1fe71b251da74cb98a57f0c15d4f6ca6ffca9027744bf7b616b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec3fe50446d3dc1a42836755829dda2c03e49b12029fcabd2a343a9453e88c2708d1370c40ee491f66b8cf5fd95ded6857b8b4487dfe60ee1584a5834ade728657c2e89c2f6a7c802fd0a1d5eb732ecafbed705380ca64e6f46a9dd520caba673895;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57b8afdde98c6ef3bc033707b47d9a27dc4196d76a03627002288a76024a4ff410d98fefec942e9391cb8d8c623cd4e2838ff6d2fba2b73083dd75e99bdcaf41df3363299b6fd4178147d0668ee7b33ccca47d540d1c3a036e7b1fa75309772a34ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d9baab19d008db52b28062104e8ae9d1e063cf8e3230c52b11f6bd175fc8a41a8c7eb0fb156fe4d85d4104c18bdb056e1939f2cb498a0bd55bd75cb73bb7bb39fe9691fb81756ad3430d5c3793cd620acb70b01d3a9caa7d3506fcf3fd17abee205;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2454fdeac3d8ef9773a14698100f5d67b28edf6926a365a8445f1face27b59cf9fe0caf590e3b4c0cbbc1ce94e761b65437ba4ae8fe607e31f1b2d524ed208f42a31bdf768fe0f03c1b96d7652fc9c5a24310d82b8a1685bd3059f9462d9c48381a9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52bce7aa33a152b379e8a21add9ee90b07fa601030cdd5aab1e05d8816051aa361f083d2fb3d0a5ccf10680be845bff1996ad33bf9458dc0162dec7f06121f5cb1d3fcf98e6a1e396ca9e3fc21d7885266ebb58f923924e61f74b9beb31170632d40;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a47a9e92649c4d8095d13593b1397b933614276648fa96c18ea6f4372b3a2e9ce00d92d86d7d8394a4d34febd6bfeb005adf58f00085e30be9fb1e76ad8c5a419506a54b30add418b1c36a99234cd3b72f4a23a5f33c342c3b66bb3fd20eb649ed5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h68afcaf6c58d53d882897903a45a3f0519d6e08846890a064b9e3e0e9396885372c4c83bc51380c046dd287e1f5bbe6f53102e9656cf55eaf2636df438df86f42492eea24225f1e8b5804e7f05e55047ae06c448288816de1228457dea6bd5ed4bbd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h810d55dc7068db78fe993b66d30c39554ea86b739cd3a95597a49eb6ac5bd2341c643dd7a8483619c8293a9c44f03c476608aaac94f670d8bc742ee590dfb00f883ced4d280c25b9c6a2e461e9f652303109e6fa5259d14ca6ac8d0090a2735f30c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a07335712d4da976b27a33adfa44b885e66672e6dfd01bfa2293f22b185fc80db333c801238170cf54741979e111a4645f753f57859a4af826e726f53ffe1cab34902bfcda86e29af987f152b2ef44378841a04120584b33601d4b5dc7366c10fa1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95e432da6e8e577ea826db680f1cb3cd8a652694f180380f26b33e92b869c5f88bb52c2caee5bd8fc2616a9b824ba9cdb5df8e448cd702389c414b7aa635eacc254c7405e284840485970dd2c92f649674baa18929d5f7e45e4939d6d4b38f0b8681;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5735fbe19fc5093d4536fc789c72febb6c9cf21216edf42831ff58e64073f1288c8cc8daf53d5c60695820c1e8a0a64212e0cd808707b785e9a6f100d2b31394eb6c8c69e0576317282b4341bfc865078bc032d2a3385f8bff4ebdb930652d775676;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he93e266d571d23b98091c2dca97b6270c0e5d64c20d2eadca802de1e0656dab748b7ec643840495210dc3a7e908003b99e524cb4ec9d97ed4f2d67cedc7d719ceca8aaf53a8fd4e4bf9b0ee244bac3c1f2a3aebfda509642b3456e487afb2e2fc50e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ef6809ea98750cb2af44d53d518d77e74a8be64742ee244475e2f432aabc2df87de24af112a1223f5e1706eca61feaec5bc8c0c77f4e54e387c6d9074238a56127ae9718a9782170476126964c376ee4a72ed15a9a9403b8ce522131c3b2046e361;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h524613677ba90abd91fd9abcf0788827114fe10daa3c86cf7b1db91f236bf8fb81ece739166f43e481329acc94345983db8e59d813a6041c24557490d701e209cca19b03f07fc7ef498e1c3809b512cc81797717f93c5cfb6dc6819b55d245f41b9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h511134fb42ee3b72ebc6e8edfb7bad74be050f242573a0da265d6806e731c82a4c851f32f0d091bd30cbd9e36b26c32a9ed5d0b81fd3462f44014a793ef67d4ee753e61b19578aac29f2db0642dce529a81f4d889cbca6ac591d1f1870357e2f2f30;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a1a81eeed6ca8e7c90e7663772940ebabb3a24b5a4bf3f42c82cd395bffeafcfcdfa951a031e4706aaea6bd469b0dbad62c7cdd43eaefae138947479447f0e5561fbcb4fafa4c32c66441401aa952a96c13980d0bb16b3c2ad1cbdb4e59d19ac;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e4ec285e1f24b92351b5ecab184fd1b36184c311fc911055045ae51fe73d3908f6e8cfd529eb3efa032f8f2e82c0eb5768f0c0ac20bba6d0af223300bb85e9a19a9f0c0e2ce11cf8610b70ff2c397d84a168764d1aa073f79155ea139335acabb82;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36fae831de4bc7cc4b6e610b1024604dca78cc9cf1ab50258ea8c5b8eda27f4c5b03c82ecba97e912b1c81d274fd78da9aecf079d9fbfa0b86f2d0cf4bccb317f6e20143ddc086f217364fb2c9238960e71a23dc1b3adfe4907ac068e4432b8106da;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfabf42b73b8ed14adf1b096b78704cf64b2f0b47b7d768405309ec5041e7c55518c6f60c85a23b358e868108dbacdabe70b521c9c2282f6b8c666c4acb8ea42fdb9004d29873cacde546dd91b856ff3be7b4f70bccd222d7a4120126fa9b0ad6f46d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61554b3cf2bf2c8eb6f595f94c1cd9a74788a1b330fca5bef4c4d315cd810765b52af511e2dc493a47f911c37d654c8ee36d023789f8c423f2619645879056639b24f43d1359eb719e0bc160c0e9a4f45988442603cad29f5b78208d19715f8c506a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6cc8383218a642cc43de752998b1732cd714fc356058a0ee1f2498a74769f7e0e55125e0586702a3aeb806ac07aa2f947b29f62d959e2e3283eae5c3d354ccb1fcfa9d0035e6be55c3a1d247e5ee633e45d4b69ae8042b88463a8ec447c2d6ad3827;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfae3e246ef4b3d911d98ea476d7402221c8c91d2aabacbc70878298a318477875540f1da0435e95d96235335451597a0c1d3df20c06f5c8196ab4a1a75d997597e7141fb20f937e88a17a109183361491125cd143b394be7a75c87680e40da522b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h111f951471bc95d3eac99c1b9942a3e740efc4d33a0072d505790ad303ce591032304e0b7230660063cac5522974cec543d457036e30907178e9ef83fb47d6cf948f97365d0e97214b6725254c02b1ad89b7a3566c34f728d21a62364fff1ab5ca66;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa95e8ed21418fafd6bf868fc39db1f6994539ad898886a333dd9b540aff35a5548b107b58285f2ff1a51b9d15f49b51240d06faf0a32d9ca4266b920d11c003a37384136cc07f6d1b977e408ed7c568103f1a8e1e3a88979f985ea09b7cd7c60948;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86cde67070fd5cb9025c0f820b382c4d48bf9dda807acad4fe3fcd97a630e091761c1d34124fcce4c9896644d08ec241980c66261d5dc0808303dcf418c0b2f1fde39ad01776217c32e81a1e67717d3ac7575ea07ef6afdd142fd01086ee0b7f3bce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd52d5ab6d08c2cb7ed89a9760bc832bce00ff7937e81d7855daf346b6dbdb3c653ec088c4c9641999f7df52def2f585feb38ffcb14240bb3c79b51e74b255a92c185a7b0904377ce8ed51d2ccff0a1b5cb4536ba295e1c9369fd153b2e57a4f2c21f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had58240307c6d9d48ecb700e3be721d46a131f5421c099625f57274e087aa4593d7ba327dc941912d5d585c6f6c1125f0ddf25d76b267377e52a9c456869d55f32af62a61b818ef8529c6a31438163cf799aae06f89f23ed6addd045a7318487cc49;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he17b0bbd7d5eee0058da933156855583a31a01dbb2659e36ffb8379165b2d3ba58ebc1e2b5ce1caecccdcb44be719df1b3a55c55eb7035257c6b865bcd8a45cb447ee60a741e5331772880404f45a6b0b3f9c607eb67374735fc02096dc8ecea5716;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h253ed966258fa6b2d7b4d385ca0133c5c419151ad5f044462c735a231ac860cde1867cdd23a897f65e816ed199482d9f14253a5a9f6652b7d578d88c5627b7c41ec64f45ada55fdd1f95e9ea18b8595e345c615e8bdf910dfd9346309ab79d004162;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ecff4fff8cc6c1947f6e888b6457f80e5d4161598eee419e38e82ccdf9b97dd07923e04621285afbb5f07fbb3d2e33bf8cc2e8ef99a700894de711f264ce2ca113138af142a9fef40f7653ecd8dae812de780ef54ac07448e1334f50097ac4c1dd9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h479944c3bb3fdadd2572d1223e0d83a9069bbb74c5a81f137cbfcd283f945a0a329ba0c39c2ecfc5f39b781a10099dce3420d3bdd1f260903d14e88a56007ae827e860b18c2dcc2bf6e5ea0299c68d8cb44b409941f660ab69b040ff07d7e360963f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed99df1f4ff7b68a86376f5930e7a905031018992259631123d992dbbb388564ad0b39de30dfa20b78cccaa4436d35053820c8e0c9fbcca42a6d8acb3f5c829529cc6f63c49cc6350456d88fc1b11dc828bfc68e6c99f6ffefa7da5631ef95253178;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd4aa42de2d92773c7a479f358374a6efc980b4400dbce9f4878d9f323775da21ed37a19bfba0bf7bad6f9280cc94ebc628c62b9519b430722ffd14b83649950d53d659d09b1e2fd0557209b7870abbce2d1b5194d0c1fab5b5e9d1f4f7989c2eef85;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34007be3910abadc387633191ef0adadb07d63f4535d232ed7e3aee44a57f607f1a0a9e4ed5c8d0164d99d43a75a812bc9137eb2dfc50603055e298aa2dba61f788fdcf7dc886f4362c69d4d39f4f144f5ab4edd8eff6a4ed0db758c6333141da525;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a2135c6b62b36a2118cc49a79275d660825a72c52b408fb46228760a831e2820608e65f427d114309d7fc52cb6f4f31f1f3f69a946cbc3cf49016e733b902a2cb8f7a85c4197bb888b807f109f08f5db1b89e438ae8ecd2c3d451f5287ce4321f15;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7de4c64671c3375e0ec592ab8ffd5e6f678df3fdd8bc0cf190d26de2be712961b8c381c19b28cbbefdd7ddf8cc576fc56bc186341f9684a989db3088d7db88e0f60e90261958c1d47ee5371980b93830ea1020b002aa7e185bebdaa7aff2fc525262;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h859b8b141be832fb47fb957231b8d5c404c8dca1a50704f8b4b94b395a010ccd0369d2ef29d02eee9b1629c15eb2888290f2035dae0d1b7aa83ce2812086fef5cf5137d5f7e67a86782da11644cd07d9689ad0393d1ef1b045fa84d8774f67707387;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95c493246fac9a23464e6166cfdc28dc5c1f9d234b86b8b9b34fd77087d85486b6e8860dc829316fd18eec04656606af1c8977579419a3f0b43b5748e269915cd9e0dd2f0c745a00d58254713562a9ebb8846fadc0ba6bf92f7e4f31ee786fc7c533;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bcd25233d18e408c59f6663c84a5e38ca5b0244a5659723764598084255903104878a1834986241ec63b37e4ab520b6a5adb3e454edb755745e234548cd52a1ac956304b55f1c6a3f3e6da3b48efc25ccc565d0155c6482af945b5d5d5c926eaa79;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c2209ac32ce03f1aaca69ff1878406330b38c03724b99eb1ac0007f0276ca3bd94eb690f57b1210ed35df2b7e99e08efcd4609b776a8586669d1db1953068e05a4045a40b4c654374fd103afb1425f863499c31451944c1879b1e66160083aeedd4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf604de53dbbbaf17007e4e465dd7a4a554ab470555fb0930607cd5f08bc1d4064326169c7564f934d2394ffb690ee4ba8afb525ecde9c3a48cecd615f5476558211b10adef86e0bfd1707db095dc287b4a475826e571df2825a1d53aa302bae10ef5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67f8e6ea4012bac4aede821177111c1fa830948e28bc053c7615cbc7e53890465fdd5eb501ff676962654e35074234e52a829db194c1902c6540364f9ca3241df7010fa5d476f20af940935b786001a9a3ad00382cc8381e37c180254f5fa823e8e1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbac49181dde84de87e8789320ab0a83b0adf5a6dc8eeb420bf5a0b8ab9650081769d51a844ee6e7438028d7bc47428ce409d7a093e9c2efa216ddc6d6f096a351a67799e7330a89619b74d1f928f293c5c361e01553b00cfaae6ada8dd1713be0660;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59125ee666af8c78d199080e72c6673b289f25753f5673648d28719219082f5f231ba1c852cebe88085013886168d2835ea0a7679d42ddd30a656ac04212f9070d74c732250eefca19ec94c6782d8f050e5dcf86225b6348d679205eec5ea6b8a0b3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h912786737180addfd8a430631415f97986adc00da78097bbd455b9e8307bfa65cd0688613b67592b332a8015b1f6f8b78685fa5beaad8709bc98cda0e01bc2b58b47f1e904fcdbfb2d8750cce024f786e83c85fabb0b24c83b7821469fd3e0c6a13a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a7dcf6f1a8202c7d6ae7d76d5c9076f9a7efb3c273bcf6c98e80d06e9d3f125294797aceaa87b620486d8fe57676e2c9715b40bca3966d82d23b6a0b86fc8a25759d321ee33843c7e24cf0b20f5bf83eb4c3d4e84dd435518094ccd29d72afe5ab2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2e4a28d8736ab2be688d6a322351ecd312c990868303b4021a792423366ea9651f6b14b38f12257f61e8afebed3a1f71ca528d97dd217d6faa95890b0f98d56e78ad196501fad1fb6eb896ca799a7901a2de00faf934ece847eac0d3184cc0a38e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb95481afca91954b4b2215bd7936c8bc4a80871d5cbfb2bae5f494d17845f5a1e397afe4250ee667f2b4936f3f22bc8c1fff95536c6e18a47917aeb11eb58e8a3841f04c6b312aefafd903781dd76e09aa2e246e015c96ac1fa2a2e5d999ccf55b8c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff4c669aac432c71f5d7a4e67ff032e14bffcb03e353c1261c6583008b566bfbb5fe226bfc5d7f0838d842289d848bbb81bbfa4efcfff3baad7e3bd6876e11a7e83fe985489c4b0e3ec78ac258bbc01256a8a5005039b7618cae26bceaedeca70f21;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h621476fb5ba38fbaefb6f3be4582b933f249208c6d6c9debfbdb8bc30512c9fa942a7d665b49a84df27121199ecc40cbfa5410db7f877411efecabe1131b40a314ff33fe920ff5144b1a55bcdd042297a46e5b48cfc1f1e8112ae4b33ed6144bd20;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bb15c0c6e53202973174bc2c6a56daebd1e63ee37cb853e9b12bb02446c64c200aa3d5d5185d22ccc5a95d7225a24d44578098fc36020ef2390180d518bb1038b394b2aa82fd5309f958a0ea0c106e7a6aa0f36ea0aa907cf17df0c0240cb591a8b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6084e8dc18b064a94fc171a38b2aaa1faf95bb6b6b9314c0a3b7166c86fa8507822a02bd0acb2cd4cef5e42dd589eb79cd141033ba927df9833832fe332926828f898aa7f7c626a610180e0b1a9d4d3fc28fb19c880200b53fd3591be86f537a794;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc28023d51a50d025dff868b6f46c5785dd7a9860fd556c64884e69d31e032f4e31087169e015565a373dfe0343e627ce4b667c3a9149f31b03c26a321195467a04e94dc75364a817f0df476d50abecce733adb8033b62bc4bf1ad743def29853083d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8087238d7fe560eaee611af1cac10df4c1d087f4e138935771f9cd7757e44ffeeb2038f9c52a9b346f727c3521f8b1c72a531aa20400b43659650164971a5d117b69b343ec67e12bb7267246eca4e59edf30a4681b33597130b763c006e9dfbb9092;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e2cd49797e8acb346b38532610d5cd1061e0a5a1e69aa7a83ebfab1b5059913964d6bb8111c6fa4a024ff3d26b585c2f84cc571b2e92e63496c7346ec59e9d736a42e39f335ccee09b2d03d03a394fa2e972621113c5534d20063f5239e1666017f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8210b308b478136f0bebd6a044652ad83cc2b9065001fe0734dde4aa292bf4fae007c187e3291b75e83d67b610f2818f6f63236bcc2974c62d5b3fc9363d13f6019ba7b7c79550f9cb3acf373e720984c8bb2cfe6c442170a6026bee800e6c85f7cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heccb6d92f6d7605455b53c56f9fdc2575cabdefb85b8d652ab857391316d87cc374612522bd4e583a4b532a6477ab113ff1e998627aa2f4c50d86dc0f1163e389b6babe947f7f378e7e0f8444093cea104109fd3a7a01a2adb1d52d34aed0dd69c10;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8c537d30080e01c8f1ccad07e7de043c945567f3160f78b5e12a5c7b0937f6acf8e3e8e692de355faac5cb0f8d380ae6b228ba2c90f337f45f9dfe3d6f33c6d87c608b2d92f65e606396f2ea741e03a9647d9d43e2b64a516c1abeb6c5b4273080f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f5d5c936bcb66ca1fa3620c157f9752f160a9b34d0a34e54d4bd98bfc2d8e661df1ea6ae82df8b6625ab2828c7593663cd2d0c51282872718de71f620e338b0bf1c47071668c1c0cdb3e57946839017863ec687905958ad847dccc347280cefd000;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf86b34531cd2fec8a0418b9d54917533b7a5e23c740a58192d86f4fa1f11dec597701251bf4de57f58a0c2a9943a3028aa259a33c83fa6146a885bca45d4a5d6451469be33ee9e0c26230ce20d5ad7e49a44177c021fbad29614036e90c4707d5e65;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd0e6ddf3a3ea015a2acf42b3d45ca3de87f898c92e051fde693e0ec2cd02586ee4496aa2ca5092745cc57439b23a276a985e7a2e7ad757c7009345cf4b3f9f0b5508921351824db74b307ced2d3101df9185daf5f149f294aa76546ab54133950c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h596041c344664b80cbb938e501204d2e35e977b7e60ee333b32f3a07db5e7cf7d1feaf58ce5f76cfb76f4be85dc57b9f007e1d077f6408ea9d428b8aa8b627e7216cbd8f6c09e71b3ea08a15e301f6fe60105b78fdfcd2273ea52b18b7b744495854;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h233d446e17a6603d1b8d43f652e3493a9f2361091d88a972fde7b705eab098728fa0cc36f80bdafc3c1aec9fb544640a72135f25e39b3bd238c04620b701749d8214e6191056c29e6147c0bf1c0f349bf8a8c4aadfa0ec484255aea8d0cf13ed77;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2272bdc0f760b9efe141db3f877b5638643ac5c5f29572f5d86b57079688b40c7a89087979863b4c4a0922f5379c7d8c136514283d2225cfec35a0e0e84a02ae2214c6694f15ae122ade2d2c2f218bb13d30a7e7bf2c5ce1474265861b15664ad95a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h564c88574f4d0f086c095f5f6624aece3219cef2ac852521f72b1eab977c21dc1a5ea43be3c4082e055546f05a9e400f4dcfc03e13f6d041c51bf5cec9fef3c4b3d3b72ac052db1c7c3d9b2d15bcbebe85ad683545154fced8f8ad8bf93b292fdb0f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h233fdfa83beafec4cc5715c2f38a92c6a2f140801b2598f29cd5c6f9b5253adf934a90c783497ad126dcc9d8256c733912a2d5062a8c0d0ae3a7d1c43145d80282d8ae8d98b4299d7131cbeb16be493a52eb7d74b8fb593f146bf335b11ec24f171d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha071c8dfadc5d71ea3cc274518630a963b853ab77137ba986aeb8602f013bfc884aacf0c3fc77e25dd352b194cc319b673f439222cf5f1fd153511b18f13152fce1d8d72ce7ba77948a97b1a4e261124e36f00f37544a4450c7d74628895c9cfba5f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58dd7556c93246cf19ddaac43b6d6470547d6c865ef14b45e6c292db60de7aa99e4029d1c84b68a4d1b7c1872cf03263e5d068b80f49d0c280ab58c1696929dbffb534a964fead394812ef81cdd1c85d6a16fa50e3c74825457a4354e708f31b99c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55b88f5abc1ea89215d587c59c82108f7433e778e1dd519a7b31e88363f5ac1fdeb41b36d7c4f583938c569f8e5b30817edbbb22be5ede944c07893381becf8dbcb6c1246c496f6eeaa984101f11a40119376ba325f500b4b1271025a8dae01cb2bc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heff7d236fc139c0244a25f539df704e5413ded9603377f065ce875f72465a3ade7bf9cac80e542ce63610b849514dae1364d1f449b5331f90a4f0c49b07e00cd1d27d30f43eed69b71da5050fef45f147c67f769cb6edc88bb1c565150e73b51b3fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf31b3b58eac59f3e66573efca2acf082be4939110fdfdce174638f09ee7d8a785e111d76bb2011a81b90e5e3f13ed117a5ce7bff87bacd2ab6a531eb1e6efa2a7e9dc5a9d76d394e9abbe9f097a32f09a25d03de541bce35e205c90fd015c9bcf63c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e72959a6e443da17591a257c9e3ce3e4b5b7c6265a135b11efbdff8df7669efea31134071e896b54be7448f54fdb2fe30393ff84c2c714f2caee0e99e4e98c27df93c7f26be92f3ba8205dd3c1d89764ab12e3e8ca3a0aadb77ef8ed4528ae97c5b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h857a307aafe45ca1e4ab9e5f5a39d683cb9a684631e01d20fa4c78b38c61461ac59f923844fdfe081cf3070133141d0c1cc950176cc6c57de06796682bb8539ffd334f84d830001fd8c3cc3146c9ab423843de1b5bf31dc48b6b554f6c7635c842b6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdce95fd22227174ca5a823e0f67058c60c0717e693d9b989821574a0b8fe19672207fcb9ac49869fba4337907080834931622c2413b90d31b3618ee8acdf1d0614410bfd9a548a895b41eeba821280c206377d1725f681b4d6828f71b11981374027;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d1d931308a47596eedba42c4e9c8e15dd208bb97cd62686a955f1cec0a1dd835526b1a2d23ed6c75e152b3cb4e4cf1c474a0a5b1998a151cc6f9c3739868cc25223585a74e19174af8f9f3dcb6404b63663feddbcb12208a1649d3ed6464f61ca37;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4df16911352a13f2709d58a38c2acec0279071ce3a71423cb61ea2cecc3200766496ddc2cafe88e96635aa5054eb7adbda48ec9dcb76807fb2ae3e40f1864017e4b7106b9c1e5a3f5439ae0db01bcaf212cc9c13fd646f477b78df74cbeb53d68e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbebeca17b74a6960b29b45783532897b338fa89c8ac8f41934b114fa5eb79c46f2490d26afcfb70fa24230530ea940464d9806883ac03e1c4b1e8ce12b9b94f23e66f20ad3e74b9bacd0787b03d5229060a702ef9ebdbd60da05df6a735fcf1d936;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66728fe131774805ce602467c1c24f933b8fba3ec0ecabcaaf9b0f026d31f9dde68d0f965b9fc92988ded88fe5fe16b660158302997423aa633782e3e224da13fdaa068e9964b3b86233100cdba29600dc7c4669996e3fd3807f9ec532a2bb52ae6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9014406c8fbf8007c1ffdb45297b859616c735354c71a502f7c4f8b9cf7939e15677204c6e71ea88b96ab002b162a899bfe9b685564ba728708bf81d43281d28e30ad4c8f2b9903274e48f51649d69409a770ce1257e433b778b30f645bfed5b87fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b06a1a6219aae13d20ce74931214455a72dd446326d75d26ea265fa87997b3875b37087c5873c8857aa68d74934495f712b998d7838d311c315d70d9602fe1b79d7c449514d35d08669dde4971ed181cc894ba75ce6883716a0f8e7ab3aefc50a7a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h675f4f97d80d1113e77ce36fea99a99b369c542af63f516a8bac85e3ea80f8c2da71902a79a07639b4248731d9ccd1431c0f9a1e58b2a363987f11d0e9954731350b738d4ba959a550ddf20504654634013581ca425f5b6f70605982a6897f8566e5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8af9d3cbd5af8d26292b11579387849d51de36b954a079206a2f8203d6020cd98745ad1313099d17c34b6fbb54de55e19e6bd000363ace65c934f00a6e820780cc12d20982619b80895c71c3527aa88d4913f909ef19ca23cd81ecf443ca6793072;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3f6a06fb760e2a288fb8ad44ef4e10a5fc776eaeef332c97269b0c103ea21b4616e7d75af10a6a72763d34a9688c0a7d1d95537114122dc81b284a69f4a2c272a3491276c91a00029cd3baacc4d4bb7a8ca70dfbe17068965cf3fb92ec5b17277f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f856b6ff51dca4e7e751d794c28fcfdabaf900f16331aa551738c5920aea2eb1f49db1ae2ee2d19a51abfdbecf8dac04bbbb009c9318453f3cf2aeded504c81b9684192af06d0ca66ec6ab2422c9c88b0e3e2d659075ae3c3ca7696472655a53b4b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f70db01f64888f8f44c09a510f4002dfb003d968d8a8213a7dfee1275b5d26ee1f9e975ec6a3dc3ec683b29bb419bb08dfe820eb33b281bd804f49eac15c6329c0afc7238f5f6b940bc7fbb15ae9e11a720d79c0dc68b157c193778dfa22e4bfc18;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e5fd47f56d127eb9798b54dc408477e5f295149797985510d66fa674f2cc7db53f8adb27af7091b8c6f13047d8324c58da3bc918d4abeab85147333858ff2fb95e099352c375d67561e74f35037e0a59bd3569bf0cc3dcb92a79bcba7a6f1b12d30;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc72ea483654ea679e66ab465c0c1c2f1e3192583ff8b5512f8a3f0fdaf389014ae3c39f55deaf61512590f0dbc293812d1b56c0801bb6e702c284d633ca17738f6226dd9ab582aee998141df4d9f276e3db1679149abb56c9ada80e6fc990da7439;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefeb398b808ee2a870b8465e13f00885150235832d6389d84cc7ab3b59b40760399984a43beddda5ac1d69f77905f46c56b9055b344500d85029ffb38846e2c7822aeb5970d99985c76b1913e71453925c6197117564cbf75d97e4b9862faf11f5e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1af58c592dfe29660184244042640a44bb52a317af31ee57b787e724b304bd1d5323d023c4f2e71f3149ea2d10145782eae1b2269901e0fc526a9178aa17d04fe43b4235de0548ac3d39a094edb8e529925b53d636840985c7170a3a44fefeb4212b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd1fbc75f0c16244428159ef5b9a75dfce82447c39fc953d8f6ff13dd648b1a84c799602d4dcea422e7f6d339f5c6068c479feaf55b7124266611ef7545121b2e851e983ec51542bed7617c61ba6c3c0b52625ee44ddd0f232b17b61d0c5e515916e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54d8c27d3d35594e4e51ba676f0705af644e61f1a77d8ab4600b3af37e4ce306608bcf2942d0a57b0486865369442071dd79864ee1292bc5fb4bd80d102ebef15eeb2e872baabe190e010cb7fb7ac0ccfb6d842c5ebb598a02757241ece75c0e40e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b503ac6a1b1c906c30a87083cdd8e8153ca84410b1c3391da45d71279b0ede310220a5230ed009ea434bf298cb56ae8e91963de999d3242a296a53ff268dda9208de8e27e324d6dfd67695405cce6ed9b1d2177508cd0e84fa8f29729428c64dc0d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6f2c0ce478a40903d2af1b8498af866a323a0bbda649ecff8766b1ce397dc54bb4edfe7988eadd67382400c13199b31103c3bcf2e2a4199af11fd25311624cd61260210fe6981bc65b4b968fd5498716a1fba159a0494daa13087b5b0a5448c459f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11a83bfcb6df1fe92f7d840313a8171321855cf56564c35e91c30de65bf76706b836ebc5bfb958495a571cb88e13e4e62ac7664b2c6c237aab38c0249d9402a14dbc5f2a4766f8476361194ca3105da6b0efc35d075140ea15c7ba96a52731ea5225;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fbc1d124221136d01e1cc02bbf5a1ca865f7829b24f89729c13d65af914547955d052e4ba75d8c9ab2debcbfb453b00acb163dda0c278fff78b7f29ac0ac918f7f7ce3d9586b867bd8fa3813da9cac91b2f7667126c7b611999b28329d1f065149d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha43758a72d4199eca0284d7c1a33bfa2c8be69b226a57d4a2bb593c1e8f9c7e8b5e5e41f3bfc01590c7c95134fea51afff71b51bd113821e9e7501ba4edbb52fe125280fc28a02e321a8f2bc34a0bbffaa3f2f28fc55ba6b2cfb091b6d655357ec60;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfedc0d28f7e4cd6c01fffc650d3416d00dc0ea4b96e61f9b440fa1968c0e7638dfe07c153cccc99a615888ea6eee45ae4148f86a892df1f3b2a09f3911940036bd09ef0b54ad51e3d954055ef922d3a8618f67919ba0fa1d120f9b1dea438bac1641;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he39fba1239574be14a17e63d64d31ba99bb7d9f207d9361c32565e2da2948b56fa3b52f501cdc3da2e737b463cacafa75b27650eb16fab95b460e333b66f8c9735d643fc5975de23d383415fe75712326867e9398904c30dfa978d7e45ed7c7c5dca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc86db9200236e1f4e71d018d26c47b3af8c0a8650affc64ab9411622d69d26f96cff12ed4a6bd40ce129c0cc31ce79b937a8020187face5cd21d6e6b582ec34ff2c7e2abd5902a7364a500ca396a7656d41234f582a44067e09cc44d5ea41a6947a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d044b9edc5a10ed68924e56f2037c49a7c27855de6f5437180770d12c402e44fd21730ec385928ab8ae2f845b4ad0a43927ad1a5828ef5fd942e0494b4239fc383c00a58f149af9f57f4d213afa0f74034402f3d501834b2b1ecaa4c63812eb142b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd81333b33d8bab7edd120eda5db736d868e8252dc5992e8be9eee1cf2da2e40f8547c9210617bc9f41bedab67de08edc84161cfd7b93fcd1fd92208cedc5c97d77cefb18fdd081c7632bb5ea7f54d0212a6e6647c1ff788c2c6e955e2a3459a71845;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcebf05ece8913d6043eccd88fbceeae22a34ba77e397c40bc24a69f830cca465a32086db9091985e86103ad567995c01429152a83f0335573b67385447b3a959bae4c67c07ff21bb35db2a53982e10c3209c51b43fd754f0be1372c924f895314847;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h257086830368c024358b1d57fb6bb91f6cac527e2b18b26f652fedd9e932db40f16463a11ff1cf55604b581af70f9f18e8162790872777dc35f83a60aee18994f3ad3e13626b53e04dabafe1fc477e9dbc0b0a77c30128caad5a0d100b2ec81673ea;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h283c8736f9b8d1b4bdb23f03c48608e63af2666942bfef792da77cf541b1fcc36f04e67077465c275e417479e59a5fa90a00603f6ce484f5eee791a510dbb3dd04c15f3f1586c63f7f2aef6956a6ce66af415f8685238c6a0d39906e98acf3ad27d8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1ee42705dc28453e5a332834ed983c98fc4a84c8f90ac0fcbf9bd9faf4e035ce5999dcb88b3cdc11b25062ed02d939029d95d828220bf22c343cc307b26dac89fadc715be5f2dc55638c52db1443b910b141c747ffbb4742ed4938e99cc36f93e4b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d14f71aadf904165efc01216dc114f85ca916bceeb51f7e87472d085e7decab5100a873d7fe7f17a40bb4c65d8f15f3260700aa3b1d1d2573b25db9d5fb6e1a4ad0ae1a1fb32ad2f943aff0a81aa08089c7c3d4bdeae210d604210f4103400a863c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h213aaaaf206bc4382fd5c8e423491db4ab2206714ecba768264b945cdf1615c97df6582ff9b01d7822ad5dcb932a8561cadcc9fe0dabda9b7ec7144504cd8ba8ade493da97c32e42e99da85e03351ef4d4c1cc296f055420c5dd63b8b78bf78411f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3e74a894055a2a732ff9123f9f346f63796dad6d86feea472a784faa4de7a52ae6898d5610d79c47b2c6a15afcad5ed9ebef6e8cf2bf85dc3b9dff703efcac65b33a3b9ca3f9a4170831cc85b870620803d28f922ba9ee7ba31e89b0df4655d22a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e562f27acce3a161b4c8f09603cc48205e18449168be135b4eea0bca2b0790c417e838f57d9a03911f381c443477f603b47ccb7d180a100df46f5c1b7949e2bc84d12d463ae149256011707d8d329e5ed1ca2b4a572ddd381b21391191229281984;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7962d1b559821e06800cda916c08724bf09113fc58d2bf9feef087d1cf51e19c547917e53d6b5cf0531874609fc67e23900244d611a6a691a77cd46851f28241c05b258b11e7b1cda5553887762cc8a0adeff08b9297e606c20faadc0009f456f0e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcdb09ef43c950517ac8cc29677f10a0e2268afa96244b22e8b3b4b8d63d5116a62b50b2814ca6929640af2ece72e52208bbd1c8268d2b60fc729a8959b9f8fdf034c74662fa01fe7a8bc2025479377c48c46175e609e37c29a0f62ac88bfbc4a8081;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90df98d2ace1948b201543765cb2a8dbb15bdf897e2365ee4d8e32a24e091da35012f7240a78f46fd95ec9915006d6002c9ab4b76edadfda8db70a1398a46fe8ca628ab7bc9bd9e826bb653ca5e033b3276e3f4e531a49afc28304faa10c208f240f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c8b80eca6df501c690af78eb6b72e7b76c495cdd0f3b320e44d18caf8a7ceb81734333b723d767e622941140b1f35c170cf9b125bda9dd9b72c434b9eaaeb960be1f0646db8ac494549514afd1e873c0e7e6d9fd1dff8b9c12e52c473e52cd82f82;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4fda6379f47e42d09e137ef30170e13e079b7fe9cc18ddccdb8f2f8550ca160d08ecdd37c7d0bad152b58e4674bc815440b232157654d6ad12a7eaa037407caf1bded30eb9fa7e6cfd6f82b58bd778e402b5ac8c5d6dd4f76e053cf0889eafc18fa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf85c3c226d604ba7d0eb035eb645bec729fdcd955a8b3888ef750e3a9a41c4e070a162d45129c6a2a7b073e5bfd9f35b976be7566e99801c98e86799b91437ca1acf50cbaf24f116280abf3d5164545635976bade8f0ff1fde9c6b27de09c643656c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa771065f299ede54003a8a6093e1283277bdce380c69ab26d5a4efbf8c847b7df893b8fa755f4c0ea2080f57eb5d019c02d60aa063cd1ecb2e3bc761736ecc021eebbfc4068bb2f6586baae8e2079d02b1d86a4b05b7dad3d85d479e3f43d1578c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2119a168e6ccb344e987fc7cb639b3cbd7bfa2553a496048c30b0b6db3378128a13547868a3382ce399027f99ae8d6f4989e023f667bc8292d7c33014a24b8552b090e8ff95ce68bfbcaee3401d9a784b55c31c9d4957b516b2cb157d187d71b4c67;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h979c3247a1fa94ae37d42020fc6075767c2491edd7cbc0b99bd3174fd9e09318793a3b4ee671e136bcce543c251f57742342f0e082cd5d5dd044a3e24c95686111f43d19bff60a453d21522876b7e5a2b482c55637af1c5331430d2a2e6b6d7700a6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d52ac5d07d17aba9422327ff07e8f2cf1358818319ff7d91055cc74b3f8b85fc15afe7e723cc5de6a52e3856596df5420e1c4cfe84251a2257cc77dd6e924f896b4f8a8e63cfef422f25e8daec887127019c762b245a55253916382a6f15bd90dad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h850cde2af757e54ceecbe20ffba071f7836788624bdd0602a8a398ff0bbde800b050993723592f7e6883ce509422346d3cc852c5ffcbcf9cae633dd66706d50e56e49aabc6620dd9ee7e3a621625cb3dea261c1754c1dfe29e2fdb08b7173080b21b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf3fa2ad6c6b9a39c490af3d276d5090098f08e82549a22e251296071bd4178da284a6008d76e2698a2ae3baf414581c34b10c07221a30aa6237294ceeabda14cc6d1490ab501f859b11bc2049d4e133449eff3d2c729c5ef5d9b994b9658d83718a0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87cb70b077aef0724cdda5bb6b983647ec9a9b825db25561f5983de7b542d713ce943818b400e3f962e0028931ce31b7d0790599ee338d84bb397d29198e624362d110082e0f637488ac88eaed0fa11290d562156789b738a12ebf26867444a5e294;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd40a662cf626d5ff8c35c92ba52f6258c848f6362b8ee60fc313451b2b69db105266dad5430f1ada7e1ff926e052361703fff0df1d2c58f370bc214b8c77b0f6713742fb3d700795d2f2354d34eeb1a556f184e1784e7e7b6fa851f55f2a7af48da;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b3bf801f8185d431e76603cd94fca8cb27f4975d090cd9460fdc5ec1b1c9737f01d125b3a0aa761325f7b811573036ec12235461a5d48f7fe04435d854a8d182eadf80c7691010d9ca1c8297231de05e2e486dd322e0bff7453fed3acb97337867;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94b42e26c8323c58c146b44dd09847ba4e0a95fda89355d3bb2dbbe017c1c5a9872ff840ccab1315ec935f220d3446602e6ad6e7be0249bb7b4163f62b95363b4c5c6ee3c8aeae63d4db0be9bea86d1bf4ee7d79795cf10f5c6712cf91eb7973b3c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h940ec8241b50cab9aa10dcb7a1acb7bbf1ed56818f30d1181e809f3f96d29e14662a75a7c58e09b09e1ea4208c8b73f387d5fb1b006308a6cd901ebe27c951dc0a5e667b446bc68a1ebfe889a8363b5bd98f377a24a48f9121b35777cfa55a8529e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8224193b8be6460b6a8e1df2c4d1b624877a1111e4cb50ae55d80a5989e9de0146ccf9ec024a6e2bec441e0448e225116006f2855b209fbbe892e791d4c947a181776b474868549f958328f432924634a702b5a4612a486061ba830580d8cc4f3ab7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd21b8546005da0082e2efd175cfa8c775194beb5ca215a8d673f438f1c4c92af3ec9905a3680d0da99d852dba003b439b6c9047a4ac1f217df599dd35ae994c781494419ab5680f53c60ba38fc22b6c9dfcf81d9d26cb366c62944e736ec1b24fa2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b9a226dab0621c68b0356618613a77c20076d8887fd2b42f5e0e489344e1b046a0550d8e6cea928ebe7b555d0366b9c9de282fc5a5d68676c1f58a250d0a44b37cba93325e52b1796808b010f60047e47a0e6dd4c4a6cc2f09b8075f85319c1d653;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6171fbf8ca37511900ba38205b94ec3f557d3842e80f8813ced08050eeff4f530611c4f23e94bd5c89f9e114aba63c28e0d09d734c820f8c8870968549cdb2b338284cfd857c544ca3743d8dc7193c9aed6c856fc71fd10d5289a029655e2a3e8d5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8976617aeddfaa26d2785bb60be80b4ebd61a2e1694a4b9adacb8035098a90eee4a20aa0592f4048d53180381fe286d3f63377977b51c271ebc6b7e98e86a6052c9d1f747f57fd3250bb2fb374f6985ccd014e08fc59375796aae3fc841b71b997d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37cd1271905948e613a1aa7d5d9218e6a5a88004a66dd9d81e95e4fbb961c2be1be43dabe1ff34678c6ded98658e56996bc23c97bb4aa83e5188d3623d52e35bbf0045ca66e6d28490e989ab5bdf629d92310a877fdbf61da27489b8dda882a0cf0d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e16e1838639ce45241b3796a52e3d9517f474e45ba20f27d3161b77ff8ab5b04cfc847ce13378b658d3eaaa03f5f3a51ec6054bd36fa0548a98ddf10f9e044757cc87b07de96494a59084bd42c22ad9c6a2a1272267910809fa3b997c40a3bbeccd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c291b46de05d9f523708b08cb73afe8db065ef946ca1611e24d25529e0ec5d3cc88294fd438ee2538ed69eaa71265dade9793d75c56278e0e5a2127aeddb8c29db7abbbdafe43002e6c529f747780147d2a5febceaa09d2f32ac5add2bb70625323;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81de25490e19f8b8e15083545db2c97e5924c8f9e6c9a36b44dee4d26ad36f1aa924991cec9730bd49a5bf7ff29d270909b6315c94c67c50f7ec3d846653f6f382f740e30fb1a7b2214034b435614d988a85b0d44e8e63fc73daa0b3571eaaa7d20d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha450266a920de1e43aeeb21925e0440d55162a4e2db61e040a9e13cae927860199a3e34f6394f83d9d85ced332e4add824be8e886bf04484e24fac18b44b4ad335359342c6d571f818820ea7ebe98ead19829b657d72c41b5ff88ebb73d56fe7fd34;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38b1c62ddaf7d30f33a24c5214f3af7c18e7095974f653fd36c20ff37e73b898de1046f35a8579a0cae5cfbb53981a16fff31139ce24d68297df374262b57fc3af8c56459e8f78eeeb9a7169971025ca513afdb3fdf208740891c61977b1e8e5eaf1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6bec894e25301f22744e6e486c72d93505fb0b57f6cafc1343e06e593a2c155be4f2906d88a038acb483f8d749e530a4f90cf613b09dac3f8b5c903c0d2f64732287252afca81f23625b7d4806cbf9966cd77567d02df03fb8278690462ee5f73cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a3c9dce7fc469ac5af7466332f874c5868c2891b7a5a36a8243d570293f582c84a1689af7f4469513ef6db03ac956441f4f21f1b34b0a5e0b4e91ee6c9f60aa7d2970cee8bea30f4cf954b654627a5a8376602481a588c42fe3054306008a3c3037;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1d4570c88892e85ced3dd867eb1d39fbabb11ad09e1843677a7db8729dfbe842a1acf28720e8991e37093917aaf452a25044702bb1bdd920c38d353c9d9d27762885f742688dde4c0f2711172fc5146538e7c13ee8ebdfa75c4c99c3a65ea353866;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d4bbe91e6137b231120f07a3833336443779ef394fdf7f0624b0e2cebe07b5265db7a8549141713d6169ea51066935d3756c7fc13d730e78c662173f20e20679cbb96fac51b74dfecb4b846e3282438471bd31f3fe08d20e7d66c7dc104a64ea4d1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h906ea66b5b0356e23fb153b223a34106851bb8a4314a73bfd323e72b47839cc1639bd0c2ebb15f633d001dea63ed7e1a484c3e8a4e91fb380dc5669cd1eec5197db269b48bc4e3dfb21b996f41778ead0d1430ae2d9fb02a30d03be767f82f20d200;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a927d81facfcbd86ba235758c38beeb1cf2eac2ea63db50a971e7e69a27204f817fe82964306f310f55c2d49e19e9e837cad8112676ea7b71a0a31c1a4f8b6ba8b8e79d3d5e021e3e23cc28a74d070fdf9124c4623d4eb89bc31ec0b0aaf9d714cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha81dca86b509da53bb63cb5269bb1e2076d08c40e513c230c5862cf439db51fece7c08e701d302fb88d7b157b8d0bd04cce124d0887733d3e2def5a8b70a92d2d498c8da0bf318c018ead786ba0b2ef2f5f7232beab1defce4f5396d9f3842d6a46d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a1e4e8c119f50bcf55bbec0f15145091feb3152bf77f82f19003ac24c61ec90b1c75485fe7929f051fa8b816def93806c9918239e9909d2c44162b9e16044bde02477cad233a16ff5cfffccf32021daa7d11947a0aa659598941ac270cc77896cff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1be146e3fbf0774a0af3e2483dae75733a928f036de87ac3d0ea70b6fda25444a87bf8a2425225fa4b1832d92741fdaa19e7b2a4d508c4125b5e03259d5d9dd122d525c72702661b022c9ce9f765b85859aba7cfa01f31e9e9baf923ae41616810a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf88c978027d528d85c9c192d1ee541c4dd30b7ba270cea8d3fb98fe622469d216f3ee04ecec39fb1ed422b7e9069e65c118c9261cf83d627937f4400837111e72ed817095d4329615b583cb2bb46712f5935a92994931b9d64a18a2139ed19585097;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5b03c1d2c5d0b663481150e852cd031bfab855c266a52ff1d4167cf8ec01459d8ba9edeb96e1d8db047a020edbfb991ae1d5d9431ed898e7e87714c46473660b00416cda27fdb16bff7675f3ad71482dde1c21b666cc312bbc69a34f4d76f3794d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1eb6f1268ae17611eff75c6f30f127cc4060ca49fffa04f47d04966bd6f3b83e00b07b5d327e2d058f375998538c24e3c2ab91294ed877109c9933564cac0fb02aee3da1691e384389c46359fffe6b94109a6780bed8d9b0635b98989ff262b72ee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34cf4429b636e6a079e4e946771c5cbd61faf7e8dcffe389115b6a449c406457191984d7eb63716aa51c78e70721abfe66a43f624a7edfd8fa1aebbf40e0fecc92b7ec45f28c6277c25eff872c08cf3fd27b996d04ea48e3441371685ca00cfe7f86;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16af190446b77aefb4c3951ca0c3a557377cb4d33a58404fbdf516cd02e67472f50c21132c86ca0d043d259f21c6516778c894b4141f87f26224a126fd5ec860e4a8cec09bb82d48861a6624a62d69aed4a7eb2b80c30dd2260eb138243ce2015837;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h460c3357cc1f38a7243162492febcb0e5b74952bf252c567232021aab46d01b387ac6c80a8f00bb2be97c8cf27de9a4efa1587a230670560e15908132b1f8b2b84d62febe22c6fd89c71e18c945e1887e2508e6d2e1669a761e4ef294592087ef52a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3633849510f35383b72521783f3b681061ddc66a40a82302aa86c9b7aea9cc8e375b95be3fd8ef9e89eaf95186c5ae131d3a989623ea669acad4c214f803bfe363bc97728f357dc0c0856119402aabee3a60012e2985d1308c12ffcd42dcec1ec83d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h405fb63b52c3beaad381b7a247bb72ee6468758fab3eab061909782de40f8ccd8185cd9eef451323771c1d7a0e2cbb731dd4becd37ab975d2c0df4c4d347b3dc1fd44e10ec915bdac4cf8bcb8c1982f5fe045e0a4296ca94cf2194a78a825ef6ae6c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h461db2c26c3c586080a6f127f768655ac5f4a073c99c5c838f27a17717f712ecc02a20f6e5348a845ed7fd19ce3d159968194e49bd9fce3acb43dabb3ff58ec3c806f792c65f2b7533ac28d8f4772054ce83351780d87de49552b731bb937a2f336d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf567423cc4775ad379e6edf8fbe0ede5c2c7816aba72f932bede910aa5dd6851f25e7592e7c42f2ff30c2ee94c7534d2517d634e3b4e200e40a1b95d82d84af698d2514ccf813f3d6973c704bd3f87b8c958d96df28f20d697351d1c62a47a2c2195;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13df0bd37bcabf45c1105ed6d181633693d244e0706c16f37b1ad75d23a01792cd1536e7958a6e2030c408eb2378062a02e1abed6646d53f0c7e6046aea0fce269efdc55e566d46cc5d354ba0e87bf4745200f3a39af9a38f2a798c18f54cfa2a0c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h65a187f30f0b206ecb69701354768db4b088f95358b4c8f35ad1c0aacd8d44d256c6acb873a381a8da91678cc57d07eaf937b2728eee062c5313248157bec6d6834e4590447a4d5fa352ab5d6bb8cdb983a4cfbaa4fa9936c99ab4d7d309e23dec5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63c309bcf6e72dc43c7391bccc589fd0fd27a3bcf4b04ff41086251d2f36910f460bce92655f9982433da259ea3fa194387cd6af63bd0c992467fc2c12a3ed078fe65de7f67cf70c26285eef6311c85c73bf2e88f24ef6e7b12e42be9f4e1cab7371;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha627facd878cf7b63d79ffd8e22b6a9a66de402821a4498b2ca21b1058b0e619e09b1d2a5a1cd232f6cb08495dd46d0ead1d48e6bbb0dc89ced2c68515e03fab29f70c132572d41ec98d3b7026dc3db3b305930415579fb75c59c061c09df387f3dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fec1f47dafb914a6154a2d7240f62b65f936125d9c4a0e8e620f7b3c49b25a5d9483f7fb2b563426e602a6ca42c8fbe66538c75084a0a7c2cb2a9df8275f99c75ccb038a8e98464b6bf722db145dddd6caa794feaecffdb509c96c5799722040fb9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf091dd2372bf17847371963cacf2922a516a18d0d412e3631312ee027715cfb7ed3fd87f3487f16f3d8d4acb68a4e6aebf01acfc76382efad3a0b805f707ca2c49499bba8d3ef4d0ee92709ff2b5374b18fc2e51aad803823042428deb945bd47e9b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45e79d9f834b74fa43f0f539aea9ec2c808f945b46f3a575f704e6cbcaea094eb36451ff681d7b8637f4b2155ad597b47b10366957c4aecea833d4856ea84f615af65f3327270fb2e6e49cf62b20e951b15551f23161959d9594cce363867d3b271a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h86e0588fbb7339651614e55d1491ff38bfb27d1b9837a973163b4bfb0c13a9bb0f20abad545ff221c0f0e377ce11a200030ba21171fd4d7ba44db579b875ac170e25e0fc93b53cace309fe21b81ba52345627bdb2d33301f054062f4ef1639343d7c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd855be36def4d636d284d6f9e4982dca12ecb3bde3359dc62114e0331be17feef28f89a7aaa79657303e0fc6a680eb6a80fe34f202fdf3a4b03b1004669943a4009b98ba47c1949d7c57b951ffaed43b62a14adbed6d6e9648afb0f1ad515a4178ad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42ff9d16a2e4c1f8a4a0a20b4544a066573c90d4d4154160bff98b51e122a12b23d394c4089ce27daa33f2fd39a53db76f0a587eb4972872b37145eda4a7b9059aaa40fd7a95776764e0500c6b558c0301fbe6ef983b514c03f1bc2ef966bef852ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1789d17a4f3d4daf43b766695310dbb6eb20b7623a158124d86ce4d67cd5c165881c6b05a3ac57993ea49c5b9a6ee06bed164f9995188fac4e954a6332084b5f28f206d2f29b42fa777f0966bbea988cb77d0fe65f5c5886e05ed61929b4a72d345;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he79f997c0e60989bacd7906d52260320a245b23196596289d2056ddc4e0879624a14522b17f1fa7d004741846c1c53b376dfbf1d9aaa770e679746d42d67763e7bc42532ccb15f77d1e9f5bf3fd8315f6f25cd395dc3ab55f76920ea85e8639f029f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd15624182a0f22c5c198cb5e16eec2db353bf9222d3c21da6607bc25bf39237a928ac7e2f19ea48522d47f2a440fdd3bb0e47f17843d1ae29946b82f6583f41be945f2a35d2604fe71f945acd9bc60dc943348f7554b3f6c0204e065252f6955e3db;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc79d81e9fe0aa2a03431b8a7186ada7a163936637fa89fa0837495433aae093c0f3d578bbc3a9b9bca529796af5b289ac7161c2ecbd951a4a1554b94601a0ac0b60bd51a385304a6fcc1c4f7e58e59a1af8e623c41947640c0aa967af598a8d29ab8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h850284e0f448565c425612b22f9a5d6973550f8c50266f262c9210cf1465c776ad5418bb7bd144ed4407765b19afff2ef76c09f3188887777241519ec6620390581da7eb6e618de0ec9498960710ab250fefdb5d16bd41fd1da4bf4eb046e5bc0caf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf85895642246b6ff286edaf33c8007b5f986677161f3ab7918b5f1b867c8e20e79200a2bd6eee90eda9c881b18193131130cd7d95f820c113565cfd51ea29551152740dc8d0014f0511263d6a1fe090a4f69eedce559d0ec033ba87a03850d51233;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h628b958dac19d2b39130b0510774812b29ac84a7f29b43da0ae39b9c6d15c3d80222c7f6c31e950d746b4ab674d4ca66f59e00ffd06cdc84ad82b42dc4757156411725163f553f632a2614c84d3944293c8076b7d36be8a91f52b1b733d60002096a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d632c276cc486759e55fdd1862752e6bf03d030c63d5867adf184d658d98702993c1ae118cb2c639c0acfb2adba9513e52746bf95e7acb64546b28c9d9fe26ebb9bfdfcfdd0580fd66f036603423d7c7a7973f98a335956fb4e7170e42ef5713dfe;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h258e7ba5e553dbd3e937b288e548cad0682f1dc109cadb96f2b8bfd0902dccd62480b4482f29287d101d62ddeb234cf780cd9351e1c7840f13be7fc57e9fa6dd323bb12e4f42321261daeb458cb7fc3a6ca1c13a242cf3b51a39f98ac2af83066dd0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2fd63dd4a2831fc7ad790017c630789f6ebb5518ec4ba91b780ea04ed76916580eee3df2d602407ffd2108c30deb178004d3fcf83407ea884e19b0323ef1906bc4a8bf1e3399d1b61047b5e1735a5bd65c7f3db3566a601445a215214edb63c0d9c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b9d5670a74805743c493075d3ec5ccfdfd7e7066ccfd4bb316f64909422c00214af82c249bcd9b78ce1a55ee2ddc20f9094f971e60b7a2755d7292d2c13d7add11a7093ace3f5288fb77edaf9400a270cbc4976e675b20c6e4f73e8e5f908a5f148;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9f3d782a7ed9730d7fb5ad17c19959a711231f69bc182d55d84494b567acf6c79506f279d8fe3447c9f47c1b56d360cf55cb7282d4c9a8403fedbb4e0b466eec8c9dce88560acf58ec6e237a07bd84cd5c2921a874e7790cad82c9193a36996e732;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9d0cbfd2d866aa3bde0d232a3bcb1b584c0e8d16bb571abc0725caad42e1d2f23b18475bf166bb9a2b6bde5ff88fc547906f2dceb94d07795bb45abb8ead4e2316a60142f1009fa40aba77c0a696d9a6ca0f66be9e505ee87d03112ecac3ebf75c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72f2c855bd4a025b3c669316851c876f19121a6e4d8a6e29de3b2e9e157eb17fe094a3bd57db36802adf9d8a338db28ce8f623749d0fd1727a5b64f2680987b51f51282971b18c885f9449d72f35a794335336eeaccc739b298ccf4692eb3bef0ab3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h603050b96bddb744a7c6c74d4e4059efb57545056cf07ff9d4566156cf7e4deb30d9ed6fb36ba2fdfa903676da9bdc36e42fc55666f5f8751043ea1a129da2f1c6d2a8d15b776c7d02bf0e356d8355e77c2156194f97e5828cef26a9306434200c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71c2a10440aa25b3258d59fa2d5cd63e3af23eaad23ad2fde49acbbc9fc9fa7081e2721e01e0ca6cdf065c21e6a15d0deeb7f7a6b7dbd1e95607618c62233b95f92df11875be32fbb95d0990209304c6b9c993d2b0469957e3e422f7c5a2a4a9c8d1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha216b7904d429d11f436825409bd8333c905008fc40caffc21f4c0be22c411e6901584591f21137ff23dd2224b4e80d25b4544c6f19e3f5f60fc5e49283888a90bcb9f12ab6a491094de762fcde3d32df2635238acbca54c2608656d1f6785cea336;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h674a3b13a421629b68eabfaed227f6336decba596667aabb7ca2caa484f0f057ca794307fcf280c7707b2ba440b5b979fbe39983ddac647ce3fdb963adbf53d057d77c331d15f82c53e592b3500ec394d8b595690a904aa05150e2833da0433a6120;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d350e8de072b31c97efb4d9b6f2885a4b0055e9088a842d708a4671a5d220631f0ca30ffd4a266097caae0df16f807a9a4ec9f46db4a74dca120988bfe201d671bd6fe3e06d842afbd103481d33f668edce6c3c83098088a79c446729451e427ac0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82bf098020f22a28423977ee010e99f098e3738812566441c0999f75e9c6635c5d8c1a458f19df855d987e607c43a8e96b080aeb710fd030321dab8fc11f8965f054b08a73e23beb071de964f12e7fa2763c83ab118ee2d9b49a2f617ec940d24c85;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hafbc8c0d0ec1896627e1ac3667c044c67e357ab2afff0b66942a42177376479d7e5d67cfe3f6225462b2fad6995ad19ddb9b6beffc71b27a6eaedad4f9042c512ae9aab43424880ca374cf5a23e9081e71d038a3d4cdf94dbfbf6d5cf7e91573e180;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64b195a79cd5ef12178c4274b55cf9e4107f851bc5304408a7902b179b704c6ba46274eef23ea6cd02d2bb6ca489caff5ba128e26acf3882e730d4fedc1cf6350bc2997251074cb81c7a528103888a5ab831105cf9b186623fb0518c9175a71cc62b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5908de55afdd995684074afa2e31d65c94ed097d370060ac1be6beb455854eb8a315e0e458efbddd4be019689d5abd77665aa53d1dfc5c6e1ebcc924f10cf76338409ce43e4762d91a2530174a60bf04b5d2e2e1f42617b972d35d19476333e87874;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6138d7732990f15924f1f8d02f9fba631c8cd099efaffe30ca4a4f05c8b3ca702d3175832a0ec61eda61f23099e5b5b5460f135641bb3f7194a29e46449577913c7a86dbabef9602237aaf82db887fdc89658e9c5a3b00c3fdc8463c0a2fa8d60b47;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8053f803764c674598dfd2e3ff06ebced0bef1166fa4553843c737ad064defbf328320b221d965f05f552e83c0016667814056dadaaf5adfb17b410a452fd9db2be04eb6efc56a20a09e17ba57cfa71991c5aad7ec20955c286bd2026c1c662e33e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2a595ef4aa7cedd0a999350fec5f25c0145eade514d077d88d9dda2352f36c63bead09392e92a3890751280e3b96a53bdbeac2d93ebf8708f0d87a9535df482289c7ff5c6f834a27704c2458931272b4b6ea640a9207e33297b20f39026d5d01a81;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77ab5ec58fc9d2039fb36b27aabb8e27f0881f9f3f1a9cefa8a0b630f28848bfe111be48401f6e9e786367132a5fc7d86a2a9fc94d39facb00b609925ea68219b6f77c9f484568a1fead1415dc110546e6b6ef909cb0bc5ba31856b71e72e3efa3c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d6cc8cb0b2a867717c32eef1876ac96cd0c4b0edc6f3362b3f894428f612ead019aed4ae5e53490404388171c2721c9a9c253f4b3acaff14e898d5af3d95e89ad372c55819b1fe790d691cc858e21c241c7aff7944c0658e411e5cc15b22fd0e2b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d31b9051d3ad88b5c33089ba9124b5de008f3fcac035dbecec1a340b5a1a77e83de35ebf7d1ce08f77761f591527fbdb3630f13d519b4869c87202d550a88cdb0fbb2343da8fbd504d702a0d2080e65f95bca5d9e98854e6ae7768a8af08a5f2da8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36f9eb9dc4df75d93aa0bcb8b46429d9f652d85d86555a8b5388aec2c691e60e4f5d2b2eb9539d43774a699ccb5a792c270fbdaa3badcbcf4a9e5e35c567df99391b2349b904085f2944994ece6b97ede6afc28f2c5ca420f6bf9406f1630ebcd106;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a4cebad6d5cebad219847b983e8fc99ed594a9d45f1764651342c40a71504675ab025a2242be50c9c56bbf1e16f20518a8b84a1e30b3a039ac6fa5f7b42df53c186580657c8a2763494b0eaf4763b196f49f056a8b4eebaa16e07ba6c271790541c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b6fe1d87f2d81afa1678e12359280075f4762477e217f3fdb3fec91ec22deb035ccdfbbd7f3278affc729e942a5b98ac49479891d1fa8e605b7020ac3522e4a0fe9eb9d877f2e2cac3d2840f24969175b3f637a5f19f33f7f888f6465381c66d59e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h878417cc21bf4188a354f0a1c84fa81b10a40c1880969323a61bd479440d54a5866199ac0445a915f7e63e2d02d224bcf4da47600379df613518beb2d4106453f78dabdcd1ff8aafdcb5f6caf531f51003ce3310f72f70ee9914de15f4b35c7d2722;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2bfba3303766a6b4a55dda362914e75619b0b78cba17da1407992795c4d7cfd71781f9ec1f14f34581d3a80e5fd12fa54eed1521f4a82b30dc7a9e6d27d4f6fe9abce0f01bc3f02675c69c91d93e998546771a186acefa6c3b466984cf5068260ac4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc68d5a09743b4c2d052d249b354cdbcbdcd0ba1c371a52559ab94027bfb81773b98ecec25ad62bf6da8b33903f1c743bb225ee0602ed195f80ae759a781de5659e2adf5c6d36648fcdfe4f102bdf30736f773c1604fbfe8378de1b94f838e7604f35;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h165c9ab57839ac04264cc2be387d61d3acfb800a786cb4fc40084b2d4b69d48b560acf6d2279eebe383dce21005fe8fce0fa7ad2e14620e197433d1582c491f9fd8e80b47bfc23af48fbfb5c76bad20edbea6ff5aef8549c6a236fa32b95dbbc4516;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ea45c70597be904ed5fa8d5ac7b5fe2930a6c2fb2250dcae61325f16c1d8f886aad8f871d4e12385414f86564307d084b573fed8b53af6def2c620557ad79a6a1e002c4952adf4dd44e41fe9c13abd95a76df5afca83de5e50a0b0649a3fe5218bc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa5b5b9e14138893441b641160f6af01f1a22306fa665ba03b955bf90e28805adb64183dd9a454f8b2ea3567a8c6e8afb786ffd622579fd058abaa00a6e46f716de76e83a50441fe4d167468a5997863d4a4b85e04d37d96954919a9e7e251e4f5af;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a38c76ca0fba58e9dd4f933a01ace68a7e8f0e72ce35bc86d9e9bf150210748db1dd7c60512c75fd814be7dc3b2fae3d7bfb9546154a01c41f830005a71566df2e1439a40eb48f142ffb45d96304823dcd9b083bed470c7a485374aa238ed4aa0f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h172e6848ca6ddf8fcff685dd8b049244e40d30d8f9913220f4adb8d98dcb7eb393ce624890ed0be69c58adc1430cd21acf027575105b094ced13dc9e646ad131a6ec44cc4753a3d35369762e83a330e64d3089fbfc1c0dbfa34aad38d5f9dec111f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf35a0ed1347089884455d340693636d361387fe575c51d28129a657f5e089646843308e83d7ec9ce5f6efd6f0fd54738335e80376afd16146ef173390e2c5305f23ac21cfc6e36f0f54140b72f7cdf20ebbc77dfb40c4743bdeda5b8c5fc5a85b09a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e21ef0735c37dffbe479738b7ac801550c6f10796eec5962702df7369e607ae71bd021dd6d349d7f423794057e43e35a4c429a8bedd3fde2036aa403540f3b1059fe65e69076d887d46560ebdb91b3346284470e9890af1a2743a73e184e9d12dc7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h127d497d8887c2bd3b7553287be7d6c9d06defb0a86da8193b03a0c654f0ee1c09770e20b141eeba64dbdda4b074e8c62e251eadc1733fa7ddc90cb27eb8e99cba96349371df0614e50a2796f8aa2c828f98191f017095e9195ac9d9421e8e029ff;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac326fb3d77361a80d3232bb81aa3561a381b843f9c0b124700ffafd55e09f581f91cc35cfe0d9ad9cb8d421bb270e17b8e0d5facc141d88bab0d156693adebddb9da95425c3efa9c02aecd96446b587219637cf71686921ada20ab11a15163ebe10;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he65064493d3683e12c22d9d5e1557877895e8b673672f25160a79c5e849477c7befa1f657986dd6fdf62408d37e07685d6276752bb8345e248d6aa0b76948a4cd01bb32188ad5ce664348643bd5bff916cf74a6ec6c4e5745613d54194fb6acf1d72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9602acbb841c20387361187dcb696f730929a72cdfdd992eb4e0d786abfc34228d39cf7e931cd7d07ed924c7cb8a85b0cff0e4b31d69df310a88f2d36cea96e5b296cb77b118538d2cf8ba903dcdfb5a2d076046cefe1922a2e99ff2c0ef078887f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9aa128b109c3569955baaa76d986f8bcf6e1e2b45fb9e0b5d39e4573ee72dd92bb3a1e0a2067333b9ed56a7adb2da3198d8479ff097a75d12821c3ed1ba9081a874c116a03d9aaccd412fcebec14d58e0430af74dcc72dc5b7a7d2012b8466a5192;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c2dfead8dcddfaf770d12f613f8e238a22a657d3a245e18d1813171e66d5b97114c80654cb20b896fe98a373223abcd8343ef7e3f4b7c3552f2c5cbc13bb74e14702f8fed3ea1327814796d0622da3c66e7abe468ecc579b06d2792c014c49d57cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6be2fff704c29330196f07302a456989f17429976a546858a522c7079fd868271a4f01e1f4bf3ac66a5dadfd10b888eb1d6a7a736f3c76b00a22a80f81588d66dc2f732decb2860e55178dfb356650566e3c7355aa621689a5a313353b85b5312eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29e9f1ed5e03524f5657e2fc8978ef483da1beff5a576d1076ae48cb0a0cd76e16af0e5efdc0eb35c3beb6c1ace0110b16e8653f5977a5c7dd0c3ad38311a827d2004a190aac24c3d147b02cf04f792a634714f9323235738794c08d24429bfcabe1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6759bf5b79a8f374e50db93c75a69e97b908e883869ea077cf2364ed653d7445164ef445f60d8ac83d42554af7a516534cab60dea82b9fe4fa6d3116bff33a0b7d1f1525da0cb9d36f1392b96b7750b28a013f99ef5a304fef36d17816af99e4c596;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58417ae51bac0bb3a47ce98d237591b0356538e7a240b6065c4c5b52df1443426e5e036d98aac9d8777cca2d798825ae682f365bb46e82b0eb24e0b5c88520bd5c4a4df5f5575feccc62bf8c2803588adfbba431349d266deae642ed70265e147ddd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea0afde7cc4ceaba3cdf0652376a56e1f3da215359e5ec6a8403746c4a172da15f1ca598b9e7c2980c481751bfe7a84328b310e50d51c874cadc1283bdab7a4d00329e4450438c6a2d9a80922dc80148899f751e47b8d1de2b1be531c30a7acd4cb1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd852ded52ec89b259f7dea7610d06f2c2aaf6397760d12ec565078c837da9752aec33418ba606180cb2d597dd907d09114a7c2972fc9841c8bfdf739d26fea6176ae8daac416401b523429bc11699818c1573a96cef8f3e9f4ee77b18eb286557bef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he771e92de0832494598c311f5dda34e356e43398c0729583a17d84aa125ad77906faac7e223f0235f49ffda6d73d0320c82c938e7de010e155db195eb6f542fd72eb0640a87dc2a55a2deccd62b93f2e736a580190d7550ebb4e8364310d86886370;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd159a43f6f74de679f086bf85fe7832a9c70dea3cd7ec9bc11a9898f5387b91cbeac5c3a5c9a13c2987babf1857ea8ac8bf64f5acb39bf13ac7013910fdd0688dae1d0527db2bb8a1031faf5abfaf8cb89f27f0c3792a879c703ca9099a6d728d8b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdb4459e559625fed2b9e6a4d2120dc093d4c3b8e600494adbd3e319aa5ed2fc4a512e9b97f765210b76b55550acbba49d7faadf565f9f72e4181af455710c84e7a7a0869a09ce4041d4871cf15447189ce6c0d66c99daae7bfa7fea9da412990f5fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f0f1219ccb1ba5dfa8a32164a0d7106624a5cb4a524cce79c8558e87776fb87c0db008f2cac9e6ac410d17dd591ae6a44ba37a0287331bd3b5c4a6ead755edc73077b08cd56a882533b1ee39e00468507843475fadf7ec6c304aab726197e171873;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce9b43816b86e27b07347c72aa735c01b554fdaa1e2c9e1a3ac21516643f92cfa2a166825892cd3a7193edc9d6a854865a3442111b1369a334d50e9cd98cb78dae7087b06a493042840da97d34109b91dbcb0bdaf0b03f1710b53b8561aa54f33fad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5238dc68f4a9ba80e0d0ce6d72da4929ce41caef49551603b2a3319c445f6434d6bf64d7cfb624a7f2029f2dc8a563b656f566787109d55f758bb77f0766622ef8e1dc8a04450eb43b105fd8f017ff5219388ea804f709bd22fa27739b8185e43dc9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53719432462aa9292462f1241176e58d9373e22e57eb313fb6ed613fbf578b5c378e7c0ec358abe85f447dff845e69c8ac003da5972f3e8651561eecb4ec915f9911c735e429a2bd5dcf15ae593fd5ca5caef1212f4531baa34ece3c2603e26df8d7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b5476f478b2628895a1fade3052baee79d7d8d585723f5336ec54dac81a4b0dac150f79aa264c54fa5e9ebfb4db035e0402f9f65f3022837b22439ea949de78f23ccc9619a5861f7815dbad5b7771105abddc7537f99b96668a30f0fd91145c38d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4ab0d310acc5e2e53f9b886523d12984b2dca34bbe1c6668a4c43446ef92f5feaeb5036dc804cd5cecdbc541f299393badbc057b728aa469cc79b5d2f8a63fa7043c7230c40e9fc4c1a735464bf2498ad20e81cca11239864093f5d65cf0925e10b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h229b040e1bb31ec1066344793e16e6c4e3603b601eff850dd5931cb22728a3bfe97ce6ee78f871f9527e078134b75865fca2c4329aa8fff38ba44529bbbbf33b1f866159335bcf87ff7bfdfb94e0631b8fe1e9d20f673ad4dec54d2d795e794e1b4c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cb69667883ff3922458ebc6e13d8737f12a895ab746374ae2ba96c858b2c1dfe3d3d9324e8db8d97ae58b35bc573245395b7388550c5c2467faff2cbdd2a2adf11b7d8e5c7f67007f4d67de05bed35505aa1dd5cd94681861bd98858977628abf3e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he369c77527e0972078e4aef0678067e53b0d73070d59f0f8c965c27f401fd9c77e52959ba5ea91ef3d41bb07cd967d890017f282cfd5620065ce332d58623e827608a9e6e95bdc924e59f47db2976bf062b0067be9f0640c8287a052d542b88e6d28;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8aa4fe2f3f5f35f863c004536fb2e7b4a0396b5278befa006231a364df61f167880756e8e42f564e4022e3409adc976524c30c09cf1e46bc18b0460759bc48a66188f1914113d158d66bfa01e04afb707bbfa33cec6e7f69095d7c0b245e07e7e808;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37c645ed4dd234afd5d33d9814c9151fcd20fec40a5a9f37b5ed18245616c4510224cc2b32b72da8764dc8c3cc19b4a4c2c51270f5d46ea95689ceb235d4311be4d8f349241dd34823b70e660574bb6bb0193a69e3495d7d94c5d7b22ed9da5d69a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea3f90516e43301b1b49b0aaaf6ee27be148faa81ebcf1a872d6c4f0addfdac83bb38f03536e751b9fb963f70df14309e456076dbea51e24633c41b8a06a98649335d2fff9e59b51164af82dda0a2dc5f56d8f12da5f55b338b97a2388fe778755b6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc85cca9cea815d9a7c72e015cad930370b0e4fb6b266c42f1ab26bd270c161a5bb2df4a0b0410a3fc16b9d258dbb69338c346d710b6078b130b50c6bdc0e543328733f3075e937be3c3ee9b68afc39301011c7627d5ed638b87c758763cc2a4e0d72;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8dd101a14f93cbfb47f88c9b018d94b7cbdb7e76ab5416ba29ec9870e3e104c952687338230f4608e2a15f3f9386fde2a4aba7e71440a7968c137299e3b1d80367f15ea1f7c533247e4b53c70d7ddee0995f0003497269b6a3a3a20b69471ab4f9b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfed2df80f5d14a5456f68e502ba4a33c2dd7da474ca12156a61c02d9404df03fb1a9324bbce498cd1c818267449e3e92a93c8d40c684729d752b3be634da7b0e776c64b0a8fd5f57fa41e8515a8249ef240e313b5cd86e00a5ec3657a2018d51ad4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7dc32aa12c6fd3a8a6709571a0fc3715f9f9aef969de90c01b061fab8de010d6f4cbb83641594e6f5843cb205147fe8f599c5dd2cf76df73a609228e5624f3c7dbc72e63271a5fe7f8ea04f764b64f110769d6834c44e6aee92e04447cd7405870dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd59a37ceab4e38f29e528c0cd1ddd1211bc407f464b990f773b27c8c955b4d069319bf9c1d888b98bd749952304e3c4b0322f35238473add4e45ed975b2bbdf492045602387a77f57b05ee04cf8534da6ef3d8be0ddb2300438a2b946fb0680e230e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4c8baedb2b533c8d0f7be15da1206d970a2d6ca5280212bae3810feebddce6c3b604d4ca254599f8f5f628557d92b8c9c88046b530df6dd694073a7bb244538ca41b24d4d98917d477bff594eab1241b8fb366238301e2c8ce0bc5f6626fda5dbf2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18dbde78fb9730489d72c77e98326a2aac43d2e8bb9efcba4b1a69b2346eaf30022cc83eabf4f1876d008ca7c7d93e1eb942d38b6885e4cb09f82e51037f03b3c0a8113da99ca267ffd345758794f6b8cfa2a92ff6c49f3b87eb927e459fe8c3b66b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcae28efe25ceb3f34b4c80bffff5709c9f953429bc1edc45bd16484bfa3929ce96164b9f32eb35767246b171097ba182803a3473651f4630178f338d660ac31dbbb052bb157137dab6cea8f4bf2de265d91e0d600416b3e2b082db471d77e4ec2b4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bf1366ee6acf2927e1b8cb06919295780fb42f4afc37d9e929701923348fd5d59c71cb162a039bcfb54ec42d4534b36a2d490fac9eb647978e1ad713d7f1c3870aff9f952f0c158c8436e11738211b1584e4c10df69b6a37983899bde403a28ca4c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80785f1173b8e4b607f8761b64f6f47ef7f9be142b66847c4be160f1fc2738a82a0b9c21a2ab5f343c912206f12a3636cfaf414f2695b892c1591a0e9e66817ccadfc628680e0cdb142e56723157043a6c727c3ec7e1a606fee7a14d86c2ac92da2a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85126ec8f996c5500f4f7ad94da584a5397811f22021cc10c5b99d3d3f37c3c0ce57697623f9608dc4b73a0e6de72111cdfa1a47960273c263e31fff1ffee2e0fdc771399dc46179d66806f080b2272c0534ba676718e87ebbe7d69adcd27ca5cd37;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb075ba9154d8440589352458dea317703b13c87bb05c6475e5e1e076b108a0c4faa3998400fdb99f9c9ecc34c5bdbd8b6138d5e15d2c949eba3d1c8a4a55e32380c5427ef4648d86fd2382cf24b00ca5210856234113216db3fafebe07f63553d7b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a6558d1a9b9ff9d26fe3340bb6beec4ef5497ca698a67b7805c6b7d22ec59e395b0ae32cc4ef8153b0a4239a1e5758fd6cf874ae5785958c50511ce17fe1bd6654dbf88d70ff4e800ddefad643e2a903834131cccd54d5225340f6408477fcc874a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h625d29281c54932f0977eff42aa1c61a0799c96ac29d48fe8aa955dcb73b7f18dcf8871a73828f2dc43349dc5d0642593fbb97445216a4a9437d20e12a91f73f7f71b5ea9c095d30d2362300dcadbe0799735cfdf362ff013d70600807997611f734;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcdbecdfb67fc03bd04f0fdf954a80e4cc14134356a8f81bfd7e06d67c8b6607844f0a799524552bea170cf7785d020010d39d13aa207510ebca9db6a570a5b5fa9f209898c4eae0f7bce7254ce27ce77dd52c52476a1e47520706504b5082b4519b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb5c36574221903c0927edafee5419e2c50e90a04d1b96ed334f15f9e78ec33a9a0febe5d1466f73f6d61591b356292f6a8a348f3af4cbbe7d7d2098c752cd394a470d09737e6f0f3a84b2b57a67a6379583baa1d470468b7f94693f97142fc9965;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf2d7476be026a89597d0cfc822e4fe6ecdce5e0a62cd22955e4cf5ed4ca5e8783b1657be838a3b48c3d38d229d4b3ddf03a713868b621dab09f0f11a8666af95358fff7c84e27be29806bc214ea5793f77db349d94eb2438c0727fdcdd7a76d0d27;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47790d6050d6f79130a0671997fe76d04c47178324b002976ec958388e5ee3e909f5e54fe35cebe753482428eec42bdbc757dd0cc06b2f7c38ca5b51cf1cfaa4e8d001203e3dc3342e9c588b4d71eec9ce2c2db88ff892898ca0e6df8c75ff0d6b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h162f3ff43905654be10b19355c77c7c04b08dc48033c62dda38d49a646d5b7500ea6170ddbecf9a22bcf6d0849aec713afad9bdc7b87f03ee6e7ef0b3baf42afe4ec882a299f26861592b075ae879d2ea2290b3cda5127777a690ed38894e7a2fca2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e1ad44d33c77c07e8e5da3e49b77ffe538d5962ab405b9288d7c711bce63f7ca2509ef23739830c329902c3b6b0301b5d541eb8229e9472983b640fed26c5bce712038b8e87123a1fda3693624bc385b2959d5892bea15fdf749f62a45e87d6f37c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfae74a1d283185befca48e087aa2571800ced84a3ff277fe9ee2a081cd40386c931f8227f56eaba6cf16dc8f97103af44e28a176de9d6b389a7af5b3f54fe4f90c5272b7ddaf97c7101b59b8f60d8040dff79d7f66953b17bd267d037fc679dd88e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h842dade0b4517607c98d79914dfd6d4d7e55c3022ba4a8dc37adbde9ebeb686aea05ee6f6b3cc534a93e23a245b617e0ae4efe54a9a6099b8c76816ae441b6c6a987189d0bea218e50f724f508178f5fc4298da108f9eca38de4d1c54af13dba9934;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e50253e0ef45adfe4e7b4e5e08c7e1c32eba4b75d11bfccf12c025977f65912e2c6352c0bef7b213b7aa80a99a43860aadd341ce82c2073cb82999d4147e00e381777f7abd644a484ff382c231982fc2e69436835ca9b1f0b2503d7f266c1585e9a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he646e5d8a655ceb5be91e31de4fa36ad79b21c2c1af11fca96adc1dd6a1218d885277b9ff713338282f85fd5e3c186ee8c857b62a63f1ea05f8bf28634f12a81a2b23ac033bb26372c683fa99ea6ce048304fefd137e12e0fd4633e7dcabbe243c82;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22802bdc979e81af55834aa0b8a7500b220144aebcb88773fac49a3bb734afe34ec56ca61586bce26cc4e6ef0d2ede3918fb511a6b6496177bfdd83cf77da6c13ee15f01330d59182e623d44e8cef4d3d322fc3bca4bd63e6196adb9be15f31e1a1e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b328276f4f2d20aa6f9cc17e47308923bf245436b75a80dc2577a15c771a92236495603edd2212cbcc5836b05bd330845a150fc645f904eee53a3cb7fd0b867fc30af7c5831fd3eb6022f87b48ab114a077f82f82f27e5971f97d1d3d403930d854;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcc430119fb3a5811a80a8f677a7db4a62b131139c11932ebcf557eebbf59216152d22bfa0e9deb406f0bef39d1c93e7f089bcf3651b699c44ff4e94ddad327369646ab0d3c6b21b5b48f4042e8697351b828ef93d21a0f01deac214c11aa06e64cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1250ad263102b81d9fb6c462ed467161770f520e6570dca72ca23466ee183af00aad4cf9245fb1c0c5d6888f5d5e0fa4f7f47c56dc1711de907d1535984d7c4f4af1069df1544113585cc8cae3360729db9af56d19351f31be37684b7ba0aee3893;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2faa8c311953ba822fa540bf2b769f095d80003a29c5de0bed9a6a71de4a1afd68fcb7499dbf2dbb96af41a721f5badeccdbc50b6433f8a1ff6dd10558f0bc08daa28c0a440aa97341037de9349361f2eddb44cb9ab5379311662847ded4a988fba0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c3e98dc894282c2afa4b520a58e093e9cc212bec56c26d343ec379d72237187422e97def8dea1c2c8f3e4e3b34398fc947eb95bb546e6f4bc91ad2de741837e62b1a21b6ec33386b453b8a7bd7539bd3b8ffaaca6fb5797231792ca2f624a9d6de6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcea89f96251565ceb38c5bea9a85d8a9d0d78e614778cefa68dfd99fec3a314da7c37f645e80057d40dea02082ad20ae5ba321775b80c526eed2cad806807ea546b9db13ce8907e2aa0c84f6adba1d49d99db7b8ca2206861d82365bc175a62ab4e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5af96ad003160b74d3dec21a215754d7ffc12594d4f8013a2f9487ff176d64e77f89a335f57dee1747f9215f45aa2089650aaf37859e6b0a6ba46c68ad43daf759cced5b90cf787cecac4fa25f194a1e1ce26111c1f5f0a129d06344a22e4000ce31;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19b07d7dedbbc339ad7b79101066f33084a86dec6edc7ccd27dfc36176c2621c567f2a59b95a69a0bc21e5d8e360433665a645dd5d046fe165486472ffd8bf69b9eb233da4c7c24b40c456ae8f3e0879b344beaa9a79019d91b00df00fc7a5cc87c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9700d010e52eceb4d158b5e6c22955f390eb140c47fb7660fe429b109b18e751e2796382e1d90e1dbaceed16330f8d4c6532eb823cc053312ab457461deb967e452a30562c5492f2a923d1e6ac6f7862ed39d5ab9cfc6abbd58abccbbbeb1d6a942f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe50082fad3ce0deabcc6973efa2800355b2543f34c5e0e4de96967f821a461f01bbf8976cf7d4d6afd31e1447b3c111f0da7bbe59b10e1f51fdfb96914c7e7ca3f85477719a0f25daa0cefcf0115df9141c87e4d886599dd5a355043b702027e68c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h53551ec4333a77849b5712f9adc0c9e176999ac05590f937c30d51824baee6f72f13c350397624a4dd158b656786f73620e4fd84f15ffe459c60cc6960143bd5183b58fcf443656c5539049fd7464b4dd15223072515806d910e2cb83864dc7c56a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb7db0cff949e9e5c6d21bf5bad9edfae97397874291123dcc8f67e14b61ea688d5b54777cef22f7ce820158a520c79041b00dfb8674e53390f4f8e97b26992bcaefdf7e690c25b03fb7d70d71cd786dfa3ae448b6a2328d6d4fdba30790a79b15c2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8647d32b7ab6a8ad392d4309b70387075abc03db182d4971e44444a0a557b60c8da7be1e7cd14fc46e31acfbf042bb05940114ece2a3b73715b129548a339dd72b03dcf7d10d45d69d3bac104cbde5485e85776877a6df758993092197c7a2e947c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb33b500f04d0ae9cd0f71b99b54557fc6b5de9d9c31817448ef18cc3404602f0146d1a7dd3e7cee379f5b8c2e4a07050f88f1e37cda635963f50b63c9093dbf697817ffd9a7fc6014907358abea53fd8c6293553532d4ae15e0ea1d9c3775873bec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3896d311745cd2f135a0707711f8a624f232b5753b1b87cb60a0af4465f68aace14d74b5239e1192cd8d1ebafe95ec4a2e7ac705dce170d8eae868a7f574f10e359364387a884de8e55176a047eb8b2307ceb20c3f1a2af47e6aefffb48384083d97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2c528ea08a1d8d1e10817aa2ce6f73a8dd11aec1d6fcf6413606655fc0c424377ba232b3756b0cfbad433bfadc32ed196c0c3febd600852bc264cd0370c6ee2325ef07f990b054bfaaaf6d142bd8db0f1d6736008e6e02e3f6e738bcf1c457f3c3f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83f2846605ee16e41178548f55b233346ea01b4c8a6005825241f500965e4ba048f6133f1bdc0a0bee7188f4b9dbb649e643159024dafa03d41adcf2fdc73dec85fa7f80f62bc5905708b9b11c055af8b19f6d934e8aa81507a19fbace78f86b7c5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75b724fe66624558f82cd71a1511635145208c74cae897495a1712ed4c021a02e6df9c60f3bde43d0a6679eceda54c151e7af905863c9b1b6c79cd052444a7f910bc0935e27493de262202d06d179541a1a3de81a39ffa0fc0eda82630cb09d7f6fc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbba34500b870cf8b54ed7dc2fc1b8a52de2df8e3f3a54d05b671fadc7f66501046ed3144ffa048bcc7e624d09cd414e31427ab089e8ee5f3f6a87c5b185fd65008031beaf0b994f80fe3d5fd53b3f4fe43fd12c07dcb6b528817ecb11ef42ec15050;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7936ee88e3057a273bc25566a30c49e912c56f4e10a52ba59474e5fe4a8c430caf408487415fa76b3bf16ab19ef2cd73ee9996c9a10b94424d021c9a2e6e9895403ec2ec384c82a08b68bf37f3a333d5811114a539068156ed337ab1dc96a654c4d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1ea0bcad5638e11d423115409ba6709ea21fb89a5eb963ce71dc65c643c4f76b62bfcabd80e6acb10d1db352a67ae8c525acdc05cb2bd9485ce4dddaa8442b17c607345387fbf7eb645b6e3578e3235e6acebf68266a30e2a47d34a81429f75d5ab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc47e3119bf6e322330772c5163049f801330ca47b98c2264bd770eee5238ba9e86e8a66b59da9e95e14cbb75d252f1ee0b5b0d5b9f103ce3d6dbac155b8cf41e2145bc52d1e4f40d7cdbe6d45b5a1789af390fae8bdee403d350ad33e99bf71fd37;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e3e81866167bc5c384e24742bc82ebb33aabf9cd71a3b37e9f152be9f5766f50177798698cb2ac836ccc96a9d6744b8051999298fd79418dc08b0db66dca8e8da91b2ecd16402b9036d6d46a9629cdf8b8a2782477a84a4a745da24138b58f94eed;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1eb587ccea3f160c504b542ebefb50994ed9dbc507bc091a4259de71879d0e757000db37c8a0378f12e35db2265a8c7e36327a88f5f58ad959f03242da3d7ce2b717201d117ef65344554674c40220c2dac9a69a6cbbdfbd5610b5500fbd91bd0483;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha84ff8c40c9aad557251b6d560232236a894062e08328b0861d2ad11a2d75e0079aa4092c3b076d8dbefbd39d58323ab295101417c93e411a0a2c74aa7080f1b668373a00e289e9a2e596d613a826e7ac5aa13bc3575500c93b419e827a9ae147698;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8817d5b2e0dc6664259cd5e2266302b76c94aabb4a757a3274e68f6ebe0a5ff07a0c1609c1cfb27d34cf0a7637e64cd9dcc3f7cb8f36055c67253e8aa8949b00042e57216d73c9be8bcff98f3a957f65eb54537a036efa285c7d591ff821ca8f2f6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd57dc4b0430984f55bd20419d946bf57532f37e912ea4cbc4f24790bd908968a1274c7960efaa7b708b266cc17d5634b68a76ea2939fb739fe5b790e3951a804f1bff00ab22dead32abd52595e47850d1da7f8e5995d191b472f6eedc341e9f50e63;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc768123966557cc22d18620c358aaab015161bbcbc0bbc4060387c85231c3ca92e59815203f1381eabf8d1c263f318e4a2cac7d42e66789e9ff0b5e7ea57dd218609f6a166e01b7e2cf3c42eb1dc27d3cc44f737153a559a4c244707b6d7260ef4b8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7da68ceff3f7ecd08250f9ae96396e95d36cff2f2cb03d3ea985eca2feb562bb22b442a9d1f57bd981e7c2e5db381e2114ad09f1298ac01b1491881f5e3a9397c496a9b6750da0a8129847be12e94d5f5c1ef6b26a41fe6984f7c75e4e315c73782;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h118349b36885ab147da40bc8f201a2453a389e98383b9aa044d704b68b8ec8781dfcd8364efb31d14f384dcb711fc3f8e547db9a25fb69d96c1aab9f5ad55338b86d08db6582aa5d07ee2c0fd58a8d26286f991fcbf0a4afecec821b617a8f6bb393;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd6249d57b2265067b51fc31c0a904d1c301f96275451b3c357d241afe849c256203bcab42481399d28a43aa3c7c8f06877707d35110766b63ed75513ae4e797e36ee2693b9891b05ddc46bff745ba28d1d52b5fdcbe49bba7066255cdc99d6eca77;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fd09b491acaefe4bd673963034741b6cf92ae5a3ab534801cd8551ae4f86054c0408fa3c473a2f91eea57944de256834075478cafdbd981f5e5ce5048425ebd4d7e8a8997888799c92125ae316d77fa985ea95794a43b956e0681a03880a122cccb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h752e38905c08cc32def1561e49a9703e770de38285b9cfceecb4b2d145f07dee2fecafe751cdc33dc5bf189aff524533fdfb9cf0131b36dfa7c059e0d06c4e850a0c77092076c9747b4ba7e2f0b1bb63f6202e184cef74e5aa95e289f271e5ef2115;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98176db097a00efd5c1faf8a557c3e9a12352f3e500fa8394da77c70d39d54ffe8ed1f0a5c5385679d4c4f1ebe46a8f25fef8f02bc658fae7dda02d723c6e6bdfc98521f82b27c95b1df3336ca551b9b12002f4c3ff60a8349f7baca772f24bdb615;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec406380b8ffd46132e30d9e961f55ad5c325395f52cedf8809f7258c450a8a1634e994ce91d629ccf16084f037b2ea48ac15615d6c9689699c99cb2a2a56deeeb5d3d707d4d238cd6e7b3e04a98702333f82541b4e77f8b2efd178c9511129e63eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf818b67a3111db9ba5b3a72b7b6db358e7bc715fb5aeb2e534afd9be9156ba7d405f3f4e9481f0475f7945d8209747008ed5930e3260fcae0c642947d2f7f0bf53e803af8de4f8e21a20c4d7a6e8af6c0e3ff6908d156d40c7d1cebb73dcb100abcb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h487a528740d66c4425337c50a133a64cfc0795456a4e26d7d240c7c91c3129199b169dea767c154cb92946d68eb098f1b500d50e2c9302f98d744affe3d1257b12fbcf6f618ac70a81ee4b82681cfd9063b21e3014ef8cdecacd0f443c741cbb730f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13f4c883800fb003f47a802731fcb4047d18454ebb4afde9532bab8558e8b71581108717fefcb89b44ca04119744fde74e7adcb833ecd5f2e2f5a3b98813a38745f2e4e0bf884ca33ac9a0e143cf1f90ae5f5786a19213c0c47eb31ef3b354cf819e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5567e5f53405f6aa173ffeedede37da153bd63da7124b946b28035602683a4eb8ed3f41d4cefec17de37768fdc796558ccbe8f787071b53be24f7714c7320c3219cefebe6d04545ecc90682eeb80a89f70c274fb184d6203eac324c04ac5cfcd0d97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3dee88c397ebe34e5ab89bf56299b086539d6844b413c78f0bd886818a9cdaae8e8e3d1abd70e83b8256828a6e35c254bc46783425cc5e4f7c453af437a52606c2aef57d2461821c72de1e9c92fdabb707e46c5ede4eb5f3c4e8a6ea863873bc01ec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a52b9a43b9eac04ac5036b199d8acf9e60e1420d26457aff2a66574e5b4ed3bd510f02bb2947d1a3d49269194620cfedb559a7383419804dd62ce30b7c4e3254970952748ae90705ddeef4856c8ccdcd442a448f99e1c286e273120d846db5e60de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf5c0bc0ec2742aa52de0254c150c3e744e968e50288a0be50e33f7e05ff890384854f1bfb8012cc0ae258263d641f11ee6dbeac322f72e7e24b8359d3c423c05f2a7913718e2c2ca5ace0467744773169393f9b1b43f678362f20a51a7340d319e9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he922961453761ab9460b1fb2dd886bf4f01584aae2d3dc80cfa884eb61c45a19a5dc6e1f151fc63efab4f24439a89e94d5c3c4dd19bc0df09dba90271b3ec1c16eeeacfaf450d1d91615ad4641f8cb6fcde05a1cf3beca083f75a64396ad43eadebd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c51eeb428391164f647a091c8db2a4dc5b57e611ac014823c497d1287cf940b62947424439144c25db8489d020c2bdfff8cf4d62c75b91c2aae1b8dcf28a7028370e346c3560512ac15c4f4ce846a5f885911148969f76ae533791ae9555bda1b21;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87a04bfa6a9a46e1830a9c8f49cf60ace32a3770000391679a8ddb75fd99dc2633febb00348313608986a46462649618bbaa3a3628e076db731e4cf83f7da1de7a9f8f6d843435afd25b6ad1397225a7a51de06dfeb892025c2aef98f8445dc66d0b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85e6b684ea83f2c40f13b478c6c15191b452f8f37c5f8987f956ee693ae8d278cade1f1d307198b63e856a9bf234f01b651fed8c167643cb17fed64d2c6a0fd261a0c9ed1506cce03a755b793dd0c703847c026ea999bb605e06b04d5196316a583;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42e2f97c0f19d3c18bdfaa619e071743efc1d9c16c4148253e13112257303b123e6b5d6e74627cbab268567981d42d63bb9df3b5c0135fdbf208646715ac0680209b99f1a1acf5cb985bc831e4266514ff4fc7c31cc8ee41936d6d3bb98f8c81131b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72c29f4fa58ac5f15be2ef98890208c6a54cda87c8f8874a45d3397a7eee587be36ec4cb58cd3232e505b660ad784f4c8aace7bf554b7f1b4b377813a840c33b1ef8f1c52046d6903e973a689320e81729c80f981ea446dd848c9082531e72ea7474;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b03a5207dda7115932cc2ba2de7ac987d6af2768e644961896e46993843de31bcef0c50c23228aae9cf004402f1c774283d9c35c5eb49a5f1a2a269d31a076f3a58ff63c267b594fc212b96fc48ddece28b03324ed6f36048e277cf15f680331b9e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39c81293d1bbba70f3166ea4de5c79a520f92f16ac25683228159677b3cb9a84b2b08838f8ea9c52ae00f11e8e21613207edeb93626ef41ed11e2f8980dc2cd11945f4de1529aa66b55c7a5800554e3ff42b671ea3bd8f12e77eddcd77a9f0ad5c18;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb31dda8a20c4e15748e0f8a02790c4f0557b555848fb39b6788ce47f76611cee359067f4ff793c1bbcf44af56fb038d22a32254c3bec31ceda17422d25548b30c49513664f57e77dd0cd7642a858b4da17c2ca0315632a0f7a91a64629043251aba6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5e96f950de84ccd32246d44f2cc7c0e8dc07ae559272dd5d2c8e018aea142bb4296d5b47a5a60907496ca5d84ea4589efcc18440a536c03722a0bcc67a594cbe154cbea9cdb7d04c6e6cccbbc3796fd99a052e50291387ac34867ea5cb840aed6f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd806660ca6e2f2662ce6da627856a59c1f5f15c7992af1785886fb188b28072bbb6b8d777454e0276331a615dedeca2a684bd19345b583300a7000d61b879fc8410ec7108dc90ce6b40c91e80786e8493014235467ec6b4c7cefaacce4d13370d89;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ae3ba2568d67a232c1121a54ba1c2457c15ff2ecceb9482ba98bb2cd33d147d74b3315badbc664262ba0ce70212e3ff6fa88bd4c4c210cca48db337b248fe93fbd322784ad3d0288fd3b70b95a59a5072e2a62d8d4ef10280dd5d71fe5947379147;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb3746402ced2898734a5d54df61797677c661bf79c744b166ee46c3e0d7233b4aa6f1a04b951d5ae3e942f47b0cd50444384de8005f4d5b97ad21c0977fe4b1fba6ee9cd7ef3f1f60630377a9f07a7d03c27b81bf2a50df95f052c9ef3433e219f5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40b8a94fa376e0d7cac6179c68b528cfafe7a07730a784599ff5ee32b8f1448c7a0ec88feb8e4e9605966a486b042ec1e101950ba084c0cddf4669db744d47d0e5017e124da0a745bf82c4bb6e163aa1a8567b0718d80ee5ea2f4b5d2d8785a4e950;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c399eb2a75e78d8f10d4c148d7762f6b41f5bb4fc72e6ba5fb3f619d3ab495d584048fcc98c312c59703d5ca74bd4000bd7a353a53cc172ca9503fd3782cac6f1a798ed11cd26e9dd7552d050e06777ef9c42afa6670081cba8869993802c54e39;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8213f2948a3f2a0d11a4314cab0d93f230d7e2c0553c0fe5d2b5352bf523daa5dc2db0fe93c58a39208c241099ed9ecac434b2267ea49b96315293dc314ca4fe0f1d5310d7619f7a78d564e42331c5311aabf8f546bfac8fa31d4a8f1ca74c97774;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb548459c7906f97f054eaa2c41ea2c1d48d39e379cfaf3a04f78af14e669efd90a0b1928208816ac0b7453c59b5ba9574299674fb660423d63f976bbe19d5ec761094e01adfc5dd9611bc242bbabf0135a0607ed2de1b48a770611a52adbedc00e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacd485502cfdf1d1a1dbbe25c976f8dd26bacd7facba2c1c307c61c8564e371d63374f0f973a557e7fb8b282415b2227808b6a9fd4dfeee61682e1b8fea22eae2b78011baca0630717b8dbba90703c25b020431798d989d0ecfb6164d04cd02bc21;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c97bdbf3d247aa47898f3166a326edc86d3f77e20aab70cac9a5e7ebab0f5505b5364665d547ee7caef5f230e8b5ffd3e505dedf3c981421afedaca48f03704ee966de3cfdc26e64a312679a813e47ae88b47d7e5321e5fc469e0e80834e10e0f51;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ef6a4b31851d4af9ce776ac896f46b923eadd89733e97ed496d4945aec0907fd2e0c2e54f5063121a4c5d7aed44c24f55a5b0e8cb4544ff3783d1e84760c82eeb97fdd75c7aeab86821eba3edb0dec1df2ed13438df3d48c2f951e2ff3ec62c264a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51926dfd8e214b1503c1881ce13d57e914ed23f5f5640bd153ff0da74ab19d41b17886b048c1aeab7c6a8bc55b6db001ebc762c14ffb36cf58ff0dde4ce9a3cf1f85d61a223715f47e827a69ab9cab16faf1520f59c5525eca560c4b693c8e3bfd27;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3ffb91880403a38c71deefe80acca1c03e1e5bebea12223331bfe6bc74348035e7bca882c9ca5dc44f9bff6f69ee871e2f229030395aa5ed2cc3a0d71a1488c0ffe9a45796b32794775aab8ad6cef36e433bd645d89253643f2ce001c7d5bd37715;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1c7171a8ba051c0033ffd812473ed7fb8050b6474d3a1102d3eb1e6a1286702974a97569450874e3905d6b9dd379adc8d6e80de1732a48db20e3cb8bd0e67cccb533105521b37583c547d6cabb60f0a73c515c411d4ed5737bf4e6474103f3dc01;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b8c4faac3e6ac6cdff26b330778fb0693a715b722447487a4ce6425d402648073ca82029985780188f119019b74755997ecebcb2703af9213701f72d0bde2ffac294c7a607a9f054b8d6713f5e9f9ee523b7ae43e24d8f8b574a643984a8e8a79ad;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2590b9ff1c9175246a1d5bbfcd2700f2a40fd928dc435c3c763cab5bbb82a0f266b534826834b0c64019b2d1a592b72f4556eb1030b92e695709b75b4f6f442af88ee2a8d8969b935dd58e81be9beb5dd3e053652e83102c685d7cd46f9bd22c444d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9ddb189e530a6d75fe50b6207c38b6e3be56a4a12b850141166fca87065de57ddab2e4bbf2d0d450777e8f696c695b1971a189aee271aa5d3d1fdd4ce0eea16218104e015fc462be1c63f68edd1fe4ecd2d287722e7788e31c3a1d6452bd68a2841;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h150b4f5216679dd2751dfe037352b01629c5bca849403d0599fca54b7ae9ab0120513ebbebc95f003988b236f217b03397ff753d8580c5a44bc990e978618a7100c542cc7913587a208c1a9966665d882bd2857944d8b5cfc55887581c34067be364;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h12536d4bb6ca595f44a46d9af4d407202dbde8b21a642533d09f5be0f9bfe11e5e7d55bafc8ffea5fa013535dc45de3d334e0b5394c5a7c23eba7e3da1aa32cf4e4326533fb5c2e2d1a433574b4199da1e4c1aa79fd0709a27519a8fc3d14ec31e45;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30e7674434edc357eb334ca8f9bf367c919ad7a16558109b12084181b23aaf0a50c3e55468adcd09aaacfb10aa808133c9c8dcd37fee1c121231789b5c21f896a2529e1caa680b22938f7761a9b987bf6527711c5b6930f8b98733bf130e2b3675fc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d19084391842ced59fdf280601e04f4d0f101c6f83f63bf266b126a6c13ca69409a71511401fb22ef61b0f540fe018ef6262e1710a4e23b40bf324d8c7d4c6d63de1285629426d2f40fc986bb566700ab447c430721ea9264c5db24f8100511448b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73b6da86f7218bcbbcde016e0d378d1043d64d1ef9499234a972bdd0496a4b0e41ed327fa256d0a80c278250c17a25fd8f0b0f2eac0255e9514290ae2c49bc4702438b1324d5fbb6a31773f6d4a51393562fc9d9d65a894d61cc6138e8d03267f719;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb838f3a7467145926879ee4a6bbe23324bcd942d956d25cc949e3f25ab3aecab29fb70cbb5ae541929cf7c2e579f24584d265bed9940e7677f52ca4729e533d21b9b4a902dfcbe3c79eb0759dc46f9b923aaa6f9aee8469f9fbf590a44b3a540e8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38e9604537273b23aa0fc2ed60ed475162b51bc9f9442be111ae5278d9ffb4aa4cb2af3967cfe1bce8aef3413a3dfe35bae7467667d442ee0534b4519c3524f0072ffa2781fc326ab933e369e838c65b5961575802fff5c4b4b0c13495df505db768;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1deb76d1ad0facfebcc6c4ecad9e3bc3354ec7d0de4435daef883d1473dbd6924817417383e579def401344ad8e49c3d2bdbe2cc903913e199013356cb472763d36d29fb96dcf89b871384f444a335ff13b310e01c3ece53ba517b26fe7eae8fabd9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc27cd985d85180dfff58a95ea5c7e7b84fc0ebac50cad34d16f0680bedbd62ca2a01851b0df63fbdd4d3a5ff2027c9593199206dde2b80874952994622f8e18606374b93c5d6498a26c6e69d3ec9ebf5149574164a58aa163e1e697e497c9ba3147;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4820510f590b3d43d5458ba390a1292e8e1d3163e06e9382023ce429c6caa85c0cf24ca45b1b25b238d9c3c6d1376502f5f58c715d758ea43e75a5f45e87784d7031ce78ac70ecedf840922b38995d95510f28824017b86b3dec8fc7bd67b9fec2cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e09477f940a1c429baf614f77b935fbcf557eadfd5ef3a0fd25ba64c5d970fd9507ef4cad9428e075ac126a510961ca0dbf2d33725e09b4300ed9d09fa9db4110cb929261d5ed6450f039441bdc845dba3700fe3f61b4f127f0e753f817e04adbe1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f95ead42568cd24fa82d9de79303a5d82c33d41ee2a8a1721ef73c5da0cd21357e265d5846098fe0def4210cf844010b3e91d5d4dd60fd4bd07546cb1c7fcd92c8a3a7a03553c6104167a817bb8b81c761a1a10446e4fd1df9ca48849bdc69be872;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32084bb158f503575d18acd2dab50e2f1559aa8ebba57454244132ac7e648e1777fa667e144456d7927d98a79a9915771ae75e130e0f355ab9344c39dc8e22a12bfe8beaa2fb3e3c6239b9544e1927a5673d1350c7143f4b6aea21a7ebe07e2cc0c0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5831357ec765622ae6ca303a55908edecd52dabff8ed2a1ebb0ba5e99daa47f0d2845768be449cc3706312ee0695432ffdf36dd426078886ae896a93fcf3cfca1d50790d93918e314477f9367b8176a2c0b92349102b240f23735ca269a2bd344530;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8197b8056b025470bf06ecbc6764bf98cd911ab36a6778fef2f3c37e06abef34abe5255d30adf0c338a80d8ae1d84ae34b5d7f31eb342166d1473c23db5ce7de92bfd08fd3411907fddc6c2abc76a1163a1c4db9808697884a49decbfd174ebd3189;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f3b70d9d107b80cc1291dfd4acf41088bcb88eae7182a68701a26cdf901b19ab9f4119fef6313abcb4e40753ebf13dd9a919c6c2566d728b95d09e3ea6354fa8e682ff69712f58c191570c815cbe66ec7eee0b471e9159d71b8ce00f381fccea4bf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fa3cb648ad62f7c8f6867d37c1ecf1b593039fbf53bd72edfe471a1aaedb29d7384cb0683618e12484f0ce39a8328e7ad30d736ab5d52db8a6c123e2b300115fc78e7dc585199abf481d4770136e8e56d91e59ef65d30360322ff9287293a3ab802;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6c8a91c3b503a6eb4701b893f7a8d80bf264c9d0442842b29d30040556b5f9ceb4be4fdd7a9f5b079f5ec6d29ad0a1d23eb4e59b70a3aa72cda00ea46231cfbf1932a22ddf74c65c5756202f76056e6d771b51e14fc4226415f037df98870a54736;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha755d92ce391734d6d89e614c811b8da3eb2e1bc7edc7e0bad60b3507a6b077cfefd528efb19a88bfc65199de683931662f037c3fbe2262529b21d258ea76b4c1bf587232f4bd34681bf64571e0940229588b6463dcbdfc53c429271de4bf5fab4b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8369c28c77ebfa0d168c7214ddfc19a08d25dda8eb91e35f02d01a94c2d3c598e27ae1cfdf0dbeb300a21209989478eedebc7be3962674cc6763a11b1964ed75e378f3ad72367db5559177a53877b2dc881ca7ccfc01e2a932555ea9b5fbf19b7b83;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6a59366c40f6aad567e42d29cecabeb4473ac72532f506d12a50bbd3c6c7b12a0c52217615a5fb742edf046634425f30948e7a7f82a28186b25bd808eb17e9a1c8bcc28f06d91ca4f4ed25b4fd793bff931b3c76c23a81a1a17b39f76a4faa670b7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35f2512cae7e1af608ad1c30baac221cb73540ec8c4f54d3df0289d7fbba7dc468b6143158fe02c5071e99326f5ae96dc624a5b0187d100b14156178d1bd468ecaecbcfcae68d53a5930223707cfd2493faf24b05280aefce8d096e4756feca7f1c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3df3f32ff3efe158c67003ed3088d67c22eab9b4ca4c1654061c679603d2b75c65411fedb77f3d29ee4ae28e2655022048f9d63bbbbd782f7ca9bf92482b43f58ff8676fcee93f94e46aa48940a8ba3a24fcafadcdb892c073fb5e1be9e80411384e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h839a3ffb588f3476b446f8306b8a0ccd4875bb9a61a1c489045bdcb63581e1794d61156d324d414db9a3e08ee65cad6786a905bcfc363b2876883ffaf5c1f7781f0ae8edd475201a7d03ba4c9c994fa63fab8761464044a9cfa59069bffce7b8e0ce;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3cce5c4286ff6178491ef528417773d62df58c506f53d093d79275cbe5b23a81959a344d8cfee5bfc4256512a69bcb1df26e54a0d1a354b148281c9a91ce7aa62ec6d054af7434d8d5d94f41451b5a205b9068da043d5515a64c5dd7cb43a5af955;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c9d3460d3044488d58445ed972e5600ceeb66275ed5009100126484872bd578c3654d61a439e73e117b87a9d7b7669ad75749bed9843e7cdf0cab39c113c69ecdeb598654912d8d4b16501397d34cdaddce1cfd53e23a9a400da994f278b855a79d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h46c504ffd8f9c2c6d5d7a877780ecf91692965beee51569251cea0053eca1d8b3d9a8b670b96a81deefba317b6bf4470a89826417d326051cb47d1532f124ec132096dd7ca70d5c5ef465f002045b9927ecd72b24de9de224023760d5be093319943;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99c2814d070327c17367d4616b0282b83a3a29e597411c4ddd2cfd8e266b0908580361b1b225e1d376ff965f8d6c50c2cf98c9d51c4a359b52864b9960b8fd9dfbf7d56d57ec21a688a55b9f0399083d197a0004d94151480f620015925fd9c0ff22;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18e4a1bf7e1f231344f1ddce0a6c6606d0ddac329516e3618ef238a39595c71bebff5d68e9b23facffbdef247196208a79cadca62bb04e1e4cbe1d3643df9aee697b723f7afc97b9e1d5dd47aa4db2cf8a7288950d77f218aaddb47689857e9a3eb4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c00e50b59cefbded068d778e6850ee0d8d25121c29303fc37b6bf9158c1ddf33626bd599700d7ac79e3bcab1011778674d22070a227ab58c3ae74326d91733c8c1803e5264504a16d05fef2b65e77374b44d29c0f7e299762350e33fd6b3c598482;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha323314c7418aab799ae1028ef70be554c84a52543e99914a120c1a6e74c165fe076802b1d42fa47d40c0815bf969aa7f075108035f04d425f3d9783a8864ca28b722e8458d79fd7b8dce4dd82c01a7212610eae4ccf7cffd18998eae44a2c37b48b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba53f2d251a3448240901dfb3b6473ff61f1009dde6f415703ef7ccd19e53b5ffe93d35d597b69b494f8e4c056cf1262d861a6032efda850d0be0455fad0b41c9ea4aac9a04003eacc095a5e151a3dffaeaa0c3c56ab792f544d2169322996057613;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc589407ab9c263d8c1c176bbf3326e18747ec23fe032a9e344df3da402d4b2380b8f0268d7dac13bc768a5507c1db896728b7f6d73472cac7b7198d460241dd6ae91a5daec19403b1b600a7abcb9e6bdbae17f2daf9736794b10e51f87da838b24e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27649d2726e827baf699d29a9c2c7f93506b21f37e61e866aed031c8c49c774d75fa05a9a1cde2d30c4b25a05b0288ccf538125d25585953eac0732a77512f6f2a81b811c4a126b59c2eaa01a62205ad183a267a25b42cad8e3f12510b60fc9e011e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b9330f7638c74299fddd3d74bf8fb54199199e3cf69211cce139c877f30ba0a503d47b3b5dc1dd53112ad1b5b451c37dc61b1985da0a8ce65057b42ef13b02014cfb2176defb15f18763abcea444f5e3a91d6d018f981b89df978faffd0abb8043f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84232edb8e991af3521d78a558276c644460aca622de8040fe957006c8cf84fbcf3f1f7752e4f7d2a514014bafe9a7f845becd5a0a2db534666b377358430866e34be2d1a60e016e18c4634c5d65434520d92585a7eda1edae88cf170c2d3003ee07;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5de0bd2d5a4928ad39c1fe7f1727364821e2b65b29e644cbf624f2e8e8a1daf7de389fcaad649dfc0eea55d57da2a42cf44d25343f32952e19ecb904924678855e7ed1915f122daccc348c06fbb3a1c13abca55fe0e6cf12af54489b001e605bf2f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d8f648611fa68f579c09c309dbf7579ed63026ffb4c21523a204bee3315413e6af2aae7e53c5f461ca2a9ede517c5847861b2b2719a1b920171d648188176ceaf1dc16efb9b6ade239660dd605a05250ff4b7d3074245f79b4c076b8294245912a8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d1ad1b6e6e4bb9019bfba52409ae8c1b6eb06f24fd631dec1a49622a916071ff4891ec11cedc95bfda13f33e61b26b0bacc9bb6e1a7f253d34645682926f0008f657389d60128d416865131ee87cf94973b58cc365c6b2c31bf7821f2215e68457c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2425ef4ea8302e002e9d41651496053da7534f964ae30df5f66d501609416e2ab6e03f4f7a6e25d9ed24da99f4e7f3b4fab66ef3540d7d010ff6b1c0030427b05049f0a52c18e0c7a13e61d939bf7cdbf9db25422ad1d76228986e65cd3d66875fe1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed29644740336b9b3970226c9e44d4e8879befff34999282b182a60de3f261265238f314dc61755e60a0f57416fb955883ac9d63a761bdc57cbe64901f57d8b0270e6250efd37ce72b48f288ac2258d86668ae1a59d09a1ef1f315c0e296f1a8448a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h395344e527e10475abe79cc5ff7f68700b75ebcb2d07f42fccc26cb186dc2df3b301558d590dd34a7e498814b62d233c22ed46596da80086d49bc7348f1543e4ba66646028a1112cf8910aa81ed9b555635360f007ec9d7851d977582d80146d039d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h788ed4417a348a91e892ba1a1fee1b02ec104d33b2b584039c8ecf978510a7e272a9a420098023a19f1e43dd98324f7e7379e7efe403a01709fd9d277def15d99200e624fcc3cd2a1078da3c365e337424de0031d989bf98d11722476128af870dc9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78b48fb9cd5464817d45bdd6155ac0363dc8a0b414e56e710c9404d19ff57b1a6a077e498debe3c28cee505d2c2a11bc454288ccd230c65d9c592320f2eaa82b4edd2b6cec71ff0b02ad15f50d6b2d942bb424de860591c9db44880c962f856e57c4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h879afbfe2572107ad4714fb1eabe75d05bfdfd8d1dfb35341ce4faa9ab335b14dfeeef7a87de55936758dd9f6210fef8bdc72db523febd720984b2eb391cba5d71f8e6d110ffc6d617c2088878fd890312a0a32d4f6c3e184b09225ca1daa8698865;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacbdada591e5c61f83df882d3f0269c59dee90ce241a8528b915da83bcb050379bbbc3c7f52bd81ef138a330aed6bb52cd2fc34becfb64b518d1067cbd3a5355a566527d08585e00acc6e88da7fc8b39a0d880591f8a9faccaaf1e72e4f9ed7c9cb7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80f9e352d8e020a66a15235e58ae7456968b949a00cc3fc32d945034098540b982a3008c309484c8df3ac43f186c0a997810d9f60bf16298dff0f24abe788ced7c577e79f33612d51aa9bec117dcd8b147cd709ea2fe1d924ecd4f52962867de6b8e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4da15009e57a0c359f69843e61fadf6d4002ad25d0cc6e52b54db32dc2fa00fb35a290710fd67c17f7bb9bb2324004b649a301e1dafae5d95fa71ae6a2ffabba243d9f462dd9bf54da9499d1e20c1082fd5080ec068b136bef9f18f9480b184a21a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a752271f8b49e7aed1ed1b61a11983dc307317946872d5de62a45ea19b34cde70c66a4eb9e8272e2d8fb12dc50b6422457af747cb3c2d9bbaae38c649fba21a69a160bdf4fc3da7ca854b8f390f14a1f351f33c4b5876346ceb44e23b423361b24c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97f9c98aae608e6c57290f80c0c8c674b5a8470a3dcf88394783839d4f1b6d392daba6a6cc001372e400b814c4dc7755cf547edb49da3976000b652674d6fc25ee16c360fbdbbd2d40b9266344b7599799e1401b40d9df2dfaaf4110b8cb1ec69e2e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d58bfbbf30de3f1feb6517aaae932fea8859df25fc07adf257f985a6fcf70e67c9492f4337051fb0b8bcc3435f78746db6fbedad721e0e84284f3a84db9302f00d8abb8a23b84a16754cc9f88b9500c1781ad2b4562a78ede0be259dff2d32ee200;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeac2ea0facc8ee9be840a521e35b2d8c7d9d2c9b153c293df53661a14f6cd1f08b8f61c9f327e0d40d5600552752a59ac2f6d1c8563f8e9eb5b3ccd3724f2c7389490d2cb8824285020e785aef6caaf6f704db27f28cec7323dada914f3e60764cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ff4b295bc7c4f5808c95572ed3845bb87c676cf06c4e3f9a2a1ab5bc62e0a28edfac089123ffdfac52b959358cfc0eaa2ea63010a36a91252d9967493ec3059ee53a11292a609fd7b4e32345f7a15d7bfa43a942f81738d35a2ee5c1c2312acb271;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a83ea3d1d62eb15f6413159a9dcc94f9d42df71ffb0e01be07d6d2c5a3c1d839accd3f4963c7506adc8f4ac7eda54105f89461784a2ac61d17761fb3816857598f5820ae408ed36adc1fc99139e85888fb0d45f7e7d6d2320d109ecd56cb436370a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf1a4024b4bc9e531d8149f87a856bccf9bbafb00252350bce9ac36c3dc8c425ff1d72623b88c1ba52fea96649a77ab06716772e42b438e063ad197e35b062f7d49d1920e7efa370a7f72a497735f118ae9de5963d460733ebe868190d07f2bb4247;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0931f022b306de077d4634094b5183342da669512d88620383aae6f1f43dd6e4f1d70d1ce5ebd7e61f7d20ed05778c62a9a7a080cd1fcfb3f4c94fa295fa11f313d3be0a26715e0bd4445f888c0a8685fd969323324b06aa649d4310d7f393755c1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc87028b5d393ef973533019d097c22df447603ce803329cd5d55665d0ebdf2a73d58f1f9487869e4af86214e3a2c516e0862c4c1602c696c953808beba25bb077637f88a73e26edaf57aed38d050f3f06eb7d64f28e83aa81d6c5b9d0b42a20d0101;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c394db50071ac0776186613960f6ac6efa576759f65e1e67ccde3f29cd8a642b86eedd74240544ac097ea54bd1ed957881f6e1209ff817530869b5c8b9411aea3b6cfd602e4d314b8076655e0119afb90a88005d3fedf3521b48ca858607acb19cc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1a4e214e36adc1b488bca83babe33dcdf0b59a4f3ffc274632c3f748a5fef24d0378764610abcbed8347ee0d7167f6b62f3c9fbbf8702edc574c60f753156e41a2901ab402ffdc755370383701339f5e47fd277a9be9badbb0efc01765eaf8d9a006;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9bb96666baf4d2e5ee341303e4267f9218dad618ef72879bafd987c58799d4dc999843cb5ffde17cb8c418e119a3aa2d77a8ae77027d2b862007707045c1bf904491a1302cd995b8101bcbcf0c7bbce025b8a5207a4feb1fb6109b1d0d469800f84e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49516be1ad04ac239a34fa2de56083f1ad3bc1d495fcec974bc9ebee5b80a112e62711ac729fd52dda6331d658ed6c0fdc70c1a3939b9ab5c50027ecaa213b2127d20200fbceaadfbc8616a1ccd5839517600f0cb3a89f16852d9b49d51d7b9a8ea1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63bcff1a75e0f674e5d563b1c958a71e265259d7274a1994077480a38104cc3f28e137e9cb379182a6203e3d77143971a60280d6356829348277c621af3da5b81f1e825f952207fc69408494955fde7cf3e35493a751c491372f1a7677d4504dfb37;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdbe9f55afc920d51632f2595a2f96380002e070f5a8b8f180beff3acfe16c21cd90cda9579fb9bedefd041e4b50ed2d8be0edd305495b9bca5aa5ac33ea3506afaa7f04bc1e66090fe01bd14ee952c015c774b2de97fabbd7bc550c38dd1e67eb0e6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72410faf0cf734227a10807d2098f5ca8198487b7e640d05f2f3ad549ecc96a9d00859062afab447964e13bf6dfc05d8eafc5caaa061e261f40c34bf0605cfb0c0d33a338a4f04f939621e2d9655e9180deaca3f47f19d3b76520c641dd9b8248c06;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee17c20b9e6c7ee629c8743e54c539060afce8d0e8a6d78b5629d7e199ccc13229e072c3441cb97727d5dbf7b07c7f2c3af136b7b31928ac2194b5e227274e90eda72b052b796384049cf08de63d0f304b38c07353ea17132725ba93921fd21f3497;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d943d5d8808d2bf7a548249a7f624749c32d8a691e649c6cde7a7ba43820af9e6333858b4541a6d72d28ef621637e71097a866f2ad4fe83ac756129840c82312aeee51a9feef20cab96ce7eadda3dda5bcd66acf47168135a55d0176c7c98b54c28;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2685f6ba76b566734dba621650ed1eabd052dd391ffc8b8b2cc0f5f7519f7ad279e09467aea2e221ba3fa43a51fc9a651b6bc9f2a554576b7717461bc90bfcc2272fcde9dd3de73bf0e08a809725c0e116d314b37f1ebb7d2467aa094c6781faed7f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h712071d7b6097328b4753c40fa1eb68e2deb9a912078f7a387802fb339bd6957c34c12abe6b4b4f81770c5ad6640db1b47b3106c83864a6695a033ad6beb1877893b04975ccef1dfb82721cebbea689a394da47b2256111d80f87352f86f6276c44a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h832a504a3994b0d6282bd2447293db490d7fb95831f4eec28cb0475bd5934021cb0ec23cf7f02bb4ccc4d725a67e53e30271a2a2b1a141ac248833f4609e1edf761bf7554732eac608695d80319109e4027b3050e6c2e6f724dad219e99a8cf373ea;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf24db118e646ab0f423298ec343e5f5fa2988a7edb44c4dc10793f8db52deea7d974f25512c756a2082f85785ff9db5ba0bbf9dfac5f914f1ee67c16fd2086b0a41dfa32c46f63fb331ae7c54cce7f8cb13766fa43c7f7033827876ca10926ed5be3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c27d0ac6acb7fada693f15ecd3d39e02971462fba6cf96dbc685ac0d490df9554a2a82a3837c55787159a81eb20038d32040c80f85236808f8e698dcdc7bfcf991eb6277384a09897cde66d247a7d2610803011f7e99b9e17ec940ac260cff656c3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he578d9efdcd3ca6ba0b938da396294a37e2e7684c55e1e259290e03faf0a6e8e37557c7892d430ce452d1b1b8cc18fc186d7dfe290963983b99d7c4b5c4c2df61556d987693e672b513272edf16776a1b27cc4db86276d26bb9622de8165e600951e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2964ebd5deba71585fe467568d3725d98c799433f31b40362d40afd8bae8fcafb350e6cb7c16fd61b27f6de909f4d16973321f6849618194fa2fc4127b7b113c03d458cb1c17ebf1d8d9a16fd07b2cbb5e8cffe60ccf70c4fe33af4fc44f3c6ad4a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h907a7dc29de007efc6f83099555029818c00872a28a0d9db84b5c4b96cbbca414cc0cda0c94323fb235844ff15faa594e53ba0ecccb8def99dab4e9486cbb36324406657ca4e866bd90d0df6845e8fcf10a71d1d12d1bc903372471c5c782b3ad1d1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddd92efaf40e3a8e369002c52758bbf73c487adb5b3e1e38343bd9f93785c320477329b5964dac363603d2e524e9f682d16271e1e2c396ad08e6aa348037ab7c74f44d1487441c6a35774374f27e93748c8195250214112f987969e85f48ceece843;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc32e38259fce4041f1aff10b609ef37c97f1d81e083045aa6296b41e7bcf489cb080fa565497df1c5a578af274fca7c06cde1bfcf72a68892d5b69cb915829268342dab65280e975cb5b11a9351c9c6b6ffe8d64d1fcc97ba0ccf988ffc7bba47d30;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b903485c3ee5831b966f4cce2a8bbef52e556e9cd59b3ad8405233954415a10f3787703bd6ca66262848316db81979094b4817cdc05d564592785210b19ecc839d4cb0cbea0e3cde9b86906edcce0210e994440b60964098d76a68a7afc4069083f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca6faed2ab3bdf5de385db894107dbe265c2ed5f1a26e078547a010b49c31ca42d220b149ea0cb9733191f049c4950598a88a16896d9106ba4027cde4c0c00acecb47ae7457f17e97f1666c62ef540364fe7430b35df4e762b3d6b5f8674e918be1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e495a8c63cc1b1f68b3552ac56cfd113412f7dfe0705077a656bb8ce6b2dfab0fcc946baceba4beda348c12808ab7b1b4a5eb453fd23017309d025f24c54441aebc248e97252a17e592642d13713b89eb574f03f5d87ce2110f7c20bfdfd286e1e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ecef3789d117a9872c082cc35fc888c8e85cc602367b2299c64ff86a498b88ec118ef8cdf82f87bb6762560c400a3fc55e391c7d0c6ab65fa484b3fdb54611340a0adff47c3e1d6e0bcff813d12239be537b12d2a36a67c5693c6435f9c79e7e1e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35469cef004c61ce6b8893855b9b8cd526132410b6b114dae524cbb4e036e5840e295c7c1ae742abe667f40945ca0ddcf895fe38b45dbcfd91047170aeacafeeaf924ca01a110c4ab770566cf494f48ad7ee02c9da95e22b35afdda4b7cfbeb534f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf32baa5068e4840cb6383fa51f342ee92f82ecff89fe4bd7e72d1be1c573238653806ecc98d6b802c2d515dc0da25b5b760feb280687cf5721801da858ce3642f3070fc007fd1af9be3cd56eb13ebfddb8e2e67ea2042f6bafc3cd20c65b62e646e1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96a756afdccc83870d3ffa990d3df6b8b8e65927d55d6d96afd41477f4d4bd2bd510c1c77af5aada9ceb2225a83cbd08b26a60a777bb7b427fcbb9e9db861b30ff02e8bc57ebd049f714cad890de84e73a7cb12dd802e53d0b4558c3c20c9731eaec;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcae084e3f305d7c1b2c03e6bccebd60b0e6ecde0479e4fa9d1caa21d349288d115fbf6805e562f9d21c4c8f14908c332855e810aa5254bea498e23daf0386dd521b19c377731c190bbddc048fae2f652e51c598c4dadf5e17af18196c8ead4c00d55;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb676223cdda36f3e7c68df9c91ea015d9d2e6bbc557d2d4f96acc4d42f9808435a42b617422ac2d6d42387d018751e0a52610042d7213039276dbc95bf638c233384b9c6efa7cc9257aefd6b09326eb4526ddad8f0e0d4a2e261700b2ca3ccfd8ee2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e54d2f257ae0e903b6e4a8bb7132bb0aac17f29293d866e093e4787cbfe97c824fe001bb48aff474a224037dd5744cb1d0e71eac51e24e5771dc461c16506d8f1a3783ecdf15c2c9761aae63f6477fa6b9bd43c16acdb40ea6558272d9d076f8ba0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c697ccfcb9abc1dbdb7452b929babc1f798375d8b8c7bf9cd8b2b2ffb69924e3f246ddb7b5ce6e5cb4a4fd1e162f31cac9840adc1cebb11f839c90637a9eef0cd64c90635c87a8712c388edbf6564f113883d670d345ab7787b70ab8b1a994b193;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h474599b3d5571fc0a735dd8c85145a38e4773bc00c18ac184d9a384daf2158a4689035fe7f3fc9d6f0faeb6dace504adc0112d3bbae1935658f03a99ad072dd5672a0c04b02c5a391c9a42a1f46fe8455dee85eb652d8e555ade9d4ba6fba449f7a5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80c90c676ffbf313a7d562861401d12125632e7d4ac6548ec675d3d3104b795171327fb2332450b61adf7a0d648784580d1d7d7739d2e0dbdc38d690dc2b8bc9e120234d8031891eb037b2e4c53c42f602e09b55b06c3fec9518a7d126de38b21bf3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddd08e0afb99b2c898fdd6866f546456ba66c2f8d960046af73a7223872f021cf7188c9fbc87e8f364f24531e7e506216d3d062b8848c39bd1e2e0008701cb247adb7e7f3ce033c86e89c6ae8aa2eddecfc692876a094f5725d4ddee2be3258f736d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd113abf6c382384e190d8cc630ccbb5c40935e5361a1b91d05f9cdc75dbdbfc05b7fad71dd3c315a50b1fb5edeb2c3a98ea44c6013d3ce1fccf96dc0830e2672f1eb3bc5a415f207ace8b005d17148bad6ea45537f34fdfcb430b22946aaf20a385c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha531ee0b17ff4559ed73a086047a873fbe1d7c8b44283e93969e13203eba628f155490ab434cb82725fb87ed58221736b66507d5ae3611952776f9bc286d2dde865f982ca651eb41f72da3ead9ebf20d41afb86ec0ee0ea0eb2fcfc9ee81ce9840a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc79aa47752eff70cb54363363ed811ae6484d4878318e18cabadaa6c44ce69776c4e75de6a3960879c5d36f95acd9834ac96f43f21d7b88456fc5f8e1db15cb879d5c01a37dbcd1f565831691b8eddb9bc074a6f32ad2ed89f8b2e5cf575c4e5963;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2ececa8f9f96ac554afd147d528e2e379163595462dd202fd0bf006a4cc58b4ef99f6bb603f6249ef9d1758bf8f75988e48ad7e203379a66ac2c44c7eef7291242079eaf9d30df333ef5cb71663d6e04232191cf72a415ae445cc90a93b0d46dab;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0393537be48381d5b6c0670c496c7c19f2883e2bbd7c83b1fd97a80ad2848f62a027bfe8bfe558063b8a11656e1f666b82a65b9b5cb8547797b8116bf501e30679c96a34ae000c72a51dfee00c5299367972a25e0180d265a1d2348ba0551300afd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbc7f993d9ed18a8b388a1b7ff5a3028feb8edc74beb0eb82a71f77fc7cfa7ea59433c1672cb734b35e23f0b6e66c9ddb808e0865c6f842cb8bd343b647c605b48e8d66ef0a098be02304ab4c0ad19922627b2a32d00a3ed02c844c0181ca413c196;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42daf7408a4baeb04c3223a20d2641991cbdc80e36ee1f5e70c9006e77554550b1c901f95717c65f46bedb70165c153d6a081642b1f25f8f18a61fa3ad15dfa06add13c211b1357c341d1672657e2149258c7de8c3758f7bab725657d733a05ffdca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb6fe7c4a3d4514176e88a48f9a93945b7ed6ba418d3e4fe643cad26873cf43688d27ccb28c6eb9d5901404940de0feaee1ede52bb576e1ad78bfff7c1a2fb70d6a77aa2b00686a91aff3a8101ae9ba22affc24161e4abf00f3bc82f915dd43d900e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a74881e3c3c58f6e65b797f37494c903fce335b903230f5fbb465eac4847321b2757d2c99405d29da6e93770b399c5d502067befe520a2925aa5e3ecfd8ca6b0251a45f881209556f13ad9930972ca89962d7ff16af5650b04ae525867ba483cf94;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2f11637d4a5f516012c2accadfb4602ba4b51b59315857c5c13903f05146f03db0ce7fbe1d109bead434bf3c4d424948c923586a84ce06c645f138763acd2d56f973133069ddd29fd56709dd5cddcaf909740eb70b97363cfc4ab8c748eed57b25d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h726218d3ac76a23f60f67495cb692bb06d8d8f0eb759a1576e0fda2a4baf614e0b2d659919dba52e3b08cb7c909f3725b280b5eb4a9460fe813e4e0ad013ef11745998d567ee5ae5f4d3ffdd0d26e8497530ca49c7798b82beed8ebc0872c76df8eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3db5c56cfab38863f51851fd60e59cf020875066b9c0c42a188dfcf1677e63e422e6754a35efe2af152be69011abd58075b73e15f115cf942ef97c1d069cf71232a817f53ce82e770ffc9376b3cb55d6f233a9becd6f754ead1ba125071eeb050634;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde916adea5c575dc31eadded7b5b974339295b0d84fec287bd45ee5db8d83445dc61e9354b97be6e7ed322971b170f82470bf42b64e3ef1808a02f0daae3ea00b2408d487c70681ac218b40a1d7255db90271cbaf84c71b36ae06e18cfda64ede00a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h790b7033c5e3b8020f07e08b2d6fc18d72e9a1c20aa8c95436a5d702b534db65dc6c4f8fc0c9cab2553664fa6a4e0d903735265ab7306373d62b7137e6b4f43d9dd6702385461d9ec10b6c6bf2130cb6945d3242bbb249b4ebc8ff95bc04b939b40e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72a4ffb84e292e7ff4701d28eacd2431086d2ecf1cd76a5afd2e6803c4cdae0694cdc6531b0e1e75219055de0f18e48d7c31379ddcc8f409b99840ef832c2c857c3fa3ec777dd8cd70bfabe2cbf856845f78cde8cc7e2eb8975a901e04961d70684a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37e2ee146c224f46ed4866130116da06eaacf097ee55fa389eb52e03ff77ab2c4deebc1e7875c340198197eece6d405861cd342752ca952f563df8bd7bc9faa37decc27d988c5110bc585c1cf98fdbc92908e4254eac13898483cc286b09b5db0809;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6983ac2b2560c21ab1b36ba4268a4925ae77062cb2af49065bc88339289250bc8154e5a5bab5c418837e584754b19db0489a65f9d7769fe764e94c7b9828d179eeb990c050ee86dd0a37a1ccbb0d89f8a4ebc8cf0c3973de4e11b882b1cbf48feb8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb0c3eb1157247a2937fd7a51c4009b83d1a16cd5ae766ee1e69d6f9a2e0e9b1ece86e1093962ba2b9849d29bfac71b32cb4ef7db4b37f5269e9d596e613ac97822ad8e9ef8b85cc3d82edcf61657db5a211ac8d91fcd5737b216a60ee6c5e4671c6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h266cbce021fd056c37e366678fe335d85817680a6df06501e61d671151eee51126eba749f46af163ea4095374aaf48d373616a93d9c06c4806d8119e8b721f581846262fb5202dfb3aedb3eb211cd1db9ca746ee647040de56395511cdbcaeed37f1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbf62ce900aa35a04a6fb41652f74e3d90fadfa47774c68bf99a1e119bc1647e00d019c07b4a9be120b9e4d45a4a597ed72c838bd7fe4b1a605d9362a9f2c0df7f1a4e169037204d9edee247ac734d972470d3b09d55f5b7cd5f9ff9c724d7a55a51;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72e219b7f32fb7feeca9977c0c292371cabc17f2db7a39ca5fae150e3b52597452b7a6d6ce0a731d233cdb0428d1d52b95efce27d58d2a12443c04b621f3064298397d098ae89496ca1ab988c63daba3921598a356f6a8a4f63c310b1475dfee16eb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca2b7bfa77667ef724b1629341a2eca16d76da861c85f25f6b0b1700f7029ccf2221fd78fdbcb92505497cdf613a56b6ea3d6d6129127e00eb7c406a86f8fa7b1832faf399a0c929e14b19c8f6c1234774976fcf5ac796ad256e57fda0d07e76e66;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he101747dba8845d189505e25542db142f766f0fd0e6aa179a3ad8ee46f94c43188bfed83e87892ff843d2de2e540c622eefe0f42beea0ce676a1602eba443188da9c5ce11b4aa1856b14764ed33b2dda47824578f5bc81f4f92d3094c8177bd1238e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee68785d3f882b1e445a870c6ddd37f7baabe078ac75385ff9a153a79322e9b9695797ee696f4437d825efe95ae39b17cfad04235a04a9fc1fce68f7234eda3db5e7bd6d1f59ff7091c191b280541afa6135730883c538067da40541d4accae7a6cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5255c7ead217b23a3b96be3d097938cb53531dde850c091493faa6baa4bf60683c695dcfe9a6aac6bd6c7c98873c72eec6aefbc2b29b01ff548a1f92bdbf7a8e55427f612de62029e408288b3a066f4de4d8a7e71d68f61ad103622fc2cc6fe10e61;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f98be2cbc7d0b4c75b089240d3f3967501f59e95e19f5c8cd6a7ff546d6e01a1855e90128cf1455d21c9749a99b1cdfca250e0005116bca3b9a8b0f7520f630ee98969982f0df9d60b6e417520a3b7db3eae314064a7550ebcba05c3d3c806f1721;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h374ba26a8598b8abe80d889990a47f12b8a349bfd1955ed4cf6fb98850a317dbb132a0ecc530f39bb8084b4b90aa70650d2e684ff83e2d0d3a26df7abb8a09171e2a844dff48c71471fbed42218f72b12591a2b18a71efa18069237809491bc1c888;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha20e96db05abe0989c1ddb073e79fddec474c5d0ba450e0c025f200521086ecac62774149905d0a52ac07044d78d2b77a78bc3f15914a56d891abcab36c877310c4a688b86ccca15b5fb868f715a1b67e7e0676dd0bb21ed77a1084d576e0931bd4b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3ce31c781fea033473abae5f1d795e0546a28dbcc7ad0e372bd6bf88b9656dc4f828dfae30530fe629f4e209a6c804fedfb6c031540ba60a5abc79ba2767cc3d0ffc8c59f2b8f6ee756e4c07f6c9bb6b559eaa9b55f248246d3a88e8985a61fcfcf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0c67fba97bce1793c00ed05819426095d8d47403b2a722888ee7e9ab49898494e1d6372927326f52b79272dc6885a1d8b9efa2acb02da61e02ecf6ed84133a0bbce07bd7a11b9151b6f9b20481c895e346b21ca114f112bf38079c4f07e1bd62e36;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97fad12b4145191cc580a04bd59a58801508b31860a34326340a5681dc0f9951f291dfa5edb700a69ddb8d9bd0f87cff1ac9b19e525a5dab1072d2941b368897f1f347ac3a53266a1ca142ea5024c3f5c91470aa027a5ff66f41ad3b7727f19c7f03;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4bb076e31109d388ea4b31be941109f1f648768118a4d4c0202a2f7eb6822ba0eb1b2c40aa52d3ebcfc1e89c0ef6b743d10c7ce0d8a8c20c5df923d21050e863ef78b897c2317d5c35ffc305a3b37d167ca700f08f21d718508c53678604bee05f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c9799a61f34cca2adf9733be57d7271d7c8150984ba1a9fb14ac8353fa15fe0b718f6eccc1c99f1b7d933ff90c68b4814b90060058edece737d7b879dc32369f4aaef14dc876ebd7a1403722ab6596647c3fc0d470ec852cf769cc5c2a2a35ffc5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45a138eff7f85cb6ca9b97d0adeb6c80f869fa533682dc8594c2f5ce786deb8f92aaea1dd0aeea5688ac41cca30b0777bf6536b3ae7ab5d865fd08aea80570b63da29eb3f02276c1063e93309d1dffd1f2963493114ac54cb6d4815eea1543969ca6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf04ac062c4937d648687288974d856ac0dce3bafdb7547a9884a6413c874504bc13bb01f6628db2cf19eca205f2f88ebd2eda47a32d74b148804ef563d02331d70a98688cec1a2071fd92cbd62f03950e21cff578ded4288ce2d7abbe1b142830f00;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h938f12a6c002a2194c67020fc6897e44ae5347be7641825d21c026bebb21d11cccbc9f333d0d3f00d2bd89c4fa32d556c7bb1d6b4006f865882b46d08561c82b75569cfa54521a880ca257c8d7cf3b9ae612a9f3d7c6aa056a85790657fe51cf57a2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23658f26f137c52048fb6fbbccebccb9e8c6486ec29751317ffaf761ca8a943a02d595c6c8fab87d9dff025a1f3419101b1549db642836e7279c5e31c7cedec060e9901f233e663ca74afba8660164d2cd36630867dfbf854d2e01274e33fbce1137;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5267461e51d91953117d0b3891be2013df74e7e0122fe860184445f3a118a1d8b79ec2e9cfafa76395b8189cdd44e964d87588134ea3a73e7b0d2af1b210cbdd6371a2aba6cccf16b7e10bf4ff9dee7c1dca09b2129c5ae438553d333ca76c2581e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2eedde96da6e0a051d1e6bc4b7a661c87fc0ccc365ed4b3978a8408483c7cfe9074da9b4c8ef76b1e9fa5277e227f1a9b0b6799d12d9a206595e568039109c98afe0e89d8988ccd0e6579b8bbe99b1a35e75a6fba190ea821f57ed786888b6d3ee7e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef4554a69739da5076e86f87b5ffd78af9060a0856d0f219cdb2bbe289d6c52c95f5f45e1abd67c869f6958dc236736fee29532e508cfd5149c892779abf7debe1da762d7c07e8c6f0df4817c7219b5a1c9f53824a167d721bca47707520823ba74b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c5f3c6b72bf30681ac3db94deff6ecc4ce2505465d9a224caa01932da3bd56b88ec1f11c2c020c4410d9ec6a18c80741061c76f07e700fc35bbd4d92ba6c16bf0886c65fdbb61e869388156590a54fd822a0ceae535e7555d953fd7cf75903d6e60;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a6a185fe6b63de26421de965267149ec5058f547cdbb8a0c1fb3c8f1e3939d91d317f4af4b41de231a3b6f919e03908661a2b830f25fd9ceb15f95a20d267b247495a0fba1993accce38d96ab8f32e2f0480ed4f9f39ed994aed24b3bf70ba1d867;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf3518003c99ce2cf231e6437561d5a12fbf5d3ee8273a5a0be8ab8da159f61d1db137a14d1f70d81edc2fb05644e68c6c7fd5cf8b93514555af12489646d5d04f459657119a6dd8f63bd28956acabf205aeff4e42a211495c5559b093fe5ed24e93;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1dd11f89af78c441ae3b7edf8b37194266a3cbcb7e862d13c9d25ed42de0f5fbd8f9f949d3c05360937982eb4c43218f9f93911a8804bf4e9d17d21446206cfb624189a020fccc6a97af57d522aa1b7001ae0b5ecdd6da4570a678c3cf870cdd4a25;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h327bb533840d665d7c0d63204af7afb786b13795bc4e513a9d98435c05dc21714d8220af8ca5e9a86b6116c5859783c2de9c409d436662cff1f0f14e8f16554434150f7ff4c1a7ff13a05dd19b989dd62a8dc08987c22809d5c7d39377e176aaf68a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ab3ea3877b4b6572f8f2d62b66bed3b7bfcde3f97dce5741b428541216f070b37f4e4a31b3fa2da4a597cc821784708101fdbb0999fb6a0334a16e7ace0463a0ba2543465033196c435bf6d1e81956b181d583bced42975bb267ba9a4057abf67f6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55c93de66aadf5901a244489e67eb1474f92de3a20f7f96464d19689c443106210dcd0bb3abdc48cfb96b63f9f4ca07019a9dbcf941faee87347451377f5a83e1a2d133a61211e8385c02094c6fdb869d05a89c7ae304b1b55bc4366d00395860901;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf83f4c93a1e8ad679a0290fb438e34c82ac3f8d67aab5ce0f274e32175b1a2e1efcc2af4b85b4784cbe13c5f08e583bd3d6ff3ce8d7d098927b929302c2bbfa431f851ec8075882ec7b65c8ca0887e1665d20b6ddb64012b1e161f0ff1124ef93a23;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hebfb1f411aa0152c582c7c00204181e9168f164df9084b3163a2f71746a696fda630e2af6999a98a51750ea0a23b9ad938d857a7a1ba3eb5b4b7bad36c0f8405a122472ce1c74133933ef63983e50308d50989156363e788c7216cdd3aaaa5aae5f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79571df53959b61b7cd5364b676091b2d37c83fd0dcf2fe5acedeacbffe251ba574c75e6339796b59f643b136cbfce5ed767a5cf10ecfaa030a0c250c76a4f929d27c76d31e1bba692788f19d13136342e46ec63960f9f01fb4342718adf19729d97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he463c3e51457173e496a67292cc518b7fece30387b9836c8358c069f874841fc2f9b3bb4566f590b13eea3b265683728d85ed3bc70f3cb8fdf8acb96818d979e23d7a4798e806a37d660c322bcfc9a2fc626c10c36255a912403528e1d34a436c9b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab7946ae8c79280198021b41094f8c06ed381163879a26460ad565266158761cdbb8b075a6ef4c85902892740739dc84ea60621b1b85aa0d084deaa3170234814d193db4fdd5a12167f16e15cc2ed8fa48e93617830ca62d36f6402e56404dfdc5b8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2494e5427da74abe288f55b16880e858caae417612398c181fa3651298c9fcf700e3c7262e84373f898e756bf7df0f4f48d0f10cd35ad65c45424a8d54ab434a9062356e49e061e110961abc3f117bca89c12fa7876d0bcc67e9ddf1dd0eee2bd7b2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f094937e69d67cc6d3476e95d185ec851dafbbb58d59ba7a9138545237c7973b6f5d54e3598694ec8988e149c71f475f6f31a2f9dbc7f03d2b1381fc8ba9a3bca93df33e91d15fbecc7656ce124e3023a9374daa1cea3805b91e16fcb876655dce6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd87b7a02be2ed7c16b3249bb2135b3a75a0dce2c9a2c0a235d9a997f68ce84fa23737e7969a23ace3fe622da57eceb77503ce4e0c8b40642d83f508b5bb38915291a11d03a8126bf421623271883003aefec8d4a3eb2ed5f56e6f66b0d201ae554f2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h890c49dfea27c9cf7d0d358807a967b488bbacc66ac3999d7da6d3fc6533d5b40123a0963ff4ff753c0e26c3d6e238f49030d9d3b9d06e96a873eb9ebc04446124c45537722c8b138b262f5dd648e2df5756df31e7e8be2c21813777950463a26452;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h762037272a6ed645bb5f61b73e5705bd47ebdd9332f0af6749e924b83902dcb64c361ac79b4e255d2dea871f9f413fdb0d2714be7a2ea8a04d51c2b01903a33d40d7fabb1c62f9587cb5a23c83cc8824cfba521daf299a952604a264d6c13f25fb99;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bf02d4d00d985facc190936f46dd472c0eb179b95be2c4f88971b772a128d72e9e72976f5c10c837bfc479861ace8924374eb98ff56c3e0277b25321e7f249a39222ed0bcf2bfffbf780036e358bf3f0c038768134123556cf535331c3af9527d7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49c3213c997772bd10a5a428bd8ef791943cd0f47cc857065344132ae5be1ba373a3619a4f36bfd9518608b18c818ea4a912537bacde4f3ab07c2992afe9be5e41fcea7d94b0ba70bfc32f3d60690682dcf892f7c79fd9b48794023a3dcc3e47a3cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9383265b3136825b01fb829817274b8698535cec91be6c697b12c00ab0dfc893eb40f068eab8995328028d57240e640922719e648b7ba611688bc8aa75f9312c11d607f6f785579ac183ee4cd0d29c5b2a78b4b7654480a90e09e36a948e3ae27279;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had4987d4aae3fb42a6c77107110601618907013d9f480a11562eddf3d1556b841adf732429d6c0aa8da4dcf9f03cfd417bf3b6177ece88474f78b6091fdecfad297a2e313324210e734a1a97700397e035ef28071084872fdc35f13e4bfadd29f285;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb98e3f51cdf318bab1f7346d4f64233667947257205d5b319796386dee324bda654684b6f3093c686300beb088f33ff4cdc56dda81f26ec497f2282e39e5e3d1891d9ec6143d2d0a1e020869ce34e71af63f51aec2a1ca1b5dd1e712530472a48685;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h164e8e71baf3eea96d2730cd4e4d75a73cf935c193f28b7a6dad26d936fcf052c0a468430c26bd5b16e5d79a1c27f66ee7b18867c217e3bfd02413c5ce4bf21b4f5bcc09275957fbe8dc3e79df079b74ff4c7928b37ee62322f8674c8ebfb8d3591c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1b79a33877c720d4543c1df77ca9219b3cdacad2a07d299437e62ef91cf0009d2b88f3051b91d2945914a3a6acc473c50fc0f4f1aa9656e10ec325d3443235cb59b36093b633016e3a103d9f6d99a40e9eb6e35d96f834916c55344ec5924a4f7e3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64d042539935f6a54b0892b7b9753de5926291beb161efe3741434b242ee638a6f8a8f0616a79dbac879d28336921d0f01a36c92e3e30d54c0748ec7c1be5922407b1bb91f697e7392adfe97bf203dcec4fb454c2707994e54ed66e13e5814883ada;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a69dc0f78171a2879db4a150212b33745e5765ec1fabcfec9d38b902edecf137e51ee115f3efc0c6d6199f3712084de78557e7800f9c58762847af631cad057323d3829e3349cc7a8b7ffd22e49bb638fbae0bb70c19598188253b083bb97718f2c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19906eddfe3d47db69bb449276570978728e8c5b2702fe783663c044fd20ed041f1e41f332e58f7e7f25d184a0ff79abceb0fa1bbf51ebb8bec8e43d4d588da028e056094d14cd32010557c9160d73564e5d649e3e6fa04c1eb2db5dafc0f4db408;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcceb1e31176544f77e439407114477ce012075a1d1bed5ac65d5459629a6226f7210c82c3cb1ec4d69d6539f5428abc679748469b5442189b54549cc84d6e0ce4e9757dd5ffbf86e7097433f4699a3c3b965b341108852a451e949c1d7c0e498624b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h459c881909a6dc977402c9286067c0967996f0ca7a9ba564771861edd1cc86d2cd21291cbb880f2a5b13eddb547b3ef04ab99f7e04c326f8437500a77ec76152166e4050ba5584a2b89ec83b82383be01ffc3f4a2066c06b9828e3c8bb7dddb332d5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb4780e99cfd32662ee38dddba2fcc1dfe179ca140d43b2d5f4701ef482706622527f452afadf2838dd1293d2952cdc5ed31d274a64b2c1a62eddec3d343df52cf28b57d2cd4fc931a38c74acde836c472ae5acd4a90eff903773d852f9fb8c14b96;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8aafb58494319f014f544ac5fbe9db5357bd41680b093bcd256f73f7819f9b4cb2516090104350f7f5cba1d5d3b98ddd3d9ef6343da59b88e723b29f0296900d03295dd5e463461bde69ed995f6735f7742c462e10b3b9ab468673c9a7a31e8fd0d5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd931788b6f1f1907abe2c680f1fae75748fd1e590458472187bcc2a469d6eb9dd464381887b368f09fe9383d0acf3ebb3500f76665e8597ef949e34d48a6de1f65cdf46d4b98dbce707169b41386ca104c809862846c31c855f3e102fa57d42523e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e51915d92dd32d114c5877b851381eea66388c1fb9ce2e5dae2e58b9c4d3da89b371aebb0597ef8594ba0e1d6e9f3e675e2048adc51252811974c403399906391d51798f9260434169ab2c7b79eb643fce022f22c70b6c648550d9da98412af81a9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h464d37aff74f0b49c8e35bb308a1ee01b6ec6d2a68c1d8897cb146054aae0674aa49e2e5821e7612d350797e5dba2bfad6b85493083ff51f5cab8f1cf271eccb573562cc98aa9641552953e9cbe95d713107f300cee96710b256600b5ef213e09193;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c93c32b95f0c80dab04216f24cb01df60030798110f03dabda9aa8ba0fada019d001ac422a9337c24f572c7570dbadedec7a9642f8f3cb05c37232d58e74d612c051ea2dc9bb5cb0a7e9eda48d8ad84308715122ec28b41a8de0b4ac664ea87ace9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2a87cc1681c0ac755492bce26c0688656bc631aa92f6a7d121a7934c347acd2b6e76ca6843106adb9eb11081a4859cb051986a8c1b5167081614a14651c58e479975a408bb715cbd4101b61ab1e39bf88d444ae2c546f0e168453c5b338a492c4ea;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h543b7d2ce05fceabb3047816d05b0bcaee6d80c063d636690b1cde9db36145dc22423d1596179475693a37d7c60a3dd08b9330f6ab265d6d3c33b76e995de2b921fbb75a9823adbbc0ccf99770ab0108b8fc0958cc128c1c39516ffa165f4334b23f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbdbbd0a38a983dd7449e256a81fd11a6ee387de129e55d8c107170228786a22627d26c086c4e2493c500e706898e152a18c81d9a8834ce28ab02292b731de86149493269596b92a83eada82f07efc3679e9018c82f1dc86247e7c92edb12eedfd403;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e885eb84adc7f0104bad1a8b4b7c47e667f9d86d3122f08baeb2b53fd276750e16878798c4af61b70731a04288a2d30353c841bc08d55a497fff964ef8c8a74b2c247a2e9dd024a09267def90fb9e4a7e933100765da574e7d688a88319364d30b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3ea860f6bd49c383ba0ae158ea134044e87224ffd3babf369a1383aa4ffe71513b609c8b1253b72b7b329b2a8d584704ade815731d1c5a430c7df3fd8adc1b99c1e284dfb2a50ab02a9818da1b4b4bcdf60256c7528c5b1f96a72e4f104d46b051f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2706b646d68e5359f59678f874884eebda7048c1162b120d7889e690922fad1befa9c87c1b54a2cde62abf4cc4963d283f8852fe06c182fdf43c6d633067f1c63be1d051149a697e6fdd1b36a20a8957799071498ecd0c27b4f3c4979578d272e0d9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hedc1cd327f12c0b33e33b56ce22f6637139b6b0cc58659e3aefb6a82f4c8fdfc9ee8e8e81db1161dac46691692ed7aa3b044d927da136388b9659768c3bc552f41a64dffe54e5129d4bddd4c30ebd7eeeb8eac77d3c41fe5478115b45a4cf3155dc8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f8b884f750dfa338dc5f62cf0b860efba4f910ba9806314ec5adf011f80908a755889192cf527bba33dddb33e350800f263ef53ae2e2256e5fad0074b2f2294d17f8cabcf56f218e045e79e5421032bd136820691f4ee57df51ffaedaf0c2fa53ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ba841735fa82567894eb99ac51a5d2b8112b27617bfe807fdae897df933ead5d31626172ffb5dd46036e2818a01d39e211430552ced65a5fd0c8b7b7f3b357c27f83bf6984123217d9421c8481f3d2311c99b7d888faa3dd89ae8bfb63d10ce6d03;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1a30e3aac5fbea41913a6b127c1d31a12aa82919c3a4dd9ab40473cf207886c5e990c11cfa32b0ecb26b0752b61de72dd415e5113de651b203213e6e7b9268fd3475012509ee59b95c62ba238fbb2c6aabc20e3949b5b61472c638c3b7432721a1c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3851a941a0d27c630d4d8672b33c1702169b5dc28481d47499835056184a4fc3b49f943127a41a07a476be653029d2576cf1622cec04f34be90c548e3d249b1cbb322247214876ad11aea8ac5b4833efba7448771038de17e55f70f87d96a2a02fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h28d07858433507cdc37bf1a713cbfdbeae8acbff47972650eca170a342ca768e7a5c9dd81ba1a1498f17885a6597ff03fde9655d3da266c13229ed2d6c13b7f7cf7bc36b29ba04770f6eabf78b7fac630644decc03fada18e7a0f15c405b7cf02c96;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59f6ece08de567bdd7701d1bb3a99b952f4a07cb13dbd85988c6ce5e6765d230fd5f9d6c3799186f1cbc20a7c717356afc2fad004909c26b910eb2805213ca95b2a36df62ee03d90a4b4bb3a9711c93bffa7df06f0152a31e36f0f3ed966c131f5d5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ad9e1e0357ac93ef8fb4beaf806555c67002c6ec038f9c65f8807427589d8e5fed5216e670a06de24ebda51b0bcbddad8b1277c6360a78f7ec644ab5cfad8de0b43bcecabeedd7d15ddc138829f72fedcc302272c74b2f94516274e958c78ec7c08;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac4db4e3eb2969da578aaac1a31136605e0bbaf9334587cb01244c6e7b021440c84276d03f5dcd018635f5c72f8d5b64512769cb788a9fa69041243dc0602b3d49d652c17890ce15c7782d21e77ab3663f053dfb3aa2887af18be7d2ed5022cdc5a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc51726696f146f8fc00d90b7377341326199402d061b95eeb1b797ecd8fdc1123c6ec461e5138be4bbe11df3433bc5e273ae8c90f47bf55b5b36fd4e339156ca7bcfef8546128c758f8e1b00e0b6cef1ce0b16889f0435f6b6239e0025113ad3c6f3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had12abe67e6bc439b21f011af4893edf13a8fadf50ff9973ba4d50c91a12fb5cf8f139c37b33584627268883c625c1f0c00111991681a15f4627ec0c397a361db754ca6034bd2d1d7598f05d2c9b8cf03764c7ac849e58f654971c1b6656cb026883;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8330fc42d49cad4d7aca84a6f4598176f112630e5e4c5f6134ae8a36d513caec1b322a4b6e7c0fa9f2bdce6ba09c4886f505f6d48cf616edaa19979cd56617351f01fd09adbe2a07da1906731c6807ce00cb697cfb5f22331e63514d4431c34afeb2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h199118f73660db8b174e70871e627094e40eee43ac1dbb0f93ebdefe1523cf5e0baa3bc8ab22377997dc50947ffed8cfa47cfef8212768f8a3cbc785a2fb02921839cdd807be2b13e9b6f34430bf148c7b1cd98179ea9d76833ea434712e49ea4c5f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38d7566614f819be1a61f3ab57d4a7c56d68dd857f964d401db3be7ade7f235bf61a6455a897b375972a8d58b3a315e47fb188ebf15bfb1d8ad8e9db7358e17c73e35006de2b32fa91f182ad547203d85b9f59efffb10bfebc68d62d4d461d36ceca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c7587bf43e4c3086f201c5d3753840115578e1d189417bf6c1fecd2806098fd0803f9dd085bb046af35aaf363764fc86945f54b49ad45ae631c22b195b24cd89c4b69a4b55ff8e1afe9b43a5aef22c3fb8e6e2df658fa691620f8f9e09403221a36;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h686155d54a7f7756707f4b5d2de3a611a0e3c224da96cd27cf077e186cb27e0a771e1e34c2d06467b5f497d2b3b07f1b17cd932d8cbe59f1e73b4157fe834c6579b4feeed85e15a7f96feb9125474cdf11e326c35f0e9abb3b0fdbb18611c98e0760;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h73729da373abea2250d9b2cb92fa1d7d59e0f9ee1c9d0a410ecd7bc825460edb15e31498f50e6b09a4442616a82e7e44ac3577399baf38279bf76d11b8dddadec37454e29bd9ebfb4343c1e8d5be358b386094b91d6341cbf84546ac0e4793e86322;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2f4dbe622523d6494979b910e98fcf4679b670e5632e2c85b39476f1b3352c7b697ca90ea9fa2f91ea4cb77b4210c466e3861bb4c5fda1c58c1af78694a8d252597ff6556aba0400100508e0d649d558bac7b4c1e5979f917f1d93c27034891f9b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca23b703890f487726c1d128a295d3ca4e23b94c9d8f1c65a90d9e88f95e0c6c16077f02f95a1c2c87b4d2ee5707ef71485ae02290f1c3bf10e5dc27d4fd609d0a7114a7e2740c0e40d8a703cdd0096996ea6828a6521c91486c6f506d27e1c57a61;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56b8fc17306d7924bb7f4ba76ffb31af2dc1e5371f2e35162f92f197d251c2860a706cd65c93022e72033fededa5ccd3d3a4e62ebac85c7b6709616d8ff262309ec6bbc18bf9be2b9f0e87c94e42dba7af92ce61a01a0e77b114b248fefe09af0a97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbdc6567d5b0443c5170ce52a7ae4106f0e04e1341d0b975d4b93eaa86c5f12b5930c959edb8acc7dbe11f5c9b11adeb2737c925e055c027856f2793f5afecd52205612f9099b2dccc69dee578d67ccdda275f02bc5641197ba8d5d9809f31a68f0a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h776139813950c2c929e6cb5842220f74e67d81df8d09171ca3e14826f2a002b6bc774400dfa3ba04320bf0232c919ee987a4e4a85c4735d61146dcd136d39ad093cb1748caadb38e250609b34081c0b2967e062830058af1b8db184f56212f0afdb1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb77b08ec328bda242288243e87021fa89b408d873f6a620e7a0e5726e4c61333ce15232d38a27e3f26a05db115476e5ac1acd6e03b975a7cbaa314413a7a406c430afc9aa516d7b8d16a9091bd7a205ed883acfdef3756e60c6c5c204363e8222abb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h889b5afbac080e1c2724582d8309899759a832dee861425e317fdd582512c6fbc3805c3b15a80af6be7beb75553098e05b6c37ff1455f16a87b917c85bdbf89f892ac3a72709ef1959cec00585bc03d8a46433e696160ff5b0832671da135dd27bcb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd251a20809a2adbba55faf6dfea33e5f27e76609ee5dff55dbd7d311d32eafc90df12615ead6dbb05eb2aea4ae57afafa7e0aa31181782fb45687e84bb8cbedc90d8d97f8c510c68d459f3dfeb3bb3ea0559546b69d21d8ac138f847dbb53766945;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc97c996176b8dbfdafb0f226af522778caff034dbf04db714ac1fa2fc3e209adebc9881575c563b74024c9e96b910b09ef864ed0b2b5372f2e69ed359bfe2b67801f5c332063686c6369460c9b22ae01596b43c883a8be5a3520ce45e24bb0efb1e4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h189841c45668ffbf3bfad81cc6c01393d11b86829c77aaa40b588450dcc43f09a20fcc41f1a2867deb9c97cf80fb94e72a5d3d3b8b31994efde271831d42d1b9fe451c1c3b25006f8ffdce11d36e8d74a02c561c0c2675bbd40d43c5a240b561672d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1f46daa5cffb06389465996503a02ae2f6cf9a80b93268888d99c3382fa5adc761506b46b3b6012aa9cc66f06d38d94f80346113cd3b63720b438067b4f53998ed3cca3e64636297ffc548fc239d3018c2a212dcf1f22a91099572d261f5a717525;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h721c6fef588fb6ab3bfcefd636da1a7df686786361235d659a4f2683b956c407937caf81fcff8abc220457872f88297cc3142ea3f6252303a8f5792cbf1e6fdc9ae0aff9fbc5300da3db7b1414d90e514457078df9cdf351e78e0c97e23e7d0280f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b40eaa81aa3933252388666933e9d8181e3f8fae338070c0cd573daae56763b46eb7555a7a5affaee1b71f73561b04d92d6ff9f486693bc70a35092e3fc314bef57a3b3fef8e6cc51dac672dfa28e1ac4ce1073ba40105eee27a9af9670f7d4f377;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41f9557d95d9ba2ae3e7548dc0d10be26ed71578ab44c2064f098f2698c428da5e600d3de590552129bd770751bf04eb757b40139cd18ab7ed6f49764157ffbc747bd1d23cca67094a8cfb1007ee8c002c2217db77c448f8ecec0dc4895eda01becb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6be3ee00c724e32409adb586ed615dfa15532e4e2c8fb8bd31b4a78ec965e94ebb73da9cbd3aaa97352e039974d39b7ddfc32038f128fc0ef51d8d85dbeaffdc2b758badfe41ff8e9ba8cbacf9a2fc4d8dd393bd0d24ee7bd5780e4a44c259164ae5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b293ceb647786beaa822ac4111aa543828823c469b871ce1881cbe1b14c0315ccc92e9da40f3f0fc7322ffb511bc2f4ebe9c48593a8912eb5c7094b64cfe519aca50dd3a8e0d3d7494175044a92c0779fa3fa7934e9e47a65afec5c80163c22d797;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h147ff8069586a0e57d47f386a66eee362363e9448d9ab592888273509ada401a70c3822a95295511e6b10f3f215d8e5d2c90882ac03ddebe96ca39edecf2df6cbfdc06dcca286134aa37f6320600249afaac2591d1883f95a2aaea05858a9035bf95;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcc8945bb516603a7b7b9fb1a7a0b7985a85f336e6a3ac21421c4116208f2dd7877f1134e3c8159c7675ff988ce907ce4760992dd9e219db9a819dbacaa610ee97d837e66abacf5866c6ad1ce27e1748226f9fe7432b014b3a42d1acf3983ca5fb53;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5cf6c4079250503f0e84eddc0fd5b607281bed0564f8fb591a8f0f74e2b5d8d2eea5df71b963e9f6885e95115b9e84f7f7af5201d1bb1898eb08fca8b6be0c723d8a6d4910232a06093b60e701350f69368fb59d91cab7dd08b0c3fbc87e260a05b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1610d0e2c79b9f72b57d28b0155d9afec69cfc668ea994ae8fc8d40f7f547c389118ed026e9f58494baafc150f9de68b3375a2e29ecca4e9d3a9228b537ec825b4ee18d430823c0d680c64f14dc1a43477e2148c15a61bb27ada73cfd90f445121cd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ee92c22095b43e027102415dfe66fb9b064a7e70c7a285e02513f5d4889a3eafb4a2f3c1aa26c261327b4ba2349150c61e8cff521f74228409c83491cd85cd1f4683c958326880ac11e43e8a4b4dd7b6840ab9fb20f6c41e5fbcc4b136e68c2db13;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5712c370cf4a54f466308b51fd1a4101a3b346923a43766e3e686110662d7752d8e9d0c7837d5b200526e03f4092519e5a256c81a82323feca9862b61eea7c87130b6d9084808ce03781ff65dd978a54eb76d72fbf2e40154642b69e1764a41daa8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h557949ff9b63f7621713567fc1f82cdbd8e64dc85b8b3e2a2701c2a4b4aceffae86de388752284c069d06d06983e7eea1e5785288a979fee768e39abfb40f38bc6c0a1aac37cbd934b294f689981c1e9b83e1fe07e77463bf0bf59edcd3af55d8d90;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d1b03b7ede5c706a2e35ac92747b0b88d8e1a6e3c874622857dded9325de85fa80987e6d0c59faf55f1569071f4b4b988f1d736e744a0128eb7dc5511858bc5886f6e3fab27904058d8b88f2e716068a66134d03032c872718cfaeae8c37fe22188;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3ecb2345d3e568ed744a3789b7b2821fa37a7c7bd0b416179f73ffba1777591843d5f11a9c68e4c6074d2690fdb033d23f06390b4e301d001840594afde964a5c6ee9aafcd4acf93c2f9e9313b9f95c37460eb8f0a53f5fc839b388899f0ba922a1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45e713e7b189d66e3133eb521bbe02e1c472dc29ffd8b5af555172d9ef18ce48692cba421ff9664f4f8e8c678f30338736647c3a5d652e88695f2603ebe14c35293dc5f8cb8a06de3615c894c21e46d6c0c2408470ed52f4b0f2724515e242355865;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h445429cdbdbdd77f025b908243de8251215bf6c636e6e37c88d418cf60d1f9696b75f8220c4894093b43eff159cae54a030504b4a64f9e11ed7f7ca2324c9cddda6c731918ff4d129d29e748b81ab2e2c931b60f5604e6a968d342caf2dd7d788e02;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5048d547af97a36bfe2ec8ada12063bb098e6071a19eb261b127f39a9d247168cebe3d94f79a96afc5410a052553d837957144518ff66e47dd058d8bcd910c38a97badf7a7a434b8ef63d5cbeff4b463655540ee93c8082fcc912122cfb35ffecb0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91a3310423b858391ed2e9a05468ea4fd0ff187fc601c7e5a954806b82c953586e4d59c1aa35a7a81285d27fb9dfde129e7cba2f10cdb15259aad758063d818c25838b157fb8048bb66d93efeec80ac1df38b42cc3083392bc2051da0bf67ce22d8f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea933aaff305fda5d5e4ec489b4fca687466146f172e6d8ba5712915e7cf03249c54b021307f2c7175bcda5a9c0f55f7585d97fc0f052363d9094d40fae7c393e8e99fb8712fff67625cb99fa74e430c6369e38212f2f89f2f0aeb430bec714fab3a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b5edd275785c827dc545522007aa106397d82bb0d6519f180279c9f90d8afa9ae9a2b6d24fc24d17ce8579fd579eb8ceb5ca96640287dfcbfa142d7a752b21a16e6b7e7c9e81f68f20eab479d97208a037ce70d90e9681eb26f349d918e2702206f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h682ed7a5ee267d109841c86c0e603d8476139187542567559eba6596754fabf6d240633229ba12eef292c23da05ac747d3dbdf6016eed2a029b15f90b56d7123f858bf552cd20f1df45e14fa621de824044f1dae7daa168afeeaaad39186b178fe18;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2714c9e858e824856646dc64449c886e7bbe6c7e0ca8ed684da452ece9448afdfc575241546557ccde4d614d2a662dd6f3da429c80df55a695f1fcd8abb4919bfec0a821e50a7efc2bc47ec8fa6e0b1bcfcc1716d50d9e6a751479fef4727742fb35;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he59e8e6be79d19e1aeaed9133a7530e04d9eb5d873737e2332923398d283b393bc3cd2f9913dfc950283f05478a68db9142dbb585d655fa906e5f9487776510ab03bf927ceb338762f421ddc552cfc4bbe31bf8671fd9a482abf41adc99d5e56b01a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcce0f8ac3857e4a6a6e27a2d3e35c32dcb921b3957ac9ad6e96b5d4dac5ea944049ddb1398e2fb6392f87d3785b47e15b2a504de0c2f037a3fabc43030bd77ca87368a0176367903b22f6e1c13450e2a87c01fd0869ab088f49a48dffb2c6f2ea5d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67e9f0262faef7eb518368d7bfdd7c423f2fc640aa0d3ccea74228a58816753bb93af31b726cf4690e75d4b643c5d56fda8eb05b4c9faa758d6a3c0e9f24620680206e07fa4bf6172be25e9004985c37a6edbe0396b871064150dda232123fd56451;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h539a37077e6bcb31622c674c01215a730424f4d510f1feea2c4d06038caca86d20a40381dba6ee00b49801a19732235af29a98b48382d4d2c9988d681e00dfab0423819e9be50d7f10a239becf00556c98b87ca3b7cc3a0d3031412fdba2f1809cd4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hecd950521dcc82aefad9a804d87661c065b3a3fa6cffac6b0f7c85b960dfcc1ac94c1871f9b8e2ff84a06560d4dabce0d8f923dbdddca59ddc75eb859568df863ba674c313441093c6d25b1c5092d2a1eca5bff5974661aa6943a596ab6515b46fe4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb20d5112b26dd184fe99703f89ee8ef7ffb7023cc08bce846426f65c9dda5bc71b0d47281fb2fb225495cc89777b3458e31e0d3d0977ea20b3d034257cdcb46ae4bbfc38a449176f89ade39247733643cfc5b74a483eeda5ce6a591c16371bc76e41;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haede13d969f92d1b4efec280f8ccd741b7f594533a5729037cd19449bb5189ff74c4d293d21b1cb33d6f98e226459fdf0e4edb108dfe5bf1c716334d21a5a26612c0e1a6376ccab4c71cf76711d2999908261d1b83a8f753430bc4dd2c7ccbae6ec6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42cb39eecaecd995011a806aa7b9bcecc60e113012563abb007f7ca2614c03cef72e5c260ba23ca73632662db50457c4563d485a469e4046de7a64aca99834be32265ef34c2846fbc379fcacecda92376449d99bcd6bebf67d843a97ebcb84e93328;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b55e6ed7a42e4a1150e51074ab07ea7f940e5017b44eb5bdb1cf17d02e19dd3883ff2e76800c382e7658879120d9ba7cbc6e3b0df99ebf5dba05b7bd673fc23f40195c9ce99752270a44dc7a563b486a70ca89a36c6963a16b35b56b644c446cf0b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ea53db9d96c2a19a73a0edd21346f29cc0a2b071a6d798b789c8444d22124f3f1e409a59aa0b080985fda6117b057a78f3170618425b849baac4bb12db59d54d458cf0309a727e5eada40ad0ae474d4273b552d402a46a8552be6fd5e34792e925d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f39acda4eb05801277b44fe5a53dab78252981cfe5dfbf12dd99fb3d23f8b3fef6122608edae2278f88ec6aebba38b4102962d82546b7fd32b98f0cf0f774178d5b095a79277d81e159cd4461f74aea638f180844234dbbca25ea07c8eef0337f9d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20ad53c52c298c783ad1ef2644bd9a95dfff735d950795c567dc0374b554f17cbf33b5ab6a3999a814b8db0627728391bddb5eb77a34e1722399f399ef204bb5aae60e64816cb01a9acaf7602696826cd86e582aa8350c27caf1239dd400d6b1a04e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf173ad657df83b96cdb5f2ffa8fc3086e2dea39531ea172576f86b814ebc418db4e35f1c4180d36cee844cc7f3db9f1d51c1108de571a46bcbfa015f596fcf830f90133f48d5b9acbd2b081da721729832c0d86b681bf4a210b0def91be3a73ae59e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a09d5831e78c7958ede0723fe01be2377fe976384ed9433ac562a66a382c7e41c4000c40405112f5b4ca3314a0cd4dad49a10c3b8d0a4dd70556c78fb641614322376df044f3f7fe75c1b9d51d2fad92102bed6451a2f624e8d5e98b7007a34ea24;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed054f9c336240ee17c7b099f2666ec2779821257db1a1c475c77eb73b6a1f24d0822de90e03adee5ccfed01a5c81f95046d9bdd4b12fdf89d0723f89f7ad3715c973666a444cbc2fc1bb16202a889eb422de81e210f21c8c7fc87d2c8ed11d3c6dd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he08e39e5a4fb2294d220a41454fa58c7a1e4a24b4cf348a5b1a6b515a9479a44cf6ac8820e1830d4aadde974443667e22838f6613da462e0760f41d01c59903b643e7f1b0fad6dfa5da8ffeee7e0b3a8fc13e01b094acb40bc070a927b82671ab22a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb039592dcf198fabe2bd31c64d6f39cb77ce4b9d600613f1424b0badb66380704af276c14de795b5e960d7676f26f19d833a0f1f3e21e1c6ffcbf53ad5c89ec00f3da66dde3ecae6d1ae62294ac1e53dc1911f63042fd88b7663c2dcc5dc441160fd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5cf7ef3dd8af30c755be0c8d6ddf7cdd5e0ab168a5f879e762329ae5bf315c077e0d4f50747da0a813798b0be7139f1de065a931fc0a8aaff71f0d4ca8f5d9a3c2a9cae0b05ffd1dba06f14417241b455408f235a035bba3c8c12bdf69bde482e3b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9b5d2ded30197b7b4bc9c4a1f337ca59d7eff506b20ba4785cd19e44ee5bf55c9cdc6a059457f3ea67a37ec3e46ddf8790754a10daee1451093cc702b3e436670cdad437e77a20ec39953d77e2153ee50f9c166af323f7deae85cd95035bde78b02;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb07ef002aa3b1c319a91290c39e55c47bf1a0ddd2a851ea0fa2e03d32fbd7820435bc5442e69670ddf35ab3a8950a7558a9713a890480b2188107e3a2611a9442f29e785df7ba2e3118c857349e24f3eb589490f9852ffe8d7de0ae2cfcd53014e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1167a4abbbcf2c93720bd7139624f808bdcd616e653b0b29c9b9cb12c3a0ffedd61dd47f4bbbbe80ccd1f6d06a63ea3abf10db062f2b9ab9503367a8fc3adc2ec55eb1c091fef57a2fcf6626a7fc116a4f5e7bf99fb4c70b6af7b4072e7a27c4941;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26265a1b2c15c4cb1f07dedb22ca7b1229762b52111caaa103685c1698eaa30ca5c9353cfd1fe3515162f3ef5e0d279e1c71b662f2ec500dfc6d781db77ab3a2128e32da9b61f19809c4f08a6eadb9a254f81322e906db32699d5b09f72e59e7202c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93aa62751a454483043d8c3be5f001a1d18f5040aa8ac0bb2a6326c9ee3d86701c953e6eb32f9759c0b0bc378c1aff2d425eabc70dc2baabef1e7ccce6ea8064bbb69af7c838f07e328b595f99bc38855769325dc3dc3b8451153e3fde0013a788b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bbdadf817d09b06e47a1b45e5bdcc498ae8709b3717b9be537e356fa05ccf5381144138581262fa3dff3a062bba95dfc9190f101b56968d9d37aadb3c001e49a860c9a4f172f61d8a9269259306ad45f61443fb9c876fa43552cea3ce23abe74956;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb688e7f73a7f48d0ab32b62fa307f6624927af958a1b7a8826b73a1cd1944b0644c806659171599a1edf179b0dfc34b83ece97891e78aec46095bedabf7ad906972b8d51b49ac7aa14fc64997585a064a7f7d21e0c3b085fe3e240f14846c9df7aa9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habafc166d2ad4b5f822bd666a1a4edb6f3f3f88efb8a32bc77fda6b59f40859faf5c66f4dc0f30df177ba524d5d096fc7590af7c3cc14ec5cbfa6634359e0c5438213c1db82583eff3cb8b59c01cc75ae5e97fbab2ab3d53d8f1c0056342db131903;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf75467f9d8eb9a27943d7a4d8f5d9ef236a06956d8120502632259d07e94f6d168de0c98573f84bf141e65b58ff179b9ba67b77d95027d92f1779cc32f97939f6d0d0fd3dfbd75ba1d84631a842064b4c4c507d3a23dd81d26ad91ce2dd4cf5f595;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha09dd9e5623bc61455e38f32f5af0bf4ac4d320ba0c661d4d95c050bdf081848c28eb584b3f76a886f858d3e153bedde91fd80572729a4b640bb7c0aac350422a05fab64d14e2e0b7e19cfb1875f543289e6cec609f747fd2b72b40b828557b1dbdc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac376e32a75cd075309caa8eb28fa62051515e23a62c0619520fb7a51c85896ba5485f7f8640627c363711206f26bf4c726d3ab5e70f30158c9bb504b274168ceb91c2bf0bd116bd1baeab1dd8a54f15c0538b938f4c2193de25e22aed193b78ea88;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h209112dec8d825c37b6cffe203de7a29226b1285f82dcd83592b2d708cec99f15c2770305f1ed8d5dd5306105c12a77d6483e3d9c565ae15fda891167b8bc7ed53c4df0c49099d4d27aec1cb075ea47f5a6025e11dc2185acd57c03b10628357124d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c30865c949ebefd6883e069a3e2afc78e20431d923538ef6bc5ade744ca344c9c4f36b3ba46739d2529166dca72c719322e4024f8e5159f4bd8dd325089f433e3dce6650bf6e13189e16249d02ff11791c35a41841488322b6c539682c1734e11b6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3fb2f5e08e8721a2a3a62dfe1a3145c7bbb4a3d02126a36afb8b8851e9ff508d1e544a471e92364ded1b8d6079e7288ed314bd3b9d9ae82c04400215829761be5eb8cc0763127478a1034d515e2e2844cf86f8ae5524f0392a768c6a30fff21547e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcee73c3827833091b06ae28e93330bcda0e85b3995aec092e31e4b4964fe3d5fd07a8ca061d8b802d512f6c47098bb8ed0407f88c36e534a275f6a27069f9b263a37c2f7dafc9e09cd0ae5761145c1d9fd91245847d48efbdac80ae4b8829b22a81d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54a2fd2a0d91dd7bab535b74e7bdfa0b83132739ca6d15062aac26fed15de0bfaaeef3580b1636c1d23293043724bfd9f11c9a1e1a9314fe0f0ca47ac6d914aabab6929bfbb66ecf77c8d3b18f54d6de656a2dc563be40391d4dbba6a0b42bf0f05d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49e908449f4b19bad0fc6bc2ebe20a09e795575424bc44bcdeaf8351872f6a89aafd7184a1575365f6d12170db82ebff3543658aebd2b4e05b7b49771fbb21598da4d08858cfba390c55c52a86542659c829490189162537025ee6cde8af0df2c92c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20133e45194fe0b05f3d5836e7d1b535857bb001faf82b5b04a79dac3f9d553ffa0dd7be170d7b1c315980f97b67ae761d2cf5bd308aa0e064ec3972a2105636fadee229593b28ef7657067b45490013d6682967d8bf7ed79f3d11c069b6b5fae25b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc32976462a093e0a2ec6f3b1318a60c6d24e9c5b48e612598374c5ad1b420eed0e08abab028bdc81b19af6cb0508ca5a98aca20b493605c4575da4326165a02f6f8a328106776f8375717054f6b6bca06b80fb802d077e28bf1e4cbb19b5281235ca;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1442ecef14e376e6064fabd6abbae39b688bfa2c0fc7ec7f33fd1eb4646bafd8821e86244dd225b574ce4300591d132eee139e05da4ab9d05a60cc4c5bfdcd4ca14eb14aca80fc8fb1f8758234d88d8698d370a28562d0398d9cea8af6b681b086a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf9122f79d7c42642a7c5627a1e8531c51e1213b98a5623c296aaf660372b761c859f371d7329fe2db394041b735bc165aa8388adac0e3d62e62314a91dc775aa927ec7df08b750a016a588278490e28e4321faf10b75e779f6eb8a2afdfa8c487d3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he25b884257b961df133390647c83d450b311c787e3064a17d2679be67ae205dbf7affa43da0da5f45b483cc0dcbccd8901a5c060149d2f9fd2f09773293f3602f93f4fdb9899ff447a75265412378ebb298e2c8c92177ebec075321f51590408df73;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62423a9eb5240496ee83eab9d6a05e9785bae814a8a216babc8ed27a82175994b8ca177704605e16c5dc415d2e575ee472a5bc6b92edb112d186335999ddf3a363595610ebbf420318fba0f27df8c201604a947a49d88f15928decfb4e39e3670328;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea5cf1bdb9d09fa31fc284dcbcdb6ecb79d3e351a0822852f07ff1769fdc1b88bfb16ca26c5f6cb8ddcc3b1817fc1c63bbff000c26e09b02062b113f11babc1b94c0ebbdc4fb333219661265fa32d6fc5b3ce2f77ea2b5a7fd225cc6c658b8c72d58;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f2dbeae9f81f1d065af75cab3c870c0e263a922fabec58dffa5f0b73b2f44622d7cdd7e3b46286773199be74fbd9d0de7ed6a73978f1c7aab35160f36747b0a2fa4dbfab2b31589b36387760547b449f87d51f9ea9cd1443c0041604ab10a758db1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe18411eeee83f55c92601b165c6df24b200b7d948592a5cff706e23ba0bd058ee29569c06e2271b8fcf37a43b3c25848a13aaa3a76d62751612a5ae050f767cf26d643045f0a563fe3c1dee2d0a1317df2bab5bb1c81ae1d0abb4103dc22f5efce6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca3e929646659f3a66a81e25ada621c8024009db4e68f9918804b33cef9135783ee06a4c46afa28295ea689cb8f9af6bd02a476e33e113799c920b64843b06a56257d2aa38617db723bd78c4a99a93e63d9c9b994e0f289410846b9b93147bc26df4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83298a25d033279bb798d0ed9e04ae608a5d03c07ce5be83a490e00959295f5e08796f460f0b20935d05a997d056f2ed183bb0243f0cf47434b9dc68f5453f208b9869f303a87b6ac676b4f1470aa56f4f629515cb594e2d6426e59e9f4f9ee8bb1e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5cb6c693b16588597b165c3d6b834328405815690916dc1e77d17da266830c78815d2ce1cbacc8c17f8369326e73e61f99a54bd474ecfeb4268b93b236ca82c1b5d467cb7a2042bc0d63f57197d41c791aa29bb9515f6c05707aa395a96023550e01;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6036aa14637c449a80cd0d66fda18c9d79100da20c6bb2064131604c94a0fe2f0f413df551eb93a4eb2f618670bf5c07548e80d8e92824b36a9477dd8a53b6c12939b5e0fcec6fa78e5534122b020ba1f7497afef2137cbefffbcf6ebf3dbfa5367a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5333ef01f92f23e56970f0976a160d172fa550b63e33728e6d1fb5fe11b726d6b33ff2efc41127c5caa7eb5cdebf4c64af18a691b329ee7267f5967ca945e58f0e524c1b8e976d1ebc5b0d7991c8a4e4b635e6ebae47e12c33196c7c79d0f55b22b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h426fc086bc11c7c2bccfe2730b5106741fd08f059b1a36497c63bda7d4f58ae9a945f5a4bbf5ee9aef5ef88eefb9cc5e2d6b6d7f5025e6cc277a8379c189b5e1f5f1a715474c1c2be6d5e8f04bb626f8a074670af40e361e1fce00bbb75be2c4039b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h169b5df4b06a8585b49d055703d437a35667389d6b3c1ee88601adae4e916479090a459068445c0e8639095d6a78c93bbf0823271d1c4d96dfb11cd70c1ddbf9d38c04599c0616687665cf932997236465b0528dcc138e2a0b923660000da26e7c0c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7f859ca3dde9ca2ab4b22e93938c540d5722d9e87e02852fcd9a8ce9cfe7cc9f6e296a371952a7c0e48b297d9c4ee3f1a6be12fac0f718277f901ebb92d2af582ed986e26a76459c9f9dbb82416254c6af668611d5312760f3c2a49170676b1c98e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a3ab97449d9fd6aa369c9087047743bad0f7780f51c3b2c6b6f2dca81b55c10138198da1f1d5067bea772692f8909b834e75107334a3d47a93f7f654059c87f710ad4b660bcd04e193c68b20b162d0a7e58dd2c5c7bda86d706d38c440ebc56c7cf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c22a2715fcbfe6c553bd025663fce1f2a34cfeb1af63052fcf4498cf88d8a9e4a982c17907da2d11290194f131caebcf247a246f50dda87f32a42fd4eb28b4377fc85e26d215fc4b1bd4f32a5ad152d716783ca3c0c1b8de7fda6274880ba8c0dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6521818a1b18d27a5a661a4b578900f2ae78b920f2f994d47a2543c749785b10b3b72d70e2255a3cfc23eb7eef8401b91dbb3a9b22b6ba42be79ddaf128735cc72920fbf9593a66472a6d54844d4b404ffe8aeadea55166abebf6d0e2d94c481ece9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7b63c0e471b245a2d65d71fcd62eda86051c3b716067ef1ded76e4a8ea37df0db01daa7493a3fa67993daf92c4106a1e94884414d27f44178e2c153176d6af074df0e4c9557eaabe3bd19d3fa363aecf4405891db44d11fb3262e21bb59654b09df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha9c6c91f04a75c4913cd82b31bf175bdd64286255180bb0ef1a780494dac5710d02c2321b4eed6df6e009dfc47acc5ba805349ac4408d228921b416b088dbb0295da9018f379a9c1aead1241ee238603d7f975c103ef860caa02d2578ed3f4609555;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f40abb84f7d5c15c3cbec69e3ef2a8d2b045a0fc567cff39eeff71c14a50bee01f0b815f2f7314b2431b50b2de3f93612c075bb0af87af8510a9fa2c2e8459c1fe31d13965ae484f2225a83f732c20aed05406978a5e91cfb94a54970743b888dd7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd33a97a3239ec4df76d81ae7aa35bad0cd6cad0bec2a7efa6ae15e68fe2eca857e258773ee4ed93f92233c1ad2c1fd718cdf9ca29be6d845eb1daf16a28cc1c10fd0e1b2daa7d05d48b7c10c67bc449d74ae71124ad9ec402ef1218b55b705a46a9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a770bc3ac8a2e631b0902bcf443f37804373072654fcfa626c30fec99ce2f5a787f290b6970f271c86c5d2764647d45f612e37f97e3b5aff4ceb70e6889ffcbc1a6ca5731f0b29c5f41e0eeb82f772da66e5db63ffecb927e19487937962f23fa9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h783855e6c05edd2dae162e4faa8768b66ff4f4d5c5b6794261d800930a96796efedd71c4c613d8923bec2e133311383afcd591b67798605722b66244396bc23d659e9f53fdfe64695a33e158f834482d9a057b6fb3f54ae97b005bf939dc75d03f40;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h216f819cb6510602970e7c22e4e1ac2addd3ccc0aa50413691a6be324cfbeaa84be6d51232006a457b87a2d7013a8b1639064e7e9a0ce3312f3078312f0f087628887cb8ea042ab737fabe0418c67c41acafbcc7cfb7af867738938d03ad4115e91d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3977652a9867da389f5812e1d41203f330c3b2c39dc5be9fc4c55f2ac1c112fb47056b72a0ba0c56b256649e35b4485a3d3914c959ced1d55528eee7457893b63798167b9d3ec94cbb5d1b7cf07daf8b7fe68b2ac243c76bc4eb7975460ea11e6fda;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf7d8d7d69b4d75dc71179fc510041e406ac90feab996acaa590ca2c4010bfd4711b3a2984fb4447578a83e589623431681b49bda671d1e1bf41733aed718dc665dd87c19d45271def0b2fdad084a4110738998ff535360a7b319c62d000524a2249;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had5325bf46446a37dcf675e2bed5935834ab5371d7096b54d1c554e01d745fc42564c77e0900c793e7921164d68a7d947d1c2e4a1aafe45a888670440298ba527335fbef3c1b1cb151c4db69f3186e5855d462e70f7642b0f7251c910abe0802f478;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc06b653c14c95514d51dd6062b8081ef81d2b70554eb0c6c9639a2fecfecb1f7564e494c97a60b392e8a09815ff1ddaae4a15f2d7e40201be1954d9324f082ed9e6bd42c961ae41a11aad20d8764adcb1cf05d140f1cde9a3da09e8b6573ddc95b54;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c72a3dcd5ac79df457f68e3f89add84180d543d973052fad8c2d2d7162b941cea39018ba45fe6d539000a8e78997a314fd4d0d046d49a02b1058dc0c87cd2ab890078f1bc7aaec432a05995c470601abd6b83bfb51d11f6a211dd021d2dd75fdc58;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcaaf732023242d2b2bcafdc6535405c7ae63e5b17a40a83a1a1f62219479fa5dc7f4254e0604b8cb6a8f314cab806e362bcc5d22b6f48c2cc5eec94889eaa8fbc910a331e057b4ec443c32f096582d3cdedd9c9eeec8893dbaaa51f17b6bae4e900d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4be0467d711aaa0926b1a4ff67e4b3ead8692b8f389c271bd1b0ef15a74a02ad55bafa075fd72a37fb85f75bc8ea9534100d77ce8ab5b331fe072b8c929b2c36b84f7e3c296ce24c230e842acb4304dcc652718e5d9bfdb423eecb80dd4ff2a1d295;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b0a93b190eb40ee66f8f5bd9b552155ce435ed952310f64022029412d5da7a31337ac26738e7813adda17622fbb8a616848594d5f4f26a14b9e79dcc028c2f46f09dfada6d1c25352c01cfe63e213c412787caaffe32fa8a34df37a1e3e1bcdd7d2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha90463c627842ef97e13ae94b75d50f3e56973bb02d373a347cfce621b5f404354703cad2802f2f61a03c24604ca75c228890e032a84f5ee25f5c4552c3966da96e69e3a3a9b39babb3b02af80037f4d58b3a950319892cf088299561f972046c395;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c13fa51ee64e292a7d600aae8326e62a5899d125cae135754a153d6656f43986b80316efe6f3b899519d3eb04da474a223804f20d0ed245ba6cae655215aee4b04101a57b113c2aa02e2f84462bf513cbde0a048ce719b74d8d0812e65c705686dc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbd9e633b9f11f063927cf91b4e4a0d170cd0b88a11b5b98dd2c64b0d12be7293c1b60a3786ab41fc4a6e825fbca605db77f0db0dcef7907b37394cd16af0cb7b7fabad182bd8b614fc1a3a6f1b852582983f7bff63127e078448fdacc520711ff2d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ed85e79a9b48df4ddd3d769d06b424fddb2c3d0fd3c219c5932ce7fbd3f4f14dff533970a457bd6533d74a4007a9caabb6c37d50eedd140954436d6e559b991894d7fb4b47b488c0db97d685969a20878dcd8da4c32d22ed9888a538bb86db86aa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72fda4f291693d672eae33ea2deb3f8a5baddba4c773bb2070b65f5f656fc7e81064fb4aed7f19cbf05e6a526cc39487dd7d290524d68995080dbc09e5b1f8e10a1eb71572b8942fe3310852714c2e85cb6cde689d53f7600e734c1030c5ccab0739;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75d0e3d3be867544cab2c34c40ea67a39e5ffb16cf27a0fbb8782c7e604b4509810d7d30b7e7a1a0e329d07a1acdecb969a5a5445eb6a932a2dd49b4d338bc869b8eb6ba73009abbb1df9441e08ea4d185f0a87634cf246055ffde75492e1fcf7b63;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8cdc7569e24174fe13f4fc98bfd2bc0e982fa589be281bc6b9eb2db204033b01d1d7e716cc6f5054b094e086542d0a480c51f62c4f1bbf24973208f83c932e157419efac6c83bd967e8c3c239da2e7f737c19f27f16a8976989ab5be287475672618;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee381bed34fcd4cda4924f6dd7612b26b52fc929d50db1c9647e7ce45e27bfd6110c18b6c0874cf7f8c5bc8c3a53450fee1a8fac2fb68bb2af1e80aaad6fc82d3a52c345c203ebaf39df4e0a38dd0d5e4fbd959d4af0390c0beb6d9d9ae4a8482b28;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h992ae3f54a1b8688f707f9e9a72dfd2ced6be788fdcd30c4edd914f1ed15caef94f66e3064190a25bc9f0639789ca28d81566ea6ee390163de4a6f7a0a349bd16f83212e67d4a9075e9d0c141366d08cdd2fd57db6ba3468be7067708ae9c2fe2fbd;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heabe6a80c1b274a51737d57b3a5362bf65f3286155bd1c6e2acd02f3ade5d1423b041a51edc5fed8a5f441c1a39462be2921634e52484e3f6a347e9dc99bd97d47fa9ab0b640a3380dc3606d7773b2389db1cdb66b1964a968ecff5c7a02ddda23ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f555453570e86af0064e16c1fef296bdbf697b3ee9e7903f305c29f1992710c4890bc79acf9996e1ff5a0d2100a019af7e761763bc37c5fcca77bf3df3677735baaa3309ae3883b171d3289186b388f6b79ca307ee7839093bb886e93a30c81229e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc49d248688f65cb75003ef43ecddd2e3341f36d3167a0d30224774ae3700e91df614532170b13788132cdd8cd1bd98abaec3b2acff0ad1f7b5b7f1d5c4a750a9a1528c71387ecfa15ace7f7efea03154eba04d14d272c0b1f5ae0c0ccff07d4998;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he93d8f272989ccdee899c620eee06fe37556d8cc82fae841999d1ab2984df0a97e9ebdc3f36595182a2b4b3b9de35e79e629eb48033fdc07c78f3b0bb1e29dbe1c851d5f4d6f8d1b181123c4923e3d4b22d6be20a35cae92897980bb8b6a50fa24b1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58c2513e92b37b1ad5ee312b28730ec7b65b052fc236249223b1dd09859479e32e2d96ef8f7e67b2092e58669f439369ee93858ccf3fd8b79ad0474ac1e091be13fe2373e1e9d9e855623cec367d04994b50898eb72fffa8eb5399aa3d9deca8b4df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h876003d9ef4a69af940e1e637404621edfb05cad8d7ec23b1b29537ac91586375bc8a4eb558b32abca26627fc39234e5edf4de8508a63c03d582353b621a289c86755f35c0381e4ffd37b9f7c652709755ec88288c226ad72b4e7318a7f9728341b6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc39c3d4839daf7025e9cd68afd418b1c3eeddbd0dd42e2332634bab0d1de78d9e9acc4872a6e7b979576a7d35781327e98b309f5d694276cc223ed1020b6f340e42cbcf1403bcec803a53e8a6a348aec4d58e99213c28cea42c0c8f2ab2cfaecbd87;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39ebb53f479ae4988136b9f4341c7de6be74159d952651e8de16927518b2010f0279726ddc0b0bb2318c320bfcfe6e7eed8dbee0ea67c459848480a67cddc3f7698130265897b71c04b72e0aafc081f2bff179244d1c167819d586c61edbc4204ef6;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43036c4d085fb04ab8303d29b753e0d62c90ace118583936c39ef436b92c99d36d704ce9216ec9c80121beaa00da3179c9c19ea03038fcd4b5b54fd75786ca1ea673203917b2803504de0041f796e909618086ade98b441542a13226dcf2ef2665ee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h905e7b2df3dec03b0ede7fe87f4bc87957e378c62595a0b1c49917a09c88adb144721e34d4edb2716c5144dd8989c71a853cf6e9c7c3d9e36ce70ee8431b2d36ea24b542bf103fb0c6dd777ba5ffa3bb41e8fe1bc2a7d9200c4375949e183b5572e4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69980dd782fc6733ad1e70f2d6731ee2a95e9ff48e8735e0b47fdf7c6fadcb1d5ee7063fa57e0f772e72c9c5f239d3bdbaf48e9ec12a3446cf421d4b099944b21451354bb0249ec6f759aab00febe4e5a4a1354307f8de4f9667a6864562e7f26662;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hde7cb1744ba3099451e770edbd1712b9314bf256b9b3299d55b9c3d485c984321255608d62060f67d15ba6d362f7344f339724f83d68a1583a2ebb1d8f30b18fde28b0bd4ccb68d7ec9c4d707f94ef22c682e5cd3e0130fce2ce0dd2720aff9086f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1bc0b978255dc2fc287bb73174c40533bbf1d9497189ec7e2aeae35cce13bcb314bc80a7dd8641bf03700e59e759526ba2926044e5bb93a133fbd7d8799fdb58eff25213e6d6f8b13b79b13e8331f6336cd0b4355e402c26cbcbeaf0420fa7c63f9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf511912f8852a828918490b36558eaa56b3f4c251adf3db3f540d5c7b49796183abbc0a8656829237b5eddb3b35a16d23456c63e0befc8fc619d949b9654c804c887bcfac0615bd3293340e563a371f277dbd08af3d64008a986abc234672a3d5560;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h457de547bc1f48cf44d4cb5b236f8611cd5aae8ebd0cae5d61c4aa5dd94c9188accbaf7d5bd14bf89fd93e9a73b7592488afaa0172f351939af5fb8ab0fa66c9f323055e13f289e50f8dc5adf62a48157f6b255405f9462085aa94091275290458c9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd36e7ea98d399022ad9dfe2afde049127cec808069fbd0bf2da75a00e8f4ffa5c76d2019ab6d933a686a3d676808229ade4dbf0a0897d26842ae552eb56ff5c124e736bacd77ea4da009786f42b93eca87a11af08d37358bcb1b901cd37294bfac96;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5863b06c70d1d174134543c31a9a45ad0b82c18c7e55030deb39912c8a7de3b8642cdcde788b8664b18f75fcf8b930c31bf3776788f468edcf66d38da735d8f75d0d3377717fe996bce82700676c91488e02cb8ef4e6aba70d59c6552ceffad28c7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h290533c7ec5dd5f3e2e18c866b668cf9bb09a956e78aa82451f6824f3b1ebb4ce7d77234deb16b4aa2b0d37d38bbfcea9d8eff6b96f57100ca6029e0f823701c5f900c6772ae410e9eef98d6d7b7239e410bfdd23834bafbee903526a19576504c5c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b79274a1f70b19f509aa81afa1271fc087e0b880773ec464f369efbf70947a5bd176ea9079fd1c8f20103dd592edbad756cf85b3806144bd4d232a67e3af5d639ae97aba9c4a6467df1c27aceb623988c81a0065f2df1f5439051db6c9512e615f7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f1a2777875a085363b65c96a85d71e5f832756d0d6cfaffe603056f6c6c2e511bc8e6c3947b0cdb5a89601aac48b932b00c9b65a9b23a17bd0922f71a9f6f5f72387f2a6c06b2a8383ef6ea55868bb442767afd99bd0f5cf6103eb76e6778d92381;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h59728606135a563228ff1ef3e27490a02e8b8e8174b7d2d7a0489f803f8b04139144ca2aa252480f45ab66e0dab5e8679b7bfe2c8c5017da3c4c1fecae6e57b707231b6d8f84e1fb1578cc6af7b6da25b9d38eab953eaf6783e5d6eef123efe7f1fc;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a783d5a20adc0299d99f2b7ccdaa026d0f690c3b3578ddefd86ad756b6ddb7ccf07339d9b5a04c14efd3515310b9c43928a9c07e06167ee4467c4caa823942e6884a6aafdb6ab4faceb36dc54dda6964dcc32b219fc28317aacec5d864224221b48;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h172a6301c4c27cb9c5b3fbb4a86411f8a8458e231bfddd78363af877842961e0cdc0d52790f943228110b60b132dcc128ab3faf6cc571d6c2e14d42cd7f5ecd9078ff7a7aa3e7cf22c0a38902c58bd417797e46b3451b172584454170f500c5f972d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd17ba55ae80444a0e145314665a5cab6a0c8200770c03fe2ba7ce295df37495f2dde9d6ab54a1b261caf292e79663f23a88ffdfc8e004c88efa10c7e395fc626937319121bfe3f234d89354ac5408b2f99e5923633fa5b3cfe4c31cc48897f04348;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h147a2d6e28ec9953698023fd64bb482338090ad0d0bfc3509943774a467f2fa99b8ddba3f253ab4bda0cf1cacc7223f60797c5a5c8dc1dcde97b8825520c34f54adea01c18ae4eafd62c44b9177e26a899498873d25f11d32f1b16bffeb3d7584ce9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9591a958ba3d8426a56a7f810559afadbebe95c2141e0646a2d5274cdcb8e0b65016d6df63055a0eff6ea9b34f9f3d0358bfc50d3b6d40bf6f2b1840c985d01afa881bdb171e7a94d7418c8e716b5824b7df08e01f13febf396d7d25964e9d6fec7b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f2f498265145e77efcd95d96ec41227ac1d36a61c690c458d950cd3872938e9777a9d86ef54c4a53b37d359c68310b56a4691b270a73bd032abf7413bbff32794f40059fb6ee0872a790d5e9f6ae85ccec69276940ee4f1b8ed2a72d47c3ed96cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ae15c5af5649b53f4e923702762ed6f12439bb2cb6fba7771e94a0bfff0d7f8434f9cbba1a9a5755afd639f1446475299f94d9d341ae6d01f2cafae11dc721266ea2ae13cac40dd95e5621ad0895c196c216151c05296a0ca489396484324941d94;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c4e220c42d5d7aaf4c4ecaf7236dd8cc742126cd925a7f72fd74f7cb1404f4413af2baf76835a5f987c17204b6a0661fcb6c336a0ebc120d40fe2e584d6e62123fe0c355433a589875c29f4607eeb2b01d2d70426898fbf33089682271cb9f77324;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb20cba200a8f6d296acbbbf8418d965fa45a6c19d93968857f8c274f6fd5bc6a748521b2db1f41ec8c115ca5ef32de77b41363f140d17a6326778eb715a7f37c3a0d643a7ecf6c5690a8eb82115cb704e5d3859dc0e423691ab73b769e732e3013b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a77e1187cfbf4c5e103305edd879777f2ac04a74d48bb6219b03eab277f2320dd2246eec8af15c3d0f9ab06b7d35332bbf804ec5a0ccd6bbc74df0a35ceaa3c976c8991b170765e002f5bcd5711592a039fe90853d4256c030f8cb9dc50e729325c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4e1ec7430ac490a664f6a6b432fff96a044cebf128dc66cf32252439c4e4c4abac14e2c169f9f9cf5958dc20b434b9ff122700199108c67c9bc5b301065745fa4db86ed170383ed7bdcbe7b1c31f81603be960f0e1783709a97a3fc4c804f2f1ef;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bfde656e1baa00f534009f27c8a47fa4d9a25da97afd4912ad6bc3ac9a632da33b23a20fee2d43c1a983426482c5b31fee93fd73a3237d08d1b18b8c8ab94297f03a7f12078c25fd66c92cc1d20c9bba0f954aa0c4d82965dd980b89767e2a6681c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd429fda1cc38c6074743818f49bfa600b65476c685f2521b813a3fb95f31f3a6febf96062de7e01a59f659f22cfc2d3d4a74593241aa4e691f7804e2c4b68831f13776cd6323a765acf4b5aefd1fda704c1870774a4ef7a8b468c8acaca4cec3aa26;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34ef7273e039bab258e24ee7ddebd9901f670cb383543e165374e95bfa591a9766d602a83cd9b5d74ea7fbd6bad244586877117ec6c438bd9442b8df4a62b27831ac36bdf829d2818c63d4f8f7e6b28c243a381915b447beabe4ebeb07f4f959c397;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd249743e4d322b6cb8954183c0732f386f9db18d0c18aee1f31e223d6fe5c326bc5594b25f7bcec816bc472828c97918ec9cb4bc9186df6570d7816f7a487c0d14294a056908a4967f931d52703a0489c6c6653650a741140b782f07b3120a947393;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb53308f5ead64b2bd4a2e7ea3f7d9cc0aaae96d57d807ddc32602f004e58380a1a1c4a77f6f96b26afb3b7fa9e5d454dc599b92ab700d01e60ef103beac8b2c9e7ab53a37c49acb8bc79f95377ea1216d51956a43ae40579b46da46b71728d9d72d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95e22ab37c8e536551a9949eec8e3acf8a8184ef84dc00fa1200bf0b968bd1602be07c7335212ecce07f69ac273ee31567301d39a92879266308197930b91ab30114df317cc4941ef4b0b469834015c2bd2f7915f749560818d1228a4dd177226d5b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h779165a1280dfceb1e156a9a8830cf17e8390c18a48332f90970598780273d7b8de2649f3a0643fdcf49dcb3f0fc4a4f69009545b02f322944c020a9ad35020017fae9b2baf6b5155722fa19c6c0ded4fe761b6b43b64d46afd053ab7dce5fc864e7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7e037a07dd1352ad1ebce623cd1feb13de6f5d9a5b85290cc628e0793ae015d8eb3b473ff187e23ef33e90ddebb112d809267513488d8accec1d0dc0af88599d8e265d018c9d48e92b7a7c3fe03d4fac4badb0b384a57d9392d27f010f0599a9d6b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca43325d614cf8322b270f0729f3b21aa775586d8757a8cf1b5bb36675264e0477e1834e7e9af775e2d14c1c1f0943c6660dbf3b5ea697bce933d1c566cc9beff29eabd7eba1033b6b0a2b3abf8bb220dd5de248b4a7b0b0c31040a5183a0fcbcd1f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h435fa672f4f4486fefa4792d028bb1685b657d906ea14884f5ae68b3efd7d63d93c2a6e26056c9f36f6d5b2c639ff5cc58202010b5539d4106dedc33e4a705409793218a75ccc95b9b21e194f0ab59a92fb9b262fabb89b2a15976371d52e292352c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe92d898bb5414dea36dcc6d254c8fb5fa9cb0fafd238118777ad0b15aaacbfcfc34f7cc83cfd8a446229f4ffc2f9b9c52faea9276800c4d4bbcd431c6a77dd5709c78848e0fcb13305a1020b0c0b88ea52935c6d4a304653b2ff0edc3b91806399b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he924268466877c9360eb9d469bf4db50c86425ac07afb0bd671eccd14acb575a98f977fa55e85f88c82e5c674b7428b6d6c6075e1ec6f3804db052b4dff0dbbf77d0827190636ba53c6af96b5fe608a411fa7dfbe7193fcb1cf23c27d930fcc4db48;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb6677572820d395a5a0a2b4eb982af33fee1317214c4bf010f7cc4f2b857c69197245b99057d7697caebc1a21afcdfa2011f869732fbae2aec343aa3518b3c3efbddb85fbff907fe74735a1c429fb913c104a7948282b990d40b39792894da3eb7e5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha625485f2ace9f7fa48cab77c7065b5d2e753238bd953d21a11918c09cb731d5b58544a4f5102de701c28f699d3576bc87709e34544423dc6fa737d44ede7953c2c644e78cbe1b21d0b7c05fa0e8deffebf9e31b86d3ee2ffee560eab1e13f1f38c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h837db8e347ed101921f4f7b0ab7772552e7c3150e037c114ad9a846719a462947444dc9561ffc2181c1e19ba4975570a44c4752fa3a95c9ce83b75b963dd19a90643d1952d74cea595a514f2281a85db3d8fb65269b88dc06878169f299c4d805e4d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h880a1d8b60eca05b2670b7e8ea9961f8aae64c5b9be10ddf836f5d96e306d56991e8e8e5a35d3b979afdb3f481e6b78b32c6f0d90a3708071d669f16b659eb19446b0eabca25f4f287660adc9b9142d5fb56115a52737f9f290e1660752a5fbb7253;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5acb90b6d7ba8baaff93e2db00f17828c08fccfac07c151f3c64ac4ce5ad1273d4ffbf67a7486284da686c9748d76489fb373ee5567ea4ff0b7b2fed220f8a45b5e41b66e332358dc2c5a7d7974154d40deaec932fbecb3902bab141dc2f5951da6d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ce050e163533c223a3ae5c038a66005e65c3fbf2ef24328efafb3ff78b19258c23d4bbaa7b884a6622eb81fec6fa5d98e229a3dd16b56d2485a3a7e7864ed4fb5a3d9ed017b74d1f33140a5bfd12ffd503ed6c23ce57919cfea9c534278ceebc742;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15b0349999862f10f3221ae5e8b09e2c30640caebab643c4a375d895dc1b2a8c5261ac2e41e371178ffedd41d081343ad7aaa343c2d2cc1eae8624ac1ab90b766dd138bf542afe79798ecfc357a33297e6c721020507881868ed6fdadb4f8f00ac2a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc9ea6cef38927ba8ce0521a1e21a54e309fab2090526d1607c7c7ebd7a2dae63c24ac61f49fe5dd84815abeeedbe8b1c0ad5b0577ab0a4f9040d3d67ad396ddff8328b6d7a2f12814eb49d4ec9354c9ea3625a4104360572d8d223f9c9185d33e34;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32c6e2a098dd74dcd8664479baa4a5f52e50f72c24690eec87b626fd7171af526310f15d3aac46cae43cdf492d5bc787c4df416ffe093d0e232c1b10c83c164895b18a479b0828904411a328e4a393c3c440c7fa101c337d53c41865065a4875b314;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c4dbabed14f2edcbc0c41fcf077e4b0751092cbd25160486f1c039a9d1ea2a5364d8d72c5aa53fb9891382ac4a56217b1f6326b615479d546a9584ae2bc1fcdad036da8ba35c43af70dbf98be64505c2638cff134e09c1fca3dd65a74c7fb344ff7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf11fa54f5ff170ba37dbf3f5b3bd99a13a41814b28d9373b9f5593a0b73b4e160f94eb5cab61571022dae9652a481af7edb02d2c213421618f2625eb109fd471ac353fa0af93280f793711f2e56eb9f61f336e8a14e1db03cfc77f168f88c5cd38fb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43cf623cbdc4471388f6ec0c39e7952944a0bdce2a7c85b519f74446feb3bda5730c4838bf141f888b945de2e0687ec97005b4834eb746a0340a5e0e7fcfdcafd13f2026d288167d6b0c2af28e7c9ec5241d737dc0a4679454a7dfff1219b53caa09;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h563d4c1b0a198d5210fe98cae5c63f9f08222e4aa64689c68348ecf495950cfa25ba061427bba26f8cf1dae58dd1c414dfd2715be2aa6a61a63a7fd36b25d5565e8f7096a19ecd7d7d9d2e11b5e1c4855cf7d80e8079f9f995e9c927bc46da4865c8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75a09168d1de484824f76d5f37355fddcb9b3e19567274ff25cac24918d3a8a888129c1869d158e347037bc48cf63f04a9f289497b9d1ecd24b475b2917d9e8bac660869513b78a88ca63fef43d67b88976c62309a25fabea1b36a39cd5490d21457;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8cf6f3c0642c396617879608c127c55232fe6ad2ba9bfa383696696d2cf9fcda7d26107e6211f326a807ec3a123d3f92180a2215238443f39feb4c6b2e6ab993af3027cfebe36d9e65d63fa93b5988efbd7f6a4d6066bf7f3aa5daa0291887b532cb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27ee9dae0852d810fae837ddb7be8d71436a87d36ce90c1b8ab92cdc50ba8eba717c7e8db4f644a2dd4d873aa0d90bccbf2253b25fc37e23d920052ea473e9cd8b9db80c5f95f2536aa5f09b431e0367f88751f79402028b4f7670e862ecb1de0b4c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25f241754b5d0ecf02badcf143ccc3950267a8ea6403c04410a808fdd605ae478437eea4d5956cfbdf504a3b4fd8c465312e4f4331e0f0083a570b70c32a1491fa982d54245198fff612f44d4857e6d6ff30d9debc7597872e1fb4769e1a0b7001df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had6e0ee3b85fee2aca2a2735a31e8caa1619aaa98c4b27a18d0cbf8afb3a1a228dbd3ec86de31a095a613cdded225cc1cbdd65d8739975d7f3d449c183c090fa3b8e79ec084707367a49dddb465917097dae8cb6c802983a0577878a113567810498;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5809ce0267e149bad9db3c43cea28a04299e2f1ce4bf7d51f5eb99b839ad93579edaf4ec266d914633b1477694dfebd5c3d04f149ac63c4ea60eb81d24229dea512b14991f06c7b64eb32352886f205ed4345496992f84ea8c9e79241e3dffa901b0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2ebe2a625992a7c06ced70beddfb5acc52f1b0536a075f5c7214b9e8df97e782960d39bb6dcff88fc408d15f62b04ab22efd1312d7892cc30aa2202644c717e510ff499fa9b761c0791f7f42a33bf4af7c132bdc6cfe65620f79baf32b870a0cb1d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4335863925e7c2502efca6a5c8eb9cde644e9986ab35dc62a02afe10618123e3b680565f83d042ed794967bbf17bfc239d2f1eced5995270b153ff751e911f2069b072817725994cd8edc3909aaa4bd4519ddff168ff5e9d12399fdb043372b53e1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac523b24d91ebbc585af1c29c8b4dd0676b515c478be1bf60f1550f719f9288d53aec3c461bccf8b81506fdb385112884cac51f78965d0587a15502c1de59039b9401de72b985e37723c26a19b54352d3ef39a2112074c5db1eba0230005f4f0307;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bfd5c4650c1b565ecaff0f92e41d3c0815ae26318be0d67f75921bb5ddc2feed9b4c045cbf0b3fb4c7f3fef584b2ee0f2eec2c31a577fe90ab0bc458c2751d60c71f5e3a375195f0a4051a4fe7957a2ea1811f653e97087dc7d30228974e3e6822b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38ca497150bdd774cae5331b8ca98d3761978e73efe79a17840c66263907fd964d66a4c590a8c333ac99cd826378f6da6fca136f30efe9679d9a6690ee0e3093f89190c95316f5edfc4b0ed0df85270a4e810c5c715837b5f1e9e383156a024a6a24;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35a982723f080c40d6f3a79e6b56be95ee2d74e693ec60b838dc8eb3c2d0e30d04682d57e928fe6ff54e486ad782621b00d9ad397314a0726a13ef1277bf4d5e80a76ef065d210c7ce6b7ab98198a059633c47d4b1492f4e23f7962aff68e2c05227;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h393d0bf93acca09512e065e95164792d91ae776af7b7765d1b39da1f9a69b62027990a54c1864e58ce0a38fba00dd2b860137f99a3bbb56a0a1eb901a1a9f5d49b6dbf0d64a4b38c5b3a5b96c87d271772e51ee1432714d034a7a009d8c0b80c7582;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1e98b0555d58ba97ce1d736e0623aa4ab0ac514cefe92e706cb23601410053e5807ca1506358560477cd74ee838e31968f622f00f8f3a810dca03fd54008f9d51eb01c8b630a710991ab39ff462782251090761b26fd8c96339dc461dc1af7e42f4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64e405bc1379fc1615387d33f34dc2bc6889a6a60709aab791b72edd8981b07699d98421c5692e8e02b4babae387a23c936b2586d20e8d799c6448fb79f3b1ce57664617392d25c6632bf1324b99b0690a1737921e015f3233bc99fe7a59c5438634;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f01528fa7859bc59ee1d6a1c84ac3cc0cdf6725be40eedf57c7db1c3a2ff0a718f782601bce80839d2e92b846355bd9c6d0122f3581c5c11689cd187d914b97bee2b288a30af97362194176af4e284fcbe89acddaab202c081f6abf01f9c825ca7;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2b95c601c4418bec9402d5c4947e92d7c3460bb1d7f3729b04f58979797fc130ea9d2d7fa4a36d90d49c2d4ad604cb40b4f2df06803c1a139f725c3b8a81c6d2f001d6156ed526348d618e3375cb66e76dd52fcd8072ff3e9847869b1d5ac039e1e2;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ad9b67cd05cb3a2b26c36897ab19f39b10710ba260c08b7b1a63c7deacf851166c31db93e2f1ad2b54bab0d307c7b526e0415c512273cad49e5488f9010655a8ef75baf69646307c536a702f19df6f931c7150fac4caece368321df7d072000df;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h735d124d5c8541b5ad2fec943f2bd2712bae059871787d39f9ec8791b69be7343052b5250af253ed06235d09aa61abc98c6dc0a35581899baaec2fe076334fef324c8f4e7fec02fa4a201c0282690b06bbc6266cf214bf617317ca4a257c89134983;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h637a82b06f47a6ec8d8620eedb547e8bfd8ce40e0b073b51f5542a2f1ab8e31f7cef9b22de7cd91a8e2c087e3878ea36dd41ddb07c39ad95aa447f82f4b486cb04b932eb3bb145d7bcf45d9c95264c5669419aabf9d99275a752e520a6af82b7a17d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h747c543b9e450eccbd9127ae726331e5eb92182b0e229528df12cb49cd52f6367592fd9869a80bbf7a05fd983d3dc660510ad0b6b498b9e6ab43a357b220c3617f16b5635105eb7ec34fd50d55a335f104b5dd62ccdf087e1b4b6126a1c85ae7963e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc08814dfab137dc97e0be3b0d175576a531380302e63922bf1015a060c158871d394f59b7a27caf3a0d6a1bfab2ba86ae6d02437b58852902f2ac5e73d90fcc9b1ef292fd1ccbc100661c04373acb7a9b6fc370cc8316d193fbaf5ca1c12de74aa12;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8f749c0be24f1c4725535c7f46ca0205f4e6659059f012eaf6a3aebeda86bf35d22b6951ff938869c883c32fd71e22ad1a3b05f1600d0e88969c7233f325dfbbb3b9ff3396e9c7091232044806cc14fab84d2bf74118527f734d3be126a317de40c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5dd3e1451ecbc8a7052bae698585893214681ca85879bef206d0b8ac3023018926ae728acb3af224515ebe6b4bc2b768f4bd362d3f171eb5ff5fccee38c8f7b1de903f8ad3c3eea39c3fef6d42cd998db2dad7c1ef5116c9a447f0078ecae214be16;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5351189320fe81f0d4a262f35a72c52cce39305b9e79b342466a1b72dc199e5d1041d5f5376d3509ad9ff12f462b7b085b2c26c02708b62e2c9ca3156746394ea4f39f9976c776ce1b77729439ba38e074725318525d26e545d590cd5b97f5590802;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57be44bb0fd3bd7d32c4f189598edca651d2cf06970de7a74f94ce4587ff2a869d8286d808c13128b3618d80cd851047e079d1d918faf0c43011d0698fa2fdf49d90044cca0072366bdb8c7ec763b09ad96b6d5320f20ae08090c4f8d1ff74b3b014;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94374db1586ff01fe4cadc34535c95a4ecada5aafa5484de298cccd86a4c5e3cbe61a8e5ccec9df48b67efd223cd91c85a22100ab2fb8b0e8c7a5bc628ff0092afdc759abb9ae72dc7180180dc3caf234b4ddbf7186d093d04e0f3d2037db9ce4bd3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a45a344328916e9b6535e29a666d6cc07404e7d2413cda4976c4167053212446f4b17532b2e7811911236317d77f530f6e890562e30471326f69f7a91bde9e013da2b0c5382389aa0c8c027d34cee8ceef2936652ebae025b1a51c12a1f9f17b19c;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he859007bd0ef42dc5ddfeaf34819f1292a8173a7bf5617abd6afa378f00a9c0c533d4c26d282b339b7af184a3d85ba774bf90d8fee4adebff463104473d2c10fd2823ff740c66dd0aab84ec180a5b0c7b18c2be130da93b219f88ab5d97b8daa77e1;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h523f8ff4263c5cf40f9cfc48e74ffad333b43d0856955abf0236823ed8e19d802bc1cb5705534237ca2cc797a220fbdcbc88d5132d740f6fbab1589636a7764fe0aeb78d2098c7ec192a90d94b3abefbb8f2d3f2a7d7b688513756094cc25725f8fa;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e502aa4c60f5499dd124a95bae2903b6a2dad7e4971a7144e3c0f3915e9f702ceaf731cebf0afede471fb760d6847547cbe3d9eba0bdef9b1a12b6cd5bf88e4c6729eb02776786d66d555ea9288dbdd957258d4985e379e12995369e694883b9498;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha154f59264b91da4fa60ecd70e5bf4a5875b160df1df2e60a717a8d73695f54caea3db49f10cf4ce5505602139223da1017025e1c022f2b1c21cc9bfa91bb15ee47b327eccbc205de7f2efa0bccc604de15e6bf80b86a076df3b758cb5f2c41079b9;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha262fa3febbefea77a7ffb394dbb20d8debe98760873cbaba365996f53ebf2e36a1753dfe009be5a6dc96b96bcde5d4fbf8c3cf0381c9376811fddf5103defc54b4454ac74b6b81145231608776aa49cf2f08aa059a47c10d176a5c77d6bad3682b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd1201242e42606619e2ef0f7bbbacc78eb16443a43392af4d4312f26207dd7107985430c263163726239875bd7938a7befc1ca2ed4c07733f897e0d81b4f603d315eac236267d81ac153b3c4c088fa599e024dd5fecdafdaed6c4ce3cc2d8d4cae0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ca0b6d6a44d2064a91413fe7ee0992ec90834ac7b500b1e36c85b50c3ff3695b033f2c2b68081336d44f040b042334eb68129627c54d82c1e8c423b924e203d1be835a518f7b57c6d2a8de8ec2915e49555d5d0d97e1e63b65b83f1639d617a30ee;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5cfecd286d3fef0cebf7bbaa2d2fefc94ba2e60f87af9902b663d57c6950728644542ca0b4d7c6ceab4874c921658f794de50125bc23c8c68c4acbf21be6b5e1e5e38bb17e8e9b64bc6d60fc2a2ca85402d46ed2f2b4e1ff85363c8106d91d2a7ae;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce604985a3b5bfc4d6241359e9fd732172d12c42cfcd773e16b7802f982d361fc014f57aa97048bea78da799c011e8c5d60f9de13a6954bcb61ebaf691a3e295f6eef9f1ec6be0a4712ac4c570d10e55897973bd88a566199905ae58df1b666c18b5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha851ff2837c03fd5446b8561eedf871207c3be62d9c4b106eaf513ec2363edefd4410e5fe4d1d4f46b83dfc38dd58cfad8456a9ff4e9dc7957b54b0bf0413ddc0c00f05b4c99a10f3a5363865ba3aa2b8081e94e95a4c2f6e1cd2deb3c60f3c27695;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc80d8e6b0640febc2564b0c186b49441f5383f95a80f4652101c3df12e59c86688c28b531112142dc049a4480cec4c59384ac780f35f54eba18a332c9123c0f189baa55be1b2c2d31257a65b0ca9e2be97c10a534011af176ee57eaac2f41df8d97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h706e59cfd60996db4e46999478ed7545c98f07ce592cdb428cf8e5d98bcc0172d8f0d3cfb41bb063c0c189f8d098c69257eb3de2e80f9ed977eaced2cc765879f6c61248025ae40be5f7d7cff9c727734385bc5f50b7427d83910f079f260b5d56d5;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h461bde19880f331a7a003e7181a22f1b3b60381cd6851abbaa52a1aed9e223f971ab43f4cdef6bf55f5a57e06857b814597f3e0a3f00ef16731756ea2d47ea8b1172593eb95695334cc0b89d3862d085ea2cd7ba4a5b2f57bcb2627c6cbedbe2b13f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39b972b30b8d480058b9e3463ea5c2d12f02327b44f45febbaf007ab43ecee06757db7baa06abaf70e5a01d604b88e140fc5db849aa3733ee314d51f4e4d9fdee8c03ebc56413836a541f72ca5fabecdcdefe7b9b1f5076b9fda0c7df9de14d72094;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd50c22ef9548d801c0c86646de002754563840f616e390d91c49dfbeb7e94acd8c7ed8ed2c7d5e1290a53edb16ebc1305cab1a43e0030003d3ab336183e15409b6f984f157a3a820faf7fd92228f29e2d9d07a7b6f65a9047ccaadf89a92f68b07de;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca6d34b90677ef535ae00e7ce6333f4a7a1e9370f9a193e372ce70641428055df95e57bd703bbe96f4041f2a3adee61a2f479934c15822a8f81ac29c7c649bed2a57c108cfcae942519c7717979bb7e0849dfd056706dd80b5d03bddafca5450e930;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2eb89695707bff7eab83c326e355ef7666f58dd93e6e10bd06c6d69f6ac77879c134750ee888abcd51673c916d0151bf389f9e6454ba9e343d9b993ab88ec3ec6c39080e9ab686106e60bed62a043fa644546225ed6a2f472617baea0e0970368e69;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha71e5d7d2fd0cae15f3953b4e97ade3d2f87cd439d6554659c3463d18faa9ab17cf4f63f2b2ea3b05100a622f7e06a58ad847b7867a21f946c82fdc5feae1c70b9077141578b763495ec603dd25ab9295e3071955336dd9ce5684821ea5ad5ccd33a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42259eb9a64afd1ff333866fc7c4d25847ce1feb5e98103edf1fa707fc826dd5133e056ae00c17beb43642b3ebaee80edb0a8a825d8c3c971cd8e1febcdfe80b8cf15319dc8c47b7c58bede429014799f244807bf06e460a3b296e3e73ad80dde7be;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16891ea73c38be5ecc4036b2a3ce2bcd05a723ffc2f39b7bf2b60a79573050c2b0d632147f6cf03365784e4d3619e9083c88fdd2c390a805d77e1fffc2e9ae067031a43194877065ef5f231c91fa4708c56998edeffca8a2c911988429cd2c398aeb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h486c9ec9f3b27e20ebe42754861e762db884a14f876a385cfabe53a472b5cb5a95af40403e752f4efa9d74fa80fbe140a122641e520e296337c02d2aca71ee5a504a92cd1998526387e89ca880ad2c48d312db922128b7787bdee7469d985d1463ea;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90419de55601ef8b4a20b1388c9822c1d1dc9caec126329ba276ddf4455b646baa65b94e00aa41f0ceac341ca7e1df5985831ae2810bdf1b76bd894bdab241e8daf0b16411a75d3906ad6df223a7708c0c5c40b233a5877a542e7697388c99a6033f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55738e9a0cc208a3271374a33ce93bcbfc48785e80480a43999732414fa1f9380362f2d8c76eed40ad199d41cea2dd8fc3862ff2f32ed11679291268f351b84a12e58d782b296fb12fab3ce6138242127e6e7774ad0f327be228fb67ecf636790de3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37138cdbf29c08da355c9539992c690f47fdfec5474b8422c3ef73bfcfb95f0fc4bbccf15676fa67838cb810d7378e8674bd84a882d3fbf66c1e2b5d8d897032dc2f2bd743ee952ccb650f9621e58b60803f4d572a192ceb502483ae3cd82aa78240;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5008bc00af12c6a01a710cd6e6c19ba70dea9cf38bfffcb9fccd180464a5348c17138cb5866c2d248e98259268641177079fbaa1988400040ce02ba7da4a6b0699583372aa652cbb32c69eb303acd142b7964c8ed841627da2760c1de8591712c7f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cdcf065c9b8415a55076d9c8d150bd738db614efbdb54bc8e26fb48661d12c4a85778de280db3670b178e46bdb3c86869c295f54ced18e408e855a6f681439a64a187ad7c1e2a21e52ea98b778397bd58d55ba84bb2440d4b4dae62513ce51169e0;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ec3cbfd5d0f9bed8b6b8263729238aa14ab5ba006c5a1d86c52e58aa49e0943a5c1f2050f807e73882435b58f8dee7a4e14fa853529b02ce2b8b0bde0e14de84904b2fedefb433aa5610c20f2756fbe0297c48e833d4de2a544ba7e89964b174838;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h396c058b2162c470c6961d18e23bd868227d0cad3e3f4f8499d4c9787807d9f1f3f6ca0280d5a157132c2c1f2bee8e0534941a6923b985ed2b18767c353aa8a5887471be5e09a3b1248f0b89ca83ddcb101c2b97c6bc236f248f718f585a79ecd157;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a9c5c5fbfde5ced09598ce06b06469c4759a91110891a4696b49c2d06f365ad9efca3e1b2469adcd363348ea5431d7222ca0986b076783961cf93f85e0e3328c805d9aa6c19ed900a199d94592ec5f30f93a95902801c445f4240375daa70b63e97;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ee22ae53bbb8b19645171ea5a2e8bea7448850df07d5dd01aa0e97b104de3d0234ca2bdc99cc43aa0a2d94a3ea628f5f15dc3daecc00a7393b045150a613700c6d1777f19ecc380fc207fec9f185f82ad5caf6ccd44e33fb2682130e18e6c9c3598;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76c51be4e9026186ac77dcc66e8e6ef85da8621900598455ffa4b01c253cfeab4999d737190e731eaf129a7b21bab0b5b6352c811435c075f199b6b4521bd629fc3da7ff83bb2793865ec74268b8433beb88437131f0db54324bfe2628191c8b2f85;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97b731b3f595451abafdaa1540ab5c8285232a3aac51f36378536f04c5cec965fed6f399f6f6e8f7b3c112af4339f86e9ccedb8ad9ad391ed9870b868e5ebfbbaf15f349334e761dc6d170519e487e3ea4176e6094e614b8e27d25152600438d3d2b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b58e15623869c4addd7ac94a4160a13b7febc9ab106226b1c991cf1c537f759e6d998b2f7261d4f3d274d228aba65bf1b12f59ab6c633a2bd2240e0ee120ec738a998ec118af774875e56c169047e2fb6763803b4d1940239bcd46dfdd9da6501f8;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19b82509efae50ea150430be9ca146632c34f9d202eb1f1d5ca88caf281692c419805eaa71cc997ddc1c1857fb432ffca88f803cb614e5cf8a82cbe3581518d2812bb5ee91488916102494fd978ee5a8e7464431da440fb7c139ab77d46fdde4a85b;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fc97262455f981b9c33f9663c04e1a5d16af3906198b2018f045f84cb2199feba5b93d822311c143fec97cdfbebc82cc406e5820e67a7639bbcb43b2aac25212aae546f046ea4de9bfee734d688ca6d5e3e419a465c2af2a9900af82cb9fc116fdf;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5d15637f29793106d582a88cbe324e030f671d5c3cf9266db58ce61f76041308e2ae0e6d93aa374bc049ddf87ffb01c270e6161a6e49f0c004843413bd8fe56cfe4a901407f104b8a1335c7f20464c1406bd9a79e881de2e9163d5a7442ee769d1a;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c5dd1e92e03497b483c60cb1de9b571124bd6083729f378320cc5f54fd1150a463cf40e69298db7a3cfc467661cde32fd228599827ce391e0ce604cb202daf326c0d03ab6d6a7e583bf1f7f51bcdf1455d3c9f0f823398e36f7f535ecb889d6d41e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h269336c52a71092bc97d385929d47c20be45aedfc8aac16e2991bf505346fe28817ff7fd9968b9cd98eb70b112f1e20e05fadbd64bc460fbe13a5e37c76563d7c2ccb005f3e2d1972c51b38d7a7b043546e48b0f3ed821f932e1f9b420ad1cdc2480;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba08ea8ac632ea921f8ee5aa1eb25eac9887880a05e0671b058ca9e9b802a163e804eee63a22fa41e255819c286016afbbac255b7a8d97895c6ca2009a5494d0e3de857e028d69311f34004cd44f06fc67c7c1aa9c331e5c0cd45c488360775eac7f;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4402b83453de03359e0ebfc230adde8001ba86af920bcf746589c6be77c4a10935cae79389d2cf32960b87f6eb10efda7731e6a70b8c46ae39d8416e266806159a8f73732198d6a4a732f30d7a38e1d645f8d299f4df8695ea268fea5d397350615;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3aa02e8adaae2b7e0225a952f339aa57c0f1a675796604a33f96a0b41934af725143cffa52f34d9053aea23602fcdfaa36d3aa7d138d50f0b7bc0a9ba61abb0b549060c5545aca940cc4265d41167310403ee372527cccc5a2060cb4d08b9eaba3a4;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h318be0cb746f1dd234bef9ffe03f8bd1b79906f4fdc827e5cdd30d60f062bc113ca7525f3d19f2bac9b1a2ddf92692f2e30667142e402dc0015b24b944fe0d467bb3b4ef669c40331a0959472f9fac547d5753603bf451eb44d40908c4addf3e5f5e;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96b9c1192bf99fbddecbd9e7ef5783e81ab91ead60f70e0f7a50956a3a55dd43196223278c9e48543bebffba58da6dfd3b32bacaa82635a4f0fe6a7b8c1cf84a76ee474ed5ce930b3fc293052222f77c3f7f19c878ccfea9b780d560d6354b2e16d3;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ab92661c6ceb8959fa1629a6bbb581e14887866b83ccc4dbe15213ba21ada38e84ce29cf25f3bbeb1d3c4f5f52f7d51d2e59c907ff83f5fee6dc56114ea35ac7de780906bae2ccd7dfdea091e2a7b7b9ab02152cae47d6f239258d8469806eb564d;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3dfbfa610601b6df919dad14d72fd8d5e56bd287f4ce6ccb0ee1e0e2a68d9ac95b999666475c2a47300af9b411c9efa8894cdb0880b5ce0712f5792b3455bafa948d3682e00c5cc11db2226a60b6fd2219e4387b7f3f05ac1728206591fc45c5905;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7fbbba6f6a61a752d3b69eb982f2385ba61ebf5cf7b41afc9321b12f979c335f5309a9cd3a2733a2925c9cb538ad73e096e9f9f643d48b9333313bb0689bd0a5c300b54d6308d6b1ba6248a5bfd4e413342b47d8910aa9311e2a928cfb3dc59c1239;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb53f3306271c5639cdb09cc24e35a9e9889d26b9cf8ba3b8fc8e339f34a59576309c49bf2b29b90ad736905f8c6faf8413df9b661402eba2b1361d73d8ea304776a709d73c1a044a48449e969d3d89c968875a8548183ffbc4a5d3710924428bd43;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66b445d881806723a7785bb7f14b36bc7e03adb632e28fc92bad4531fde3cd39f50193daed5aaa5fc284954835a03eaa28da3c3f3d2b1bceeaeba71b83ba095d25ba5eb338303995517348978f4b3b60b6db7f49dcb055fab665b8aee037d23b2bb;
        #1
        {src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he9329c786cf408c3b0d69f3ff58137c59e7c1e787660e15ceb4090c97e924bd6a4974834895829bad5137cd268ac0f921649b1d97dca468d15db550df77b21396f486fc2dd312d2dd3e681eb4249f539854f24fbffad06d90a33b600143339689f3d;
        #1
        $finish();
    end
endmodule
