module testbench();
    reg [20:0] src0;
    reg [20:0] src1;
    reg [20:0] src2;
    reg [20:0] src3;
    reg [20:0] src4;
    reg [20:0] src5;
    reg [20:0] src6;
    reg [20:0] src7;
    reg [20:0] src8;
    reg [20:0] src9;
    reg [20:0] src10;
    reg [20:0] src11;
    reg [20:0] src12;
    reg [20:0] src13;
    reg [20:0] src14;
    reg [20:0] src15;
    reg [20:0] src16;
    reg [20:0] src17;
    reg [20:0] src18;
    reg [20:0] src19;
    reg [20:0] src20;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [25:0] srcsum;
    wire [25:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ee695b2dc72ea9944f1ce37a33bd0340d2b1fc4c6c6c56b0bba96b585b41a37c23e9cbfa800b446df92ab52b4a047548be3a87d20ab626;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17511fd786a1452809c39bfa842a95540c92efa42e967b95f2d3c6ae5a4e0f98d2b5a163f6bd4f8eb2e797e0cee9c7aa98351f82a576569;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a8ae888b8a678add7aa194bfe8fd13c4c9cd4a5ec8d16f1b44ceb6dca90e3ddbbfe62393ed504765620a7fc3b1d81f90a031990d17519;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb51cd27cd962255a69930e4d82c6d412b0fdc25643ed29eb11b8d72afeacc0a6fef14ed99bfb82b2f8fc60b0c6769ab9695e3d6720d97d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc75b45cdee34404365abe0ab9eeffb138bb542c77af81dcb791a353e4a94b09b0eacc3901b565e3b25592bd055896b2662c63578341910;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12aaad40d740d79558b3ba5dc8489be291d39dd22a0c1dd659cc6769cda3fc130205ca3c32ee149b68725f18eff0f69bec0e191dace0c37;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8dcab8acee067218dfb14cbdb37b222a4beaacaf36b3b4294b33a9a02d0b2ca1800534dafafa7151b3c7933da9ab884630f35669c3987;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c8bb4110f7f372e42b525aafd5bd0e2344597f33efafb994afc1f6d3550a50aef7efa4a5b22e2d569bcf36bc13bdd0a06aebab4a414fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h543b838da05ed42efc57c539a20ef594a9031b467954402000ddbeddda949d68ad2f5a5bee9c13a155154cdf12a0b4f69bfca2c378f350;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f2fd3c421c894c80c16e37e5ae6546a4eff1e00c74d394047d25ae62700940000e29b7b60ab144b13d869133e4325fa91bf2574e31e07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10863917696e66aa7d89399d226e1de6970597533be32b6347e6360e0a91920b4e003fba3f5ba664983d16c889de73d35b533d976c3b751;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h124430d20f24f62da2efa1303f62e7f7c1ecba4dce99d9e304cf7f73d8195565bb74ec0bbe0a67a1570f1c62df9eaf8c0c399d0fd2ae6ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2850732fce73a46b3d999ceb2d9a9bfbd08853dc80870abb2a58aada295faed97dadf143b98d0e9aa52fd3b805aea28cccad8ca90445e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbca826275d772e69f90c66b55055fe0256ed60fef0d8dbb36bb2b47108150dad5287a1baebfce8a7e4087405ad4c7a1bd2d2bb6efeb907;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h192ef8c9f625cbb3512ddb7bca4fb2daeb63d081f8a5f76bdf0e97c07157c6423d52cdd4cad5ac0d13305c655bec02411cdb91073950daa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd43abdcb8821ca21d898db0100cdc5e93782f96289d13209d7b2d9b2c482be6f4bc04980b21c8a776ef77b16be5f6eec1beba85003987;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198e63b5a64b791089f1d841ace166d03ad0d689c68b4f15447fa03954f34b82afe72266cdb1587e5978d12e6da2b3af965afc7d6f4e164;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9a99c985aea922ba25901893b15661129bcac3232311c8dc3ff6362990719fb210a2dbc8e9cc734c31a4d0f8920a70626dc494254b6f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7295f348e9dfbb9aed079cbd0f819a18e73794484c99fa2f7a9c059b843228a9a67071d8529d7c111580d899b1d96fd03a0e9370f0725c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b787b19ca6a18b22f57aede62055fbbb0659bf53dc53b619b8ff31bbb3edf24fb20826e6b811be71a26e8b2ad7ae48e510feff5a18f78a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9176d6d4bc1d0b5d312f6759247454caa0281b40ad491c36eb44dd9c3f7bb3c898d26f38f3764c6dc7bc49db4457ec26f6412ce4b3ae5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1685138b37a18dba07f9594d2d6c87845a3642ec305be58b49a7cf3f6b44fe7afb5eda85ca434e58ba921bdaa6a619d9978317277d04f64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca69a2e847a90ce2968195a83624fcb34615c2b4bd86a2e290c0a8d42c40138e11a544c80ce26ae86fffc3ea21964d3f1bdc87e5e891f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd805ff2ebebeb17f4c6a720754ee20d0b4df55e47f191437b221483e68e82592bdb2d67c4dd41c80be168c92cb1773cb64916eff889852;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1857364b6466063df5d7b925f40ce121db50ee0c54f187fb82afc0273135d73d285c0c1ed639f77562c515535aadbb079b53ba6e4f2d3b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19320b8a31ee04ca1238fabe34fd55c533fcf2aeec8aa692d9d90bee53b19e423a26415c0db3d74645c419ea1c5c15f180c4a91ef895a34;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h76b14137f495f44522359502776ceeef11b5b5ace0c1f2edab76c0a31c2a244ef6dd7edd3565b510eaf1d02e0ddcc91e1e200273b92e12;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a9b2d7fa1e7fe5ad31bdc0ea9fff65be70abd2f7fd0d8a313366f2c0ead85d224b4713e0836c8ed4ca2c92ac547d1b5957db161af22644;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17b81e743aa41a85db6636068b6cd97aa6f564cbfcce17fb059f9856d2954f862e6ebef33cd87b74c0cf518115db2c50e26a57e97c9c85f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1deef02756d77a6e88d1c5b66462efd9e1c1afb1d3d5b6d3e023aae65932e971e93f9860755cb3acd266826d1217f8076ff4dc04e437c7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf3f36c0bc0f51a26d4f1cc13cd371abad4c900146013dbbeaa91a8df59229f2b24fe6268b9df4ae3ccb65647ff4f820cb272d0169f486;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc77394621bd19b67edd5ef90ac82e5c63d2795768843c462c7e4bdc6a092c473cafea3dcac7c4edd272e967d3d3d8ca3a513c0ea5f980;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a999093c81ed4fe6dbba49db12b6a252823542e4d71c363b88995503d21c78bd55e71975f8cb39ae2f85df53898f66ac4053197f3a856;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef2d9e806f152243f1541784c228636ebfe159a824c7d6764ad5eb33993edf24ccacdfaf3fdd5a878343b5b2733bdad871e1033484c723;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc7dcd4cdff160f38be29e1ce174b95aaa306261b96a7933e64583fc72746a79e26bf5001c81f40976af922ffe303ecd71adbd998259;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4846b343d997e9f9df02e1237a5c1bf74a4c781d0d7f5259d5caedb5af985c474c94cd7115509ee6e942342e451b57fe6ca11a27e547f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde8d0adbb905dd806d4925c7b5b27f4cfe8ea47e02bc58b3ae8cc560a01d0dbe3c4f909544b45bb0fc8e81e6e6dc5e2122456b029493ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb662faf3000bdd70f01d18e1b62994f18c81573506e557882df8eac540363eb5cdd4a5fd520e24c0d0c872907503b393bf8f9933969145;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188dfd64ed241f1379b26f6535b133c1971903c26e90d23c060e728d6b44eef49c07a4f5f88adbd500dd1613378722c795ffdb0c64c49c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14fae0a388b2363ec58129a7aae1d843b2d7d57f0b214811f68eed098ae09a64fc022b542b65f92f1db0c827c854581524d2efb27880caa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a0b73ea91ea07be6d3812e6bda583a30c2fd2a033fcdd294cec1abce4d933d61437140d75d0c20f6f006097273fa4b5da52264e53b887e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h53b9923320cb3284981901447d505d8657b031478e9b060fa05a72d8490a9172009e0943adb1302c72c9da2782580af84d8970d27349a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18109aa02a1f0c8c6e03392723a8f74ff9be45e8fcb2a9b6abd56ee8ab3c02660cb68e98f8a6b0b206d442e8a0639522ae0335e1ce2978e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ecb1610387ac29ce224342c16176ee89aa27357ddf1e02b47492faca956496d064f47313a69f6fa0125aa897057e74cacbbd163b5a8ea6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7e582a8a29ff692ac532caaeb63aa226f6c8f582d182f8659688e47abe1ef0ef1bacf54b05d03477bb0ded75b1e47023ec7a95d41fd132;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf95d99f29aa432242dc0358084a3445a1b85c755ab2096fe4a4c9128a23d829b1c7c5b3256a7f9d1fdd922ea7b8073fefd5dcd894c5c75;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1108be0895d9188df9b57692ece144f78314aadb1ee95508646ec0f0fa6d72ca7c80c70c87ae9abf93f945c89f2eccc72726b7ff34598b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a2ef67daaacfb245cd2fc141f4f0c4f1333aec0607bc3b8ea65707d3d67f2e298b56acde024fcc7736c1e9ded07edc64ed7eb863cff9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15710150fbfd77c9a912f8938d2080d3f19ca04f4ea206149e23709238d80c3afbacefe44b6a2432d51359e9b743a3d3f5210b810420bd3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17e2e688d842fa0317024226fbe8e9a559efbc03a5452794b4e825eb8bdb3e2298947dbaad770dfa700a8d304a3bacf4475ddd4c01486a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1962a00427c3577793656b6a6d27b43e0e86658913edc6daaba35e796dfeed826cca3ac0cb9b1f9169e2216803cefa7b8369c630d7fca2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1368e58d46d4ab436d76fba7170b385fc39f6854b92e469a31bde7866043db2685466e7037a0138d91474bfa0ad2f523de7d36cdebb78a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1651057cb5385ce716c228525c0f97fcfe4dfb01e7518be917d33fea16072e48a3f4ce5373458e94afcca95320b18ceb3cd5b8fc1a0fc1c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b64bacf75d1afac7d5f69353a4b2e31f56162f3b131338f6bd4ae47dea874889cb56bcb2b031fe4f70eca15e13bb8c63aa29560612298e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e67006b45d3b078a78a178119b4e7e3e13c14730fce392df1f236275c3e22805d8e06b50d79369f7e7f1a9dcbf7d9a4bc2ad6caa7eb983;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h406b77a0bae1ae9f573fd8a0780b15f45a5d1c24bb3e58f57035d097fe708dcd89764a2bdec17bf31fe717e37e2631e78760d51df4d35c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac49c5f3b169a41c99b2c6e16c1c275226edfb246da3f8e13c65a62b82679dc80a8f4a70a69209eee34ccd5f3ab7d78fa060dcf56abf26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11aafa0cc1b86bfe6adee0573d69f5b1307954de0f60c70df5278820088870c2ea11bc8749b4d340e6be186ffbae934b1545c042a0a23d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11af1379c3df063833baf3500da8f8aa9d263f5171a66c910643580eee5a6903f41d99024b71aaa4c92a2c90b859de0eab34c0101a5ba43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b6f5cdbb5903fe38fea99613a1b4909980fd63433f1be9fc052894d291e63dfaed6aff003820e45ebcf52139c0931dfc844cacd9c492a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h146509ee50996590734ad7bb08a3106f0e33b777be00ad877ad135fe76559b94882db9fdfcf1b0f5d4cccd7111f7480537efc6c71e3111d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3afc2910d318f515bcdb7781226773701b7558346b4dffe905fbfdb8bd09694dd4e1d99545f2a2a2b959c425fc39ab2bc64a7b23caf322;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b05391ca2ed316a20b708db81e0f62d1cedfdb1182d67bbefe50fa3fbe6f6016fc853e82ddaaf8198fb0178b287365f28692f7646b9631;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129508d52355f0ebb7879eb75627ffafe00996530d61d1b3b13db8e17420ee4d7cfd55676e9c9835534d84d18fe7c7ac3397f069b2a229d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a100a67f4b798aa85d81bfefcebe7bb35628b47721625f6090e32669b679b442f2ff0782912ecc9866c16c4aea80af739544979e3cf1d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha93917b99188aba304c4c5b42b501f23ba37b184360ca1d2b22f2e7ee8899c8e5a63bfc507aea94b3c7087a7825cac773fd49e29690aad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a0bd888fe96936da72ba3ceaed9462bfd4f450c8192a4f0ac4c87a2d5795db22fb64215509e4f75d4a8fe47f409f7ccb04f7b48257da8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bdabda94b9244d726675068cdc5a07e9d9fda9f6715371dc906fabb071bb7adfd44e9074d5b634717828af92d26c0df7aa52e482f4b643;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h72d15fb066850a6fa0ecf4399f647aaee195e617dda44d0b0d283af49dc4d5fd2a9f26bbe7c7b65dbf3a2d60369dd7ddaef5b8d947b85e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ed28bba422191d1682ccc84e3792b54d3b1624a3fa3c0d5322f23f8119768c1c623ce2fd596f27afeafd4ace9a6f4158f3d24b9b58144;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ceafcd32ce87e617fa1a8acf0be9dc39969a35afe63608495143c1fd8737f44af9867bcd72459d4a57193eeb664d680febd9314d1f0c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he9d0717eb43b71c61286cf0e17c9e3570101ff39b9b1257d59435a4d5bb8502d2ee1912122e9910369a50942eba66653778925493a117f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117b75956fc28e41e818a2bf38732bd9ea7e9033a8cbe81d2dff3652506db732a105dca2e51f9d6e35bd03cc01bd9fd0710481a4b37dbd6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6865f51161943576640c80155eaab1e85dd21af4e58b2a572a96d28650c635178eb24157ae2bd053cbdfc7b4c70b7bf07c6fc7f1c73d16;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c0334dbf3314782f98c1c42ff301fea4b31b8fbdd236eb851c8936e094f714cee14f241cc6b29597c1dcf0c10f46aaac01cfa7ab151308;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5d48dc43e6172b21ff336b6b709eef9c5d8be99a3569cece55f8782bc8ad4fa284371938c52a945a62f79d27e10d50f2fc62448de4767d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h399c0b33269ec3e1cdd0846ed5a3ada60852dfd6e4b173f64995c7aa4b21465ef68fa1703b1155b2c1f063b4ffe8d8710e39b98693de1c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha426d856f2d7837af5709a91831fe6bad5b65ee3b4b543f6a01456f7d0f47db9fce1b196c6e7d7886f6774f05bafeaa6aee701cf700080;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfead43c8dda3c854cbc9ec24688ca2b91cc9116f0c492ed1920e824d08f3fd3ff01546a1ff49107f6c98ed298f69a0628612412d57c966;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1067ebd80b3e48eb956ec7ded09752ee4195bd2be46bc0a38974919e41aa9641cf786848e2006b80953fb38a54d48ff6d8180e2582a1e7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11656c730a24ae1f2acd3e0d50825252212227844b585930053661eb569f8fbce3bf404d4d9f2d7203cfee1c4fbf2cd3599966d7ea9fe6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10faf175695c707d477cfa2ff9ddd4942e4677d7650344f4d8bd9c294a18ff61a66e5c7eed9bef4bb0660a7f90d46a44f8ec9a8d7b28c0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15121d3fcc03ec115e0f9d4c8149c21df2ce19edec732ec3c2737179c9a12c2c55c7d5d6573ebde68804a940265c31cf41a124dd0f693e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdaef580b47cdded9155b443277be15ee957aec715949b3495e0ce8d40492f5c35285112b38cb160b1440bbbdb8473f7cdf7fa74cc9fbb8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79fffc0b6a090df2570c6a4fa2b839fb5c6685009518a2c5aed99785012359d5e2884cd3520b38168e9b299a15e60695d3ac93613e2612;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b784e7bebbc69554ba044b503a476aa1a6f13d747452512d325f3d260f8fb490ad05b53e44bc2bb9c528a3d33704c729a9d33824a96d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d075c6d626a422d82ccdff83610d9680c46af2bc1080c324a5ed13f3d272e72b42040c6a55e9ec2cd614853181bf885dd107a62feeb3f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0e23b7e12986d327bab588b65ede2b5cd4b7543ee6f0098d1e4b164f019b442a8fd0f447b2ec5f92dbb55a7268a1891eaed05f40f00e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h73d1fd44390309fe615be5bd2976b7145b4496d1335cac8bf875d65ed511b787307c1f52e631f7f1634789b7daa69a3ca8a7f39746bf6e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16934d0e2057ef717bed711aba1198238fc46b9827f2ef2eb1df1a58c339998b7604ec918ffc599e62f161a635163e2e8e83b976974f41d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164ea27a9c5696d3e452b62b54dd377ba777a6e446fcaf3d92bbed45b1b5af7872ff7b1a0c34a9a42e84cb50c02993ff18a48dfb1a485f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b6e711ac4273d272b48b8ee44a3082f07bc70fc185b5895aab665115047eb9fb222639a17b108793d96ad7bbab7b99f7abeab908b4325;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf40ee9e704bc689bc42cfc5a3ffb56e3fd08ecf7c3625777b2f6730fdae031deb3854a5270f5e6b449318bb488ccfd6337f8806cb09e65;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf91ea8dbe92c9c63a58fa0f7f30ecc7d9aa0661c78eebe7f05b86bef03213bbd5b295b5247e2ce62c5ae0589889835a69eebb7689e171b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a57acc4c49b1f4f5ef334bbcd87fae3e519ce28118f743c6083f3a161fa8b45f0cea24889fdcc2ab71345a80333f1cb215a7d4ef1f9a01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb82064084a3507e552248a2a4cad5a6673eb6516a467e54ff1343f5fcf6773dfce275422610ea2dcdfa5d6963acc688343c31d33d17d5f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d6e73fd46a79762abd58d8de5d471b8481784ed01e8dcdd98c644571b18c321916f5f83a8f4a0773830fec4aa189c13f54e7a4df4ab45;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf26c54f33b3918c0a93b6d380b9337e8d36a127db0b0e770d45c388f80da32e9a70f8cbf1c12f9506e70824899deade511b35a92355c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17fb355db80f1cf763ba01acd24d36450e0a22da3888dd131cd9db2283c7c9966af515d2b803c891c5140515141eecd0b47a9caed981a1c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a7adb0258f58ca1a115107a177e6c1a56c3c08d9a06e0b9d2549b7207c69e59d2d2353483d612b711ee440582193d70ac95f416e40c879;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h192b00a620c9d3a79a3fd8f1ac105c655be69ccd616960f195838f3fb7dfbf0c7bf944de2edfc481cee7e7627498c24b9caf03729124eba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3b53245f928c09d27240b700e31704a81515e2ad28725f1278729eb02c2ee154ae042e1f1e5f522a8b0a6a6ea95d1f09343116c03c47ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3944866c114c5dc0eea1c3f8ad7b1e4868615652bd7d40e41b361237a785e278a6bb108aed8aec40eb9dd221c82028cee841a03d412c76;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h90f20e9b59ebd4d9372ca6afd40185a024c42d0e6059d314ef1ca85715f4ed7a0e6203154bd0fa5888b6e27407ab18498683b181b11782;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bdb71a2eed7b6c08cf5e53171ff871227ffed42b08dcdd6c7ad0b539190b5e5235c033d46c171c1c0356522ea0a0a284f189cc5b91ff30;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5533d9873bfbb509d31dc57d1ca6ebc3e8359ab6ae8dab3f84f5f81ef56c960975b2fe69a070d23f0b22783402c9f2d843ae6176904198;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h112aebc3a60066c7bf0e02a6a4c90d7f41f1170d7e6d45bcc18be25460ef27b958ad80ac30e5e8a4dffc3f68289e50013c91e9246d59934;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h188bfbc7019690c08d833c99fc2107b20e520ee829586f0196db16e21be4344e5ce01d32a084dca108159f76bb50a4d3c7e8838d26587ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1116f424994caa57e2ec362983ae69f276b7f8d3232a160efc4ca699c71029ee5077f3463e361e101cd2bc111147852de023743c0133280;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h36c2d7d0968a134efa6dc613f642930c5a7acfb6f1bd61434effa99314f64bd4ff46f2b9a8ca1bd7e9cdc4553cec01d71cee3b2d0bb8fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12f50d1c30b68a4455ee8dd91122a9af2f93be55121624283d1029403c5b3a6c504f34c95563f8a5a3ea59aae465e9bed0752cbd5839abd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h658f98b962e274b17e46cfbee225a68530ed7c8afe762a5c97daf45978a3c91682e45c1e52a013a7a337cc7ba8e34d9193cd59e46470af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcaf2b2f9a1161bf91e1759c5620e07708a5cd1a786d20781195890f8dccc5f2b4af7ac369241302ec184d60a027d31f5325ca02b793271;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f881ca50dba8a4de3a015032e609ff2d87286c2eea596950f5fa0d687501d0bc68886f9ca412f546b1beb085847c71fd1479adc3ccf23b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c53047dd247111e4e717fe03f1b32e2dc99bfd9f0aa495a48559a597d70105159a162f5025908c4bc251f6a6cabaae02149a6a1af5489;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1979d99f500248da535319b141a0229fd17f9928a2fcbcce6f9b05a6fcae9e9f41c05c682b9510288a893c9af7a05d78e363cac6509a488;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h30e9c1edd9b1e7af53436ee31a79a9e20d1b43e33d65674757c84a1e6a385f6e3701b9de1841aea47bedd8aa01285c7472f3fb14611e88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h163badc0d32b41671ceb39cfafaff8b751e292f2341757d8c8ed3459ab39688e87cbbfbee87dd0091ed7820da61c75116d7fd538729eb4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he45c99bbb93be0da3f5c7460f855d45e86137bde3fbd7ee1ff7b067dc08c560b87cb88371b762985125598eab02366b5171c9860f6a6a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h44b0a4e4bde82056d13b05575ff3408185c931d423aac543bfb0073efbc86e1be0d64c7d69e53ea0dbcbbf489cc814dea5ac53673ca5ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c3b1d7c884ae920b9aa863eb6109ea9c767e89648a06a0fd2e84e46c292a5ac328d64e4799a03438f2ef17ed75b7272c48e0f3436da07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f5eee997399f8074f7956c56efe1e34e024a731d4dcfc133d1a6be240457f8d95bf9d402313e2bd93c793292e9447784d392f3e0f28fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7e70d833d6760e85a42d202cd8467a0b193e1da3985cd55a931f961306ca609301c1fc5d00636a68bbda9e01b28db808ba90f2f495497b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h189a039639605c4f00a2f543a978689bd5ed55628bd4b05d2eb887dcd1afd57f5ff56d9d5a5bbef51b960e7507b3568ec0a18ccc5fd7fa8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he78298c24cfe834945a594cf2be86de48ce0177a8820bd96f18b420a4e68ca9a1377218f59b9799c044ce43b7bd30f1c09cb6bc576e477;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0738b80520c519aa3168c0f0584aa980199989c02cd7441e17a9fb2428cd1c7dcf2d4d083c8121d020f07bf194392109354235e8ee13c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce8912875c22475cbc8dde43fe56f703d27136eb24b93e196cc4703989ec53f374047fda6c3449eae6bdbe2e33b20e17f66e747cec201a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad018d80b30a045a6ce9e2084d475c12939e85cfb45ba861b9c9f14ad9f3b5ebfac192de3cfb9536e5ddab91c7c14f8740bb23e5ccd988;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a5c66fca1866a858239c347e3bdf6fae1539efabbbac2842b7d70dcd6f5d8502c7523ffe2b81543be3d20077adc5b840b8b24c1f02c57;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf917c1dfea27cbdefad906312727205553a4bbbd277e4568efca040ac9b6fac5760328545cc41a9ea2aa9bb075bb455f7639dfc58994ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f7f0af6418a4c21823ebde7cb20aa2a87ce1f35af91b6f8bccc99e79ecc5d5f41b50a149ca4c153ee296a74c0276abaab9c553473e941;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9a98c582e5edbd50541d2c87c8204bfc81100fd4004a9ed23c4694a5cdca17d49efc0d002d9d261b61033ee18391206dd9be339c973eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19f77179864c8422e257968cd1bdf7208f1edd85701b6366bbb9a0375d0f196dd7825a7e908e103579188e266927af67e0d55c6b56536b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h172dd78cd2eb1abfe0defaaf7f6b07403aec27e462b3617da886f2c1d2fee442a4dc7a7de5072aeb9dfc1360369b97e9eaa3d416109dfb3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15af832c7eac400365db3192efd65cb13354bb9995c5bb800c3a544fc92bb215f723ea3ac85591fa94d9d78d27530abd50aaad4fe90acb0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12bc7d1669a9f0db61c34a57250a5f690a7738a30383632cbf195915d2ca0add64babd3d4d8b8c323b7512231eaebf0cc5031c972fd9e4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1e10f10f7dfdb5c40bb67a5d48bd350366e472f072a8f1958fad6c44bd94dd4d5bf8f4d2034a66e4c722f91fc30e8636bb5209ea102ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7e612199bf7f519fe8c02dc5c0a8fcea9bfb41075e0f4d0c5d6b01ca774f1ad286ec42a2c92298a26c91074876b71193d8137471ba8e0f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13a3cd0a82759e94a9b47632056fc9c0e6297627ae6945b6846dc45032c0ebbbfd4b950784b3abd7881e53220243cb419f1b51c1f581738;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c81cf422d6876754ae4d8056c53d6f2b93e5710ee28ec513073ae6d29deb61c80e31f868f056e243b0e55197cb42397d4d4c7bd9aee839;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13e065948f93133e2692aeede0a4c4f35e45837580caeb3e0abdf893d212ad431d33fdfed89a661272b0d71edd9e3be1723d20f964ab2ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1512a2dbf5bf31474118a4e0009faf1238e480aba9e9f29a82aa481fb67d4339af008befb9ece4dc8aec7d53ee7cdaa4c5fe19a2d686943;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104f0723682abcc7b31f41d7715bd1ffd1e5821f39e816d27ee0e9683aa22bfc756b68ebc0e94aff405fc55cf0ffbfa9ea98d6c5b5ea668;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5b6caa0ea1728184fa495ad7c13a5d705e22da6b7d1bdbaf0ecf985b0b9d65a2777c3053190c83e221d359cd23ec9526e490612407a46;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe272ee9d19b53105c297f34cf8771e05df9e0210c48d4e71716a75063226314bbc453bd56e6462f96128a5fab9a453db96fb39ba37ab0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7640361a14e93d5a660f6ac4df06a97ff8478741adfdf7d97a4088c82ee7a51aeb92cb1c3fa6b541ab9b28946dfeb827bb8f61323b63da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1762b774322890401f01c39063767bc2a423c5eb86bf5c0af214c86a53eeb54e4d092646f6c120ef47a91b75480be3030b2dc2213a6b895;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2fe54adb8840d470f9448564e16e469cc2edf954ba7609111609a937974d06f881a6a42e886d4f9f61b104dd2d86e6b4a2fa3c52b5341;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a61e37af1c71a398ac7dce1fd293f09193b06b790620bb9e56758ffad62d552b1edd7776f92ff9978fc9c6a6f5ee29f1290c54ad329b79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12f876ef483083f9ffcc3ee218ee64876a7a1a3628169daedcda18899bc3a96bdb161f267e833fc53207608e4dfb70a3f4a9941d97dbc4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164e29709aed8b9a557c21b14506c51f36bfe6944ac18028ede83dd4065429537e0ad1388f92d6c6f172817ab7c47e1fa83550bf8040af4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc535498de0abb30b676a0756b2a80eb4fd303ae573e63a745cdccfacdba1db8a16dc80e5833388cfc2af5fdbdbb14081ea48d61d314bba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h97da036c0fbd410436c4bc674efb520086fce657564aae1aaffea85c72bea2884ec513a527d924dc8ee8e5b86846c8b0a8b83ccad66820;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d81a133a052049d6057df14eef3ef4068ec6880dd79544d648fdb73b57422a960e9409ebaa3f9acb56812509a8a09cdda66ec4596ece;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h41b806d16d24ff823729c586eaadc89411d723fb3dc1eddb5a8af2863cd6dbea38977cd559281e77b740bd8c475334bb0408b186eba4d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1beffed39084730dc9535e0041f44dcfb10f28b0476268ab916fa53ea7ef2e34cd00b2770262204645d01918a5484a32141ab1f2a5aa73d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h556d304ca137326484a58c20467dfb3a4d31459c2322ca60ca164f2ac6562196e2ee30bbe27144ca7d41e8dbff04260c8606120c09e48a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h28ce568ee592e3b58ce93bd63b3be67f02c0b390a6feec7c0ce3a7139b9b7db2aae294fc249ab0da05a889d4ad2a2c256359f471d27a08;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h115ee26f4c3c9e9d8eda9e9a325365dd6e4009e4a8d87490bfeb52e6dbab313a963f12ac8b4b9d5bb69301c3faa136965e0ca3ea8119fa5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16a83e26dc030575d27a8b1729ae3ac31544614778dd5b55e91a8639e9dd108d73e64ff670b88ecea97a4c3a153ecfc0cf2d56deb5b666b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ee06af370cb323183e1a12a02f59ff803fa2ef465ed008805a0cc80c3aac44363ff3ec2bda5015020a0fe6a01c5e6cea8fa54a4b4f632;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h878541175e05ebaa9eef42431b3968db5470fe64e37ded388528ad0eb0ac3ba14f0a576cf398b2470c9d544fa27890ecb73cf5f0d5f5d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec9d0d3bfddd6d12ecb3769835603d126aac58c2ab0b9c0cdcdb5b942482d82739aa6580d7134ead5ffdf0ee14473a433c4ad65850ccac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha46f3625ad863827734374f248e9cd0237a0c3436a6bdfa0f24b4af85e0d7cd78df698cd089ed295907c867a346017438112e29972dc23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f7eb0641e74b0c5589b547da827fbcc733daf2d4468033cd49501de2497048e7186f62d953f4c1b6551e3d874bf7917ac18ede2046a49;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d21ee0fc926753f5ca6905132cfe7447a5e86449e9cb1448fe0bffd1d16ba43b18406fa7b2b70c1eed71f45750c3bd1e1ff7f26acfd2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5bca4d379ac0e2a131b04495fe4cf4b31e08193dcd510730908b24e64efd2789d71bcc59a9911529a421d0c21b5de667b0f7e775d9590;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc65940901ad939e789f77c0056b9e7d287270c0dc05be8ca2f3c3ecfe7fea725e4ecc3e3ada81bae7d49d124760be32c741780d923720b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c105ef0f942e8cc8c837f54c6528400b4b1b245f791c974234d34540de4b3d0dbe95f805ab120caf40dc7676d423934fdac70e52f2357;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70605df2fc810319de6def1250c9f7aa717958c2aa078c524d4bbab1fcfa2433a0649eb171024d6f5a686b2ee7ed22f1bb6f7a8d42c75c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15aabde9683ad3c41c142430f5d48dd219b300b89e7c01252b2c1cb4044797cd4f736f4ed26d87f80b1526b97180ef7d5fc3c24591c0aa8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b0703fd1e126183fe0d3cdc306499f0df15078b1e9c7dec417fde25332219e58b7866ee4467dc099ab654a8de4218370b118e4939eb555;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eba2ef3d4304bf8a39d4edeac5aee269133d3642c23633bef314d8b9a2e85d048d17783be4bca4deeb03dab39cb65707de27bd1a1ecb87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24550baf19fd8c631255d8dee9ff5a3d6afefc006e35cfb13320169ba2a8fda18dbde5d26954086c6f8ba6ceca56f0e689731105084ce9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb4a39b598ab362c01d698c6022c17f53f009ea065ec08f6054cd42db36340ef1b9f8925965c29ab5cb89ca3208f91ba6a1c38e7835f450;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7f695bec4a47b06820d385b541cc3faf093bb5034d6a318ccf85817d882fbc05b8eb647529805f2316f62f38dd1aea6272d0f9e355b8e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bee1f5e06fe3a8927259237a99942fb6052696bb6ccbb9ea265a3a7440211ba79a15dc20dedaf0431a45a311a878af02e619ccb178553e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79d80b1293c679afdf1acee79630a93298225b19320aa7792958947f680484fc92e31e2613a4a93412501e3052e332a470eeb311c4ba3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd29619a512dcd3415ac592dffb841317180ba33a9320fb6b1ebb051fa80237af056306fd1a4299f40a7b2a05cff5464e338b29b1505a5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h155e07ab692f0b7c344e496ebd60497640f28672ac4d34a8e284944aaaa4d1a26b95975dd707b2693e817979dba9b20547115b45940a55e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcaf0572d6c3011da78a21d9056c257b592a69dcc963c5bc0ee31996de8d0b020e831c6fb5ccb3b9d767820e106c8da9da27612b59de2d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d1150209917907d31c5c76c586d2ecbeb68f34747c4c5de4be0d8458b30d1e66ebee996f0f69fb7da81f775ea2e79888e07f510da2224;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24e48b251fadee5c4fa932440465edd84e2a4b66a481316f93774753e62d381a58cfa9a6967fd53fc163e736d68589cb5235575817f33b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h97da7c106faa569d8af23e3fe2f096f1ad184860ba81abed2614f0a7dfcce4e5ea72f6cdc14425521bd4871f5121384b9964d5859358b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa5b00c5d49033a5cab7b51ceab42f94e01deb9db192ce3cdff1aea1718c1eca0f4e87c5de360beeb798db5c71492bb9c5dd3f71610107;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b14b57ce75c30a7d303658f5fd8f72d63db0671b863e0f86cf1a3042b75ad5d8b8776aeaa776100b65a2c3706ea23b89077abecf5b4a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h155411768210b2bc665a0402bb3d76c51c817b913cfc60d4ee1e8238920a29345a04f226a2c6b16e56b74c1af86ff903ef6c6ccb1052244;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12a68f1043adf4cb6703b7d977fb8b2ffa680596f73ca68dc13a23708b3feced2985777b50f61d736acb6bdfde2d3a7d179b66b15c3c2c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7acfaab9661ef40a88bbd89921a67b885362ffc9de63e9d3d2141ee4777e3dff8d4899eece88767e1185f0f0ce93f7a646b921b817aeaf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b3c4ee410d2b66ee68883a9ccc23d1b689b92f813bc5e39db0e8870f0bb93a069455ae62b90995340116d70f018f13338fd59dd7c32bc9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14083305d869562a0c9964feae66a01bab49f7d0e22fac8d26a7fe2031a26f1b4b8ebdd860bf91d768b44392f43a67704690adcc9d9e799;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h121e97b9fd6b3379e4cb1a1fc94906bf322a444f1516d37e3ac18c6e26699676478ef2a37ac3b30265ab85c43eb166b67247514c73add93;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a13530be0442128e12b53b4f2c3f29e5334be80aa20fe99b79a4def4fb4196b00a9fe8f49bca3b59e5b79d32b58441ccb151637cabd61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e2a821bce02264f940065797a9a3b0200d18880a7d5576517450fba63e749db117437b91647619654be4aa5ae2d869665ed73b4d0aca61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he12379c2c9924646bd38c34c4cee066ec435c11a46456702f2a06810124b81ce1ebe75605096f5fb60830f51a0223c8c9bce934bca6129;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a385b4d02c133f93bf279ccb6c52563a567ac4ce2f53faa022652accdfe344f5da2ebad3e399ab882a2d71fa1eac76855a87a31781b2e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12dfb61b26a9b6e3c95619a3ac3a21292b248f90b49ddcebde64483f7318ed1a6cd3e35cb3a4cfcf8c170400b2648a9c58c92251528dd7e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f157d3ae69cd1c6e36e630b3ceb497500c2d5adff052f3fc66892cb7fdc4c5dab55139104c31eeec9794e3d348e7fcb602041f13ce63eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ea75f97d353043a45b146757f5a42930f671ca3a6259b016509c661f2078937944adad6bd8fe4bb549059e4baddbeb4aa45e7a7c4bde7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156a09b74176b54d912eb8b896a972820d0593049681e70a46af535f1c5b45c795e967646637467f52a7f1f7afec1c27cf192697bd443f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117b27f9437df65af945d131b99133f2ba0e7733fd592b071b76a2af74331ed77b0acb838b2c7545d1f94af542a816bd51fe7a216b21fee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b96292d705496ae973f4caa2681e87320587ce861651271cd9d2258796f2eda190c52db0fa2733c7aec3a45f7e83658e5bd78c5864b87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12644c3fdfbca5a8ffc18918d5bf8b1f23350232aebc31e4436060cc378f7d9a5e8b8b30295fe1d4d6c22f62dd9ac900a4c8040b26c03a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1461bcb179782c3e1426e16517c8df161a776277e7855137f43478317eeb465eaca52698cd5bb0b923484921fcbde3bb2f5dcf29dd2f04;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ecd98f8c945516c80cee044a1e7a5e6b35dbaa676e1284270794ca18b9a73199ac2932a87b8d8873dc14aaa37c091418a1bb71070fe4ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ad8fa7fbefb3e7c9018a1feae45ee5cee031dd3795581cfbc14ea3725641c805ff7c7ac3cd7d10d9cc0d4d3b11f988e53115e9234b6c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1550672317c02fe83bc97d0b62b3f136449153d1dd3dffac2288ec9c88823445fd619d43003baf1802a0a3d21776dc9a2bab3508da484ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h371435eecd93659d158ca0795cbd6b3b644d9559aa336ef32bc1dff26f0fc4dd4f3e6978081584cf7a82f98fc2cf504ab6f01b4bbbac47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ade057dc3493cf077c3e4ea18a209c6efe937ed336c1890a0e7143321ec869c1a1e7d701da5715d8c68410734498a451202a059b9c558f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d82c8af632a5d775d5f4d0ab6ca56e81fc222a373d76c04a52577a116a605f8ba0c8f699bd3e5b86d0a3981bdb0cf0fc06adaac62c5b4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e69694e5fe9ed786464c2cc19d63b074b8148aac38ce472c9b51744043d0f818d3673b21d608cb4b8e3b8df08a9adc2ed1226f50d29657;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa67207cea6c8b6f239e4f9cb323e370e4c7b3d40b7f73e8aa10d18ae4364fed85ffed9a3dd2f29f13751a714aba4ef88a3052db0ad4fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70986df0d6d62c4d1abe10d13ecb26536477fe67384ab9d4ea0eeac362a4b121502fd780a196ea957ade8ec77a610af8c6c8aca6c94c5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15649471774f6c6ff088376450c3335534e8eadd0e087b0d870f75ec0e520e536c98c2e23d4fc461ca7f7d2413f52e610c8134563bc8fc6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1b0a6ae6800089e84dd483cf354992dd89dd98f9b023e76e009b520f1f35326e83947ebec3381fc4348241f14f04964f148039ebef5f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h150f89c38c8c592f95fada93c097a548b8dd090942964f25fb6bcb7ca6f54233dc4eb428d2d1f65590a5f4c8472437dc8dc46848424f287;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16318c98a2a1a2559396db9904fd0fe7671e21da50df257db56bec2abc2c45ebaedf7c75f20eef4a8c69f5c7353aa1205acda07917ba0da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1187c490264c285aa42d14b8c77197d786176120ef8f1925a11b0b80465b1ed892aa24e877b67d338f6a7c68c51af3417bd2922204a200c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fb41bc12225eaf8a7ea5067d4ec3e358f5b72b8d026981d3d28ac0a3b537b25543259561c34c07c30e06b02a7f4a04039fbadff9a4ae3e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199a81bad8d660a9b72ec4adf52c8aff4e4c372798265fb7a1ec302c5656c427b65f052fdae0c2c9037ceb7d3227a884debd0f2db3e0e97;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b8775447c869eedbb8f0a8473cba436e9b406bf0412d0eb3250b903aa9f8a1bbb823b44d8bd44652a1ef3ae94888acfa2a19aca75ec9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h29a2bd427ce8ae89149cd7bcccbfec432c07a38729f626bcb1032c584341760a0780961ed517ff218d38bddd2a4154a7093df66a1d6df7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151283d41cc331438bb87d044f7115c2aa2ddc38d11c47b07a26fd45085fa44dc7af2cfada5b635bd8e7e84b95cc617f35459bcaac746e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h139e77a352416655b0991605f6bbb83afa338b3aae47b40470397a2d7a00b6afae82561117947aed847ca11597cee08e782c46e91410a7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4494d2b03e28298c1b38071539856d743fbc55a7884139b5b2faf9d3da0ebbfe324d39f2485a17eb49b93d64290dab94929c2c22c9be82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h150217923af45e5acdf72174b8f02c417d9cd9786360dd7831fe083a8dd5cba7f4a48540eca4e70b6fb0b16185e46843ca0c502c6ac979;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h187f7eb6288f32ea0242bbca30b2560b539e8029ff6d437ef58a01eac530612e0d9fd79173f8fe25cf372034a1a31ed28f90f77fdd688db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4d96535acac395ac71da63c0078454794af98fd1198bbee1cc788ba23a7714a6472d9100e9e8644c7d4f435a8b0440c41eb9ecce737a67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2e905556c3e2020ea63cddbde3dd52a0394f0551fab666b846914ec18707f70beeb694ee1ca074237077998d2eea6a5f934469c69c681;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h457ea8f30a38903307b06275d4f82b2e73814d92e7fa4d463c31c9433038bc6d613330438291ea74e2290239f1a8295ad389fcbc260f1b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e4450ef884a433073554e367e56b925561d2c49b21f2b0510af6b5d4670c63208a0bd9c96564182c473befe8a5a620f30562bbb1c8bb0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e746a44a9a05de904bedc09625f08b8dc062b608cb452a10b59bccae379791484479de11f75885609ab25a9d55a778220e48bef81144e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b2c4c0a73c0d9a6ceaf07de7dfc101a41f2d8c90e5ee2db13dac08fbe2baf6b37648feadd31a4482110d007af695c9ef6dcd65d430b02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b1509747ce3c2e91f14a0fa2595dd4a9ef6c54832a77087539361a59385d68a8c20ed18b132754f5bbe81f413aaf569db7d19b61f58db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eeb9cb5cea21a08507b3669b5ffe51b73dc9e35749d1ffb670bc3314471b21d7fb81b4b90d2174bdeb084e0d6cce4e92d0284d22401bd8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h27cb29a60e6b7643f182be2c6bbe3e5de1e1031d7a16fe4e131d96b035fce2a85f3f717b6daca02f773df2dc0acad1416912d09b75bb42;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14764a2e65fb1e876b3b1ba537f2e8cf78ff5ddfdea064df8d19b95bc80113534fa5d3949caa57c122c5d0a9540634150415c7ee7c1f74a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8f8b56ad117e7dfd77c7605ab9ce4e1fdcc28fa9c89943356c26c7a2e2e357b2c7a2c2ca3169c492f93b98d915a51ae4e78b3a78cea930;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16bb01fee398036b3baac0282c9b97d7f35051af5a1d89fc19d989f2a8fe4210a28580b556dd61d7e8a14fe6be6d3bc0804b19275e67f9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1683ce32b84ad83a1b3129caf7fc337a194f3fa282ea9b4c8ad20d295f94a11dd8b6e5bc218e3bfcdf82bcd969d67d08dc47c9f61e0d634;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f9872541aed6dae34dfc1cf2061e595ffa13185b1a68f0e7bc67452af27db3e447ca92732e4e7a6bd0720112b10f23cda3bd65a48053c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58a8ee2fb995f2c7000979a583840b4747f25cfb0482f98008c3edad74f932734041232c9168ca7ceed992f8afb7948847a2c30165af82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h120ecb2852cd7bb985f74b661ad2e85de6e01fc65ab39eca261a0fad536f638cf65867faafeb6c07cce5d03e612f68f905f2d118454f2ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hedb6b8367ec4f0bf68b7ec7ec6fdf1898c0f8e18b4c352a6b7ef49884d11d59dbf6ea91d2a8e5129427724374fdbc883d57944f5003fc0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3b885a0b473304d576a99a21ee0e6f8ddfd88188b31991fefb9c60f3b877a857c7ec34f18d30ffdb1429775712d13bf33de44a9dde6721;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a47440930a4877c0e171dfe45231287bd0eadb91e4df4117108b9258748f37eb4fc3e9f649dbe06af0a31c475613856e9560d7b622f1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179c0a9b109896c537d52b40bcd9b618145f071f591db41f5ef23c30b0aeb734c14346a76e2b15c433902e7006245c6caa18a7c90876c4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb870bbd3670b62187b82033d04733df214e0f9a587f8a2d94c5c3888aa9765499250a60f659972337755762072805d93a2867435b7cd35;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3944664a8400f358c2efb8705d7817614e3ea2dffaec3413fe453fdb0b73cb72d1511f800607800f1e62f0525eb2e288ff0604d1b062b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9470a11cbe2a0ff478f9c1d7c6540a7757674ac72595966ea2682f13cdc8679f83f77f02bcbeeadf676bef4821fa77aafec6cb0462d4bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78620a92eaa36d3b435d3fcbf995c94272e7f255dca6fe875587a2b80f88a888fd3d14db45eff1ea3314ba22bde356b01a5d2200ce13cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17587952e02507d78b5c31c1ba635fd93d6546aea2c7efc65d071ea0196f797189ec18b06605c6282f75ac848c24137eaec5028d5a2b122;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b4890a349af71e3eabd8b7f77a61722760b59a7aadf66d41f540ead610f24b48245e5e59928f3858df9411cba1cd2e35dd9f221e1b67cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c36e792ae74e3e1aee9ad066ea824826773bc9a51fbf2deb2b98e76b8d1a5cab54d5a52d5aa771faee7651e21e095b88655e8b5264d31;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17e7342b63570a3a428937234d504b2b871fcbc9d3019d4c06aeda91013a217a31f981bb7290a2973b8b85532a3f8d73a043609782c9bb5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb7fc025d07cbfaeb612e25ad7d6c10ea85554be07e0739084dcea04880e3fa6dc4299ddabc8da6b75894db39cfa1c8f12c7d6611ebbc57;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h87089baf17cda6db156f0a95c350ca62cc8f78d05425c36109144a2439236c112235e7cbf244dc0854af80c698e61ee8d7d3f1a0e977f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf0eda51fac8a6d6a7b9d1706e6c7ebcfb8f9971cfbc829a82a6983c6e859f981185190b0fd886ddc403d2b2d6fbb79384dfe7a4fb00d3c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a8c95c0881172bc8e4b4e5826bb1b774861a75bc69819b3630aa298ac6d675e6d0c48d451635b8fd92af7da7a5c9c87729b62917fa4e3d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181b1f760bbc8dded6cf989e6f583c9955416808a89377270f40cf0cc85c5dae48decbce12219e3357b566c7b8d7bedc9276c6356548d51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h250e2f26c1846b6e8371cc4ca2133cdfe862f51a180772ff9cfa32ed3bd34d3b68354bb8f83c448e22d6ba039c1a090591a06e6667b28e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd972bc7c4100f00b03ad2f5b6206ee40b5b9509a66167390eaf95bf47b7a716883f60c7be9c44b09847b24b0f0945d7ca2ecb7cb9f0893;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17964ffdf239ced75c0261088d2695ddd41468f7c84fb050533154e0ffa383b0af4145caf4f5383ac08905f244966103c12ef5690cb66c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14df3d982f0800254db8b674361dde049dd993b2f3fe0e66137afc2d69a3651abf621b123d7fb3761d156a3f07d46002936c3d1e997b6df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ceb82dac5336c7ebc018e8dc3d45e1b98f83efe233fe8979402674c96894e08120cb06740f370899e54b4bcbf311ec53af86c006b7642d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e18a88ec2f1f932243bff06265ecc0a3da05d12fc6ff5d8b12bd828d9bb926edf4f382abee066a90dad5800c5a6d2dd5346ea34a342e47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfe560d04859540756594d1be53543727a631e609bac75bb2250bcf23a3b92823cdfffafe78b3737d772a966feb8234df48ed2d1ff2c146;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125d4144802162f2ca73f5cecea58e7144fb7943fc06d0bf0bd56beb13a88f28de447916b5c561788dfaa5e7721673ef13c7bba54e22d9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf050248aa966585f0b494afd86419b400c9e937f4b98c4339e200c8168bb9b6a75760a8d32f27faa2d04d38d398bcb1af853c3b28cd488;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e981d0466b849a6af6612e37ec0829a455993cd6249860b4d856ee539fe0fab0ef30c358f8661bfceeeb441e75cf6ee58dc90d943bda0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2ec1859a002032881cbc856516cec18b9db6b782207de8e4b768e801ba27dae135c6ae6ce529b5f4b81ead55b22c011556a23a3326c357;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h177f1bcafafc924678ba984e6b2e423da471ab1d5e8d2e36c40983fbb7c1b25bb6aba37579ecdf2d1a01991145057751b0d5788dc33dae5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a82bea2bafb0ed061c7033effbdcced585477386943ca3e59d7a0faa52b382b9e31fa53befa525b8e1c184181b47f25e494dfe204f9ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e62cae5bec5ca682ccb756b2421b6fcd2c5ac90bd441042da274d89807560a62baf05d5270200d281fccd0b34821951b1920080220cb88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f0295a59f33d98f74b3400713426d1e13007efe21633e65c2ace4bdee2de3d68ca260b113c5c68bbacb4dbaedda7b88ace45e436be57e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1978aedc3da1728ebdfdf13dd8ad15799055c6944875ea8a0be1d111f5c1dea408d71bfc38f36a6d4a032973b47ccea3f905e663a7dffd5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a1717251c59d59caa0332e79427cf19d48d2d79d1391a5342af9dd00b064327a2e93bb31767705e79462c77f49104d47441749276f867;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18deecee5156b160deafc59df9c7864732d16ebcb9d72645c52e92d7c176950b92ea38861be94c561324f7d8a574e3c08e0e4b4a2c94cfb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f140f48b4ceb758fecfa963c19fde8144c92dfab20d7e2f30fa14708625e6a721fb87c79d99f9a525ba01f9a542b840e2599c5b7cc727;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h413c88717cc3d86cb57a6219b3390d79b75739940a193e2434271f6cf218d71ef398ed5af201b68e7309d0fabdd803af6412f6342208ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hebc75da4f9fb8a7c34c5ec1e95c7f593ec00d8905fbe6cf8fa57876d0cfbd0eafc3e209f5f22ffe7ae385adfadffb20bf63b64531a1903;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h330ab1e71c3c9e9895f336a9e9953054cde8bbf544fb955ebba32fc4829c9490836f9099d17078244339d640ae994e5779f5f6ecbe8d02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h627e617f43fd3765e91a2a10f7cda701db48844ef88f8e11dd511c4443c2f3d4f5794ea11313ad1010a3314c34e82288badb219839d51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f6507b8916f762cff624611bddd2d098c3cf0a8f5b30961829a86419405e553236017ff12ccb44f6adedce12052c863f58a4c214156a7a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b8f21af4ef903867ec605aea7a6fdcabe34194c0263d6844c0fa44134f79927f852be075c7aa56e4f373397e2f5ffa84eb056efb1c2b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h173208daffde69b60602505139a29f8443a630dae0caff3e03fad2d002eadfb3864f232b57ecb8dcd08d87d9830bd37a8b2d20d0e79102c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h24367b5923092ed129cb14406e8cbd08d27f25bd95730a48abecf583a21f844ad4092584e1033f6871a500b18cca2036ad0d73278723;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h38f040db5d6851a9bee38d37cd416135f936ad8a3aae8344ab775d9b18f1df4a7dc2e44302b3fcf2bdd05bef01b9f9eae1e10cd5831f92;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a12cb4921a146d49533c60149c3e6e9a86ebde990aed64289a33c9bd87b7b8c5720dd9fb17c7af66ca49fbf4999dc4d393ff75bd5de3d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18948346861355ec31c0f397e0ade201047276eea2a6721f38273be7fb2b5500f91a8b850e87b5a260cca2a86e6ada13a168254fc489537;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0df7f290b6c0e0273996ef87795f0e533fcd6e77802d107e418282c4accb9e4b76ab39eb9b9e0c6e1d4b7976ca5f3ee7a71bd17a19824;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb3a3ebfce39772d4fcd5c1a81483b81d879cae6e25b0137950d5a263d4915fc7fce61315d0d3e6f165d890d9c37fd631ddbd37a19156c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1845a24b37a2ddf31410796cd0edbe18f6e05c8d99466e25af8a136f3a98b6f4163a1d2f288339bb5637db6310357729cd6ea6648c114a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10cae847e578966193c45f45270816b84979d28ae781df55e3d521ad78ce7770b4ad44b1409dc25ed4ae5ca7815c90489acac8b960708bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d254446e583bc6c9302ef0a10901a934216999667eae8d569a6bf070cf0ec85e1a6a52f15849b6a7fdc256d5a1363d69d394b97c6dc2c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf890fcef77fa55a0e67d594eb8d0e96726b472d81d9dd2375abfd110f7fae76e7c2f73f96ce84d3ce87b889eccff67f5f38905a6203182;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha312c4dd2aa7e662a9de28321f7518d0bd98c80ed5729bcf892edae0b3d4b516ea13cf1119800e029b97acd87c161a2298ae56daf357;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79829773ace738c88ff67f0ad4b3f2e107b1a69bf2d5e3ca2c0a5f0f0149a64040ba69dc78d2df30c1f449bc270734dbb0cbedd33c8f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151ae17d4d9cab161496b326ca673c7b7cdd0dc792008bac143cb755b6dee18bd61f763a4da2a16e737f4db6341b7890d454679699baa3d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f22d8b8ec8b3b574a0133d5e3e5d37d92a4a840c8b642a6fc3d2209a5b9d361056ec9ae4ac882d7dd405966a1f0885487863310b9d3b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba765737572f5a3dad31b7208385a012c8f197c01d25f262a36e0ab642fea50d0a464dba82a378d7fa3b44ff5af2ff0991d124e5a5bb87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15afbc3aa9683561811e51dfd8841fcebd8b0f3f40f70838ed006efe6af5d2799d309bd31bb36dceb66cf6b4684db4c5c68e8ae1af35b29;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba6a6d11dd439b0a48067dd4689e691edf86b1da66d4cc16da859c841c84d7da76b42fdf07ec9e84d6f57fbbe7167e3b231cbf5d4316b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1722720920cf5fad1b1d688b9469ec90a775ec3adc91e98b54f0adcf336e91bd79b2ac0ec2c0f06cfa64cddf256c8a649c576416418328;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h167b3273748fe01ae1cb2c14a012faa55772c4e66b9bbbab35495e6119a1cadab019e9bc65d3821c616d95eada68edc804f13425d4e7c98;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h44fad7864f48acf2488f466a20fd7a76bc7035f357d99a20e269249d20b9c304f04ac9fe5b7343cf465c42e86ace4469c64a586ed487cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b6f9516b76d9c7fc3b0a97e4e00f195b3fe70abe0abb705f989ecb1e9c64ce3bd09ced15dc6d0cda3e71db910801d8dd6aaf2a853be457;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f8194535c7dbd89bedac3dfbcd4aa28185f06dd4ba88863a8b045e37ae601a03d512c22a682a13f990ef7c2f724e0d76a3205c22da32b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha35797b0ee5aa0115e4a3347a95aec37f2569d0844faf2f38c2b38e70e04d09b47434728f5c01fc4d489042a3da34c3255abc49c8950cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h62dc1d494c0dc385894c1cf6d8194ed3e864720394bb6878722e89fa8f6c78c410cfb52c369c8700119dff725efa023fa150d0c449ff88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h56f05bb0885394932654d8d991d922583833bf579e81d1c0470bef1f0347ff4d710fab1b2697b3907cba5945b69132845e780bc30796bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17e8bbafd6670d180f3069aea303f42d43097a280c2af424a8364952b01a24e60e0fcc9d224d44dcddc33892ed057ca49ff0bab1db78193;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3ea10f7603d3f1025f463d0b6b51637a7913a9927d80b3f2e2cd888ab2df6981a32ee6e4c8656a979d41a1d1a5302a89f1067200aade5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h33e6beffa8e3ddd8d2c8bc68b22d54603effc451ab286ecc08e0343246b49a692b9466e540b0c303c9b89892c2184b4265ece6f3d8172d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a9db4ad4f6f351d2f8845578b683a702df3cf960c252ac84668d205e4a07bbe8c56d2230ac0178d2c069d58ba161eaf5ab62f279238f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h153951052d6faa57555db4547360f4c28be37e1ec61008cab47f898cf9a1dcbe79cd53c69a0f9a7cd1efa9fb034c35912a3e7b9b9f76781;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1921293bf46c51cfef30162a2c686218f3a2f9c58dc97f6f025a554a7f85c275d7b910b74ed63296a0c88c82eaf8fdf91fb42861a4812e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a44e721b7da12492d14994fa5f1648308ba9feda81b533ef15e7335cfe0a617d6256da34c76f1642a195df640f8075c8b1e3111d6233c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6666abada0efb0ea5224f7b8deeaf11e2f8366f0e8eb1422c1d7aee184f5c99ac94ddf10963f85b4a8a76454e09ba1452902dec9b9f2e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc36b41550378b4164518638e7a53f4f4fb6c905dea73371bce124f0710b71fe760da22b89c115e75805a82ec424985bf9d981eac077f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12463e578dd95cb33ebb17c27eddd78b25bff325ffbe6102d292ce70fe5584d3ff1e921e733036d2fb51c2dc3c3840b9b6dcd7aabf51901;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12fb4614d12c185a595af944e8f77d7ce497ea6a537365833efc610f3f53fbaa8637fdf984e4fe815d61d7d79c07568e8627d439eecf182;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11db7ee943743c3180db098979236569d2b45d19ff67bbf3e7a6cf523189741a7b3b58d01bc90841bc5ca0504fbd9fb28b6c916453db844;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c9a621498ac12d60b0888a6fbd1d8b77006f88a7fbd42779d87c28ad6957d8827afcae35216c7a00b9e2719b35a7fef8e25a9f77f978a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd7d6e6bf22e128638a8fee8bbcff93586df7253f99fcc1b06cc5846ad7901c09550283a1ad8fd1323ef8324e0881c005c4c3e3287a3773;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0ed85ad771cdd8e5a56733e6d854700d989bbb7a2f7432211020365ba27b3cbf28f58237c6e600e360e1385fc4aed2cade4667049feb9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a62cdcdaa7c82e57b9270440ca4cd38b3452afa6365aa6ae460a822ab55caf024d31ef8d2da7154f22b76fa0e1fa108fdf401f8f0cd1d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117ae37708b08cb29473524053357aad2e6042f32dc289e9b3360ebb60328b98bc4027f500c76620107a19249fc30cfee0ba9ca3a5e0388;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1015af5fd41cc1aae88afe3126959fa89d1f582605b112dbac7fcc61193031a83366e628c6fddfc04d9cbca24f3a60135ff2872f3cb55d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h353e0ea3a89ec01089c1b5bbd21edceda7e9f04bc149f58c9164199d31d36b2e8fa6e97cf6fc2fd0c07c6b60ef563bfc05fab48c93409;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d674c73c02922f9fd5984612b4b570681a8794f9b76d5fcbd3ec954211206f83c517d2a5ebd0937834880a135410f4ce4212f359a0f03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbbae59a2e890810a0942fcf79d19712d1038ef15a9e398f2fbbe784fac642fe4c725a87c08080e97acddf9eca4e12a04445ba47cdb6029;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66c5c0227352a6769e5c31f83f5b6d185113cf71f77020940df8693173c267915541f7a8fd1d0d648c0e0860aeaff7124b9d96b2c1980d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e81e921cdcb8294e5ee1b9da3143dd2d5064516bd2762d740ad14ac37716584dde50714466ffcc671dc906cd09506d32b22dcd7e3421c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h65930b5c9001f6a549ad2527048bd26c4fc1f80da2d66dd55dcf5f41824de972afda31b57d07b6fbb5a7301719da2a264d7fd05745426b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb02aeba767b4df8f972ba41b5e048e86c68c22c53011080ca2361dd29e7d272bc942d686502fb81865ed5a8ed6b4097059b94da4a73a81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c9f97dc6ddd985eef66bcc3cd8ab1c0046a095d887132f4a1df87cc97e9aedbeb0670a8a78ca5a527b0de628d993c5819b4bf7441748e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f020bb980feca77843ac46c1bba6e799143293aa285ee71f2968f06974a96efefab489dad0458da375e23125f9f2dd7df98caf538a9264;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d9e7d605a81333617ff7c93bce9d3c1e1c7e29f3a2cb9bab43351b6ab6c55685c6cfd0368ef01e840c90b415c56ac5a4517994bdaf733e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b872a47ac5b5b6b5299b21c1dbfede5e193c86e3626d07b0eb765bcb2feddf55103624c3b5142f82d166ba9b70b27ebe3fccf20ab3b01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2bc58bd528c116f8b08760704d2d90f3ab5c2178a7984ec82d9870de1a2eee3eba082e1e03467ad5630f271993993c20162bd7888ca6ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd3d9cc6c679fecbed8cfecfa302173c85335c772af8be5cb18032173615cd402c968d8717838d3946476d374de0f631d63684a1f5ec888;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ccd1afd743e3b00a599df97260116b7569b2574f5bc0b2c94e97e239ed38b012fcaa6a651590411ba46b314ec1d9083c0531a43357174;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e5b3a6d35ee1ca48855946930a72181240d8c6563ffaaaa1f2b33c383224cc07361d781594af9706b144c3d52a5d25d215b7413c3c8dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1043b251ca55cca9bae561a63d023f28d7897fc75e18d488bbc988639e42bf5294555dc532c53876c7a080f9e102e3d6c4f565e01206cce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19c5ab8de65096b74bdf2bb3f360bd8a5d6deb4c3ac9635b49435bc64bfe54bf3baa959c18ba2b98e962d333b9e9e84f2f1644e92c072fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6178e899b2fdb3dd1473692b7d169a4620a7f25f85b8045fe840e67eea57a451e15fbd909ce0611eeece0fbc21e83a50c3e79b06298eec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef32da53875c88703b37445c048ce34174f2fefb63095da0e963819157770accda7748e6621da486704bf9a8c23b7a4d435de854bcd330;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h121bc31297ea688c6cfc36b2dc8afcc28872065db70fa72637417da2a2998cfa8970a9f91e32be80e6abfad6dc46bcaad5e1865aea7cf69;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15b78ded9610dbfe9ce3de673043841310d9fa6605a6cc95f6df480956cb4581e08ee51e507fd4f31e528837789e602d8dd71faca803715;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1059ee9a844732c2f340dfd4edd1212984de806a094605b00d0ea7f6c10c85a9ad54500361fefae0e701801c26faf1d5ef716a2b3319f7f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd7d3d8b2c284b38e65f800ec150cceb382e35a4c66c566a909e236b356f0cb2429a495eda097c0ed8cba875129ed28234f4fd2be1083e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81d73f0163cb936701f367432b4ca8defeefa2f41b65e4015b17265d329bab2c2c075a440edbc472bd02b256a723f56c9867f5dc53cddb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he51e107e3745802cf1e7fc97fe1ed54590f47bb0cfbbcec8559c2e1df0229489fcfaa0d7fbefd52162d20e3b7e57261f20799828ae0430;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10baa29d282d52c434208350576b6135d301f793a417a3e074d8ae2e11c3d5ec0f06371967575499223533df27f13d6e8178c922c57dcdb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h101ffae2077fbad01d60197221343e42a8a346b4f1db5de50f5219db6e466756ecf434c368bc12d4a9ffa932e1ba03a6f1ab40db4aab767;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf385bd21fa3689f1794697cda2801bf09a8bfbd3507b6afd73cfcf1e10a9e47ebc9ed2b4f0cd8e6107898901ceb6ea63cf0b1f1ffbbcd2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1414b15ca98b2905c17e39559df8d729108d2631a4aa7b317ae548b0314d628cec80b0dd1c4e4001d0ed0edbb7b1ee67ff8253bbf958ae3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h123b5eca8e30f37327701a3f1752212709425d3824b6422818d5d2ef8f76c153e7f3374bba3cecb3396f3d160ee7147ad7b8a8f49715470;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha8793f07e6fe1581859d6502a23ae1e1c662d26c79a2a0129c573dd467cd5ba6fd6066e8159850add6c6dbcf151eaa39e1138cec54ffe6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18cec5d247f7e9bcd43148b4edee4f5e9e3dfb5bce0393c96e1db8fd32c120c882193d42dcf32212717cab0ca87caf363113a2011fe1523;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f04ef0fe9e548158fbbb452dd1005293716ec69df5bc2da16c56c965edf5ccfde7390ccfb5d468786fb67b41a24d2dcc6fce3ef45eade;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1074aa19ff6d51516401a8c3097d80031ba0dbe3923f0a60ca84c1cfc51d98d2fa585047dedc99fc10253a83f8bd322ae283596e5ee06a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdbc29c9d1130f284191b57519d15e9fff870a7de4f2e19bf251fda60bc37896b3abb014f9d0dc8cd4a2e697bfcb7a4cd24c5c2bf43e31b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hef440fe431380bbc61e4f4051765986453a44a68e394438b820656a1d5918000ea7078fb52e176e4d528eb496a8326d0dbda3e13133784;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b13bef6e98deffc524cfdec30b1ad8551547a2a6d1d5768b12bff3e9be9c53cc6dd478d589fc32cd3889a2255fb99c54da5fd625d3ff3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a46cda3df2e6bd8fa581db42904db04e986c9d67167e4d19962787c4646807e7d5273192111fed3ad662a2ab5512102d8c6b5b5fb2c842;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c287ff94c1274295bd3a26326005b53dac218e79e278006a12b49ab7e0f475f9b7b86be52f19f5cb4d31b54bffc549e4818c8dbe428224;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h318b23fc810707a174ac608560e76132de1d9f7fd4f32665b9a36c3836d1c41cda334f95006f8b6ad5b2ab84f3529647f6fbf797f534c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h156b8990fe84063edaad27d8e58a3656b7b7a5b0e2998e95dbf3a417cc56d4d26e97794f277ebb8026224beb92de2b976f9727b2c6f96ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h108ed348c28cfb3d87b2690badfc6084fc9f0f85bd8f2c04b63f538377f1c1a5c36d6338f1c207d24c50d3a167455a0af6d9d83cfcc8f58;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5379614428efe5b686b6254153e0ae2740f7e1375729f61bc15a9e84e46139e0907cc2146ecaa2881f35a38417f0daccd759872c77333f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbdc708a8c04dd1ae98c12678b3a0ac712975083212eb42d421e06e0f09900d55fb33ba317a112fab864e8c3370367867fdbe93944a5645;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2ccc609750b105cf7eb5e766c6d535067e6ff7fedc0f568947ae379aee7aa54fcee2c4af54d954be7133d0c5fc2cfa10562b492e9297d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18652d0c87b184b4514de97bbc97b170b23ce161f980b1c20bfd6b6ac8f3c676621e6c328cf0bfbd221ade69b5366664963c8b9961738ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2be7920e1101aaa0079ca0d0667dcf3e77365fbc73de43a925166d57b9fc771c2033de2871daf2fa4bb7a698c49a1826f89ed798f3240;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ff3969932596e77f4ee9416e7fe59e24c7cbd261f838c347f0fb0460c324cdcdfd9ec07073340e9ddff9b4e9ceeb2c2048fe328a90497;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1adc166b34e01dc4e673231af3f6fe312384c29f8567d65b52b9044fd0c849cea178d4774af13f4f4c4255ddefeba186fcec497339df5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79cbcd23094f4d80108370be7e44c0c007cfa33d748e52939d9a0ceb4e761003962e72114482654ababad57744aba695370c40a34b671f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c2babb5488ea516aa86eec4700c7755ddadc605a2a7e37b7da751187afaadc6864204f30ed7b433d669b34a8f4bd93ed12132856b5010;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3adf7f55ec5ee42688be229221ec73f28ff6a21cb824dfc9dd02aa982e1001242b513e19a4e954a2843cacd7643513b5e709f55fd22f8f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d2c84831f4880b373a9de4c761c3dbdda7247c8f5f0d723877833060c0ad2ea24e0390cdf8247f96b9519d0e50e9c5f15af2ec3fa391e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e06c220d8cbf2664e9e753724f1dd78e70d6132026d03b320efab103683b643ddcabf16cf78a67193c052d6d86a745541bdd26eca5e20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f8cd2052d6b4d6eef29c6e05550663428036f22baf7c06b08ecb27732f8f64a5e5cf071592e2336a23452761d50b17752adadf9ca43bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c169d7f67f5f1fe8cbb263d8ac1e87ea1f2606194a0c13c75348fa3ea3fa680bd8d89755f47d671fc87efb0dd2a815d9fe61d206a959bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af709d3231083765111129c0fc3779f2f0b79920391caad3554f792673d3d0a5f186e3d82bbb41d96af7be1109831de84e3336c59339d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbfa0494c8ccb58429cda01f31bd8ff89d258a3d59c793ea6d11acb8ab54d60db02bc7595cbb099d6bcfa8ba8a67053d19fc529a73b29f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d2910553cfc57fcd23ffaedea625a2795a49f17eab13088aa8d139bd21594ff4e7ffd3389b55782901d38e2eba7f25d6d215ad0cd2a19b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf91ae7d30f5418fe25f0b54dba25a4038edd8d2cf621633a8408205260b2f3138a020738ca3919be2d572969283fc762048de0dff20f3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb589077d0559efad05017a6bcc65b44d155e755888d7c1421f702fa94ec46f547afb4e59676a113c798cec3c9f801af9f11409440cd01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9246678f80091fd174612a4eeb51715bc2dded172a446ffde463fecd273feb54b41c9fd5c065f90884a196acb4ab3ed1dcc386ec327d70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7416d6a91639b6da870f2bc22fa8eeb5f8a5606fb48edeffa6610f467b8fb5109c77e092e953b8c66580a3bbb0aec9c4792f58a30d67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1479194e591c383060a98c070861e97e8685faf8d045135193644fa94a4a70f6762eebe1c2b18e1796b3eb08195739ba308bce7e1edfb5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69e0fd472c4bbfd3238a4aff92621761099e1324cea7e922a3f9e958af0a5dacf53d8e6d065907133eb758f11556cff3222023aa5c221f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0384b52fcb8856f1494f114a1150e6884ceee27b6603aef4177ae5d672e624f5a3639db2b610223322a71b99386f7dbb7c32c6d045afd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8802eba37bf1a4cc76d62e00967d9e1fb98cf0c64540a1113b8a55f0867d7840e9592308bff48bdf6eb5c12000ef6618793ba0e2d5afcd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a97508b137a9d8e5e87bb9f5c0e4ac200d4d26bcea95eb2c8b5633b81871239ac8f2390101ddc243250b525e52d98f8f4472ec51a9ff2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h378768e56aba4bf6983eeb77828717164bb18a924f43b0ca888bc035a28f6195210f2d42302a7ba51e19d4a0e86b77bc2e94585eda5cb4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e325a26f5cc89365a67fda94ad74add62539db98cc4c9b5c69745b3372960171bf10c25e3b8fc6954d5c24e1fa079d91b5f6b1ecb7bed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha136e12efbd0b87f8d509966807ae7bd7c2804f833710e548f7a0a8cb48591f0958e92fcc4e6d157218901008fae10adcc50a53da3c21c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea062ce6400d583db60f5958c1aefa8ba61d9902a8c1d987523dae2f6f7f2c4287f3fe1bcaf6d5bd0c0eaacc4b703c91a6a66c090ae700;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h195b5a5229a1d81426c6a94db9bc23b76aabaf84bee861701d122f3824267409a471fb1d303d2f3d216e0e509dde8432740c783da53a216;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11926c48e9719a9db6250effb024ccd13c784e6dbe1a7c3a7edaf9fbd83db286212d0180a7419d556d579fd3595f1c57b5409198f7fc53a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h132ef6ef560e8775843fd985bcfe8854f44924e63e2840fd8c73d4d50448bee69190ab2fcef65f73564e4e3018e9aa1312261ab84e7ad0c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14bb60a0c81d6d27a118d418f7bca99094406ed8d2a94e2b1737742e0df22182044df18fc5d4fadea3943d61ec5ca4918bd0ee8bcbcb1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h445cd5a7c8571bd915cf8c6c44eab46554518802d3f506ed8b4d3b2bb6345f94c223a9140cc8e39872a06ac09f870d968a78bd25d24795;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f6d99b4e17bda0bec4c11f8a31bddd99a284fb0b6aadeb86099a13350ffa4e8d400ca6d0a89467e8fcbbb0c2d002ce785e236fef4633;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac9f670e11acfb11354a9d9c61fd5180f91bc13b0e9e75a9bdf44d083d5ea89d52db579fba2a9cb14971d53260c28afdb204677ef268d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19738968d2da429999759ea4df6f5d983707ed990442179ac977b8fea448c2566fbd20263b7fb648427dd79d7953f8dc0f300a3e22c71cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd4c2d604a09f0bdf36982e111640b9cbeab93da73ea1e4a35343b481da345e8d4e85b86ea869efc6fe70f7377f5cd075b3af9b4f79750;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb9f8c13f2ac19b0699df3918a8c15015a2a7b8c77cb4bc0a234a8dc68fc820991a15a8598b091f6c6e506ec5f972861eb39162c45ace1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h50e5264cae0ad254308a1a71cf2581fa7ecd91a1fb8ad93b781a27835dc0822131acde11adbaa11e63a6d0f452a51ac09850a1442449e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18e731063a9e4432d183a35f0fc235eaaa8a7634844638b220f1624037916e8d63a3ab4aa43558e965ea39407adbb6af6fc942676c9f50b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7095617b783e5ac594399a108c6e61800faf31f3afc883bf80dc3e66840c8ae6059fbaab268985375080fe66daaed5d2211a0639a387dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb5c670757061c3cb06e3860b7d43551e7adade6e435e9180df76322ae8375e19f227b8898718a7e9f5035924ceeda448ec0540f19cea2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7857d10e92d94b8b3572490560b6e2aed57e7b12e78895d938c75bc640f436579dd486d442e2f870d78293c228b0d5096e6d469372f80f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2c2bbb4615043f9446adfa82bbd4d4727bdc56b2b9a9260fd842c02f0cbb34d3bb4dc0ea2755df0b109c72ec4d5992f2a140dd9097d79a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h88332c3fa3cf93aeee207e20a3449cd3d48781a8b84b320f8778ff94be68e65683fabb72b8d3f0cc84dd17badd3306fdfa1d0090a4a389;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1deb93f5943035eb1e878b00dcf9c90982e93c2c84008f0c1293f49dfa0ea3d341489fc451c2e6ff1f9594cbc885fc655b2170add47d791;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd4507577ac2762f441bdaa8e9292f1b32db82aa33206f23c82e48de3afa0ef911438472e3434b8f96f3eff3cd451eae88e10c85a68dda6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h52ac56015195c7ba7a90316e63b5e786cf5c02cdaedd0f44b33e468aa393e3ed553b376589f7ba22a501cd5993887a320361ba0603a8c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e4faf743d204acbd4ba04abb631ddee5dd719a71e2e3f601d685e2805935229c556ff0a9ff5b100432cb1f43df75e00b3d1110125246ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b76af72452fb2e5680291861ffc54506769a04c510a4b99a01d6a5e4e8bcfeafab4fda79c6e70d8ed47232b11924722397b20c873ff67c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5986d15e934a2309774fd01a2cd2d2c3cae7f9c09338d10232da639092e70f698a1464a7ea04217aff1780bc12097fa5274d6f9aa62217;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c24801442565e73418e1b1c219d34ff6754029f02618ca5b1cdf11d88df9198a35824db293ae4d1f273a6006aa3ba67f6e02b1cd00daef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dcdfd8b65a403d51224fe8bb32b4ccc6646c6fb79b8590712abd41acb40d0be99084b376a3fcc153afb1270a34d4c374e7ced6ca43d80b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af2bcaf107dff1d3a9bc5a2151d2e8684e26ecc94806fdeb9a68c11831efb73f7752e3539f69a481730a079568a480a0d786a29a54341b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h630114405612c4c43a51ea98fbaacc477090e8dcf32e16cc062c90fd70fd02c47cb1e3b0991e32d7d95cb27fdd0b3fe8bf18d8481fe887;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd9ed784d728c886100cc2d64a99d1c551ce765e3afbadd1a7e2f2911695514283673d46feba53f4ccd31db4438c789b53ca368792e32d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8af0ff5bd8f75d0eaf3253f2a094e5cfcad25e31deb04805a52c782df57758b0e80a62dd56774e1a2b308f6a5956ca0e104e49e43d9c6c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h132102805533cab5b63a118a799498842ef2feda5c24ff50e207f2a8919508a655e28fe008d1b81e2f2e33d9233d1f300e1957dfa6e2525;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16349bf17d3b4bbed752246b2898340dce9293650e7c2e50a2495af2256d6816b5a496dc5073dececc5e49ad1efb69285602b0d2848e427;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h206499b769a357977ee7e34629d4ea4289780168ae3884341cd3cf6d2c971b6b2b22e84c1cc1832b7e50a115b5ffacb27dc2bb5a2436ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h605b277aa4a7ee19a295cefb75797cdcdad860ca18cd82d7f2100ae1484c391061ee95e697df3720e4c263ac3eddbd23dca3ecbea706ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fe9c0a959257ca5300b129cbee46a29fa84ae07e1601786236a7cf7a39cc88ce580ea43b9d777fe30ddbde242aec76f819107b80e2f81f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0141dae8a89eba77efed92f612bbf2000d956b7a89d9276d43da736305a27cf94ea4c96967967f119edc5f35dd77609a884eea16785e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcbdd3a1bc726a9e655c2856349161e50a053d09e8a0d7ca7637826010c0222ac87df22086279ca3731d868dbe93d09529970ed14dfaac8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15506b94f23d3da4353d9fdd025f50c2d4f37b4690e357a7e3248df680608c4e06da8ce03bd6a90fe6cea8cba3dec2567f05f76e2bfd28e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e54bd748fdc0266fdbc8f062705f330b695b35030b07f6016b7c372cef004ece1bb74100885eed3d081a18686ecab29c5d2ca88de4924;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc7c664f10a8ad9bb5466f4023f2d6c86e44ffe661ba29eb2d12d91107297776f747a8c30becba0b2580f0c783f8c574743eeb4ba38202;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h971d0fd4baaa172415f793159b98ab411965313375ebcda149f1ddbab47c59d9708c3bacf51818f90cedef3fdc46265c19b2b330507abe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164953c05ab54ad88f541797b8174e016420b2c3c92a7e8d493ee6ab9fe0de6f9807f3b4c6f1d9cf90fe5b3bfec361646ed7a8abae99ba7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h279ec2a7aa18d0ef75933f281f29ec20ccdf7527c715ab31d35d7d9fe1c01ec358dd18ba6a415cfb7e64bfd6df268f1b0f2a38504c56f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hadb223cb6f8add4c8621e12a31e2436948b7a0ca901f38adb98cf0de081b84ca480d4cad527ce99ea7371d572ab11782389e9296d30372;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151e21e0fd0693b1b5cb1a15e23637d814fe024a34c338f74f81c3288249809c0075a98567b59b55322d2a73d2172527ae1e8f0c08f4a33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12afb4de824640f819ab84db23680f84e9b22b82e06f58e5047915586869c6f4fc19403010ad37e26155f8e59cb9c1c8bbb6be8ebfa6df3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d4725c35cfbd6941768968973a33a334a4b672c123fc22623e6bebdb2fe9e4834d8425811110669da0d207be0abf143ca1dff18e13caa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e4edde2249bd8d1fdfbb97db5fb905bcbb76e6d1041bba4a3130866fdc9c3f9a5fef0a32e6c0ad012985d36e96557b92259ba82eaec2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8edcc6c0ed8ea3e3e3ed541a58b69cb5374030279d0d3811e5e6d1a51eba353b624fde27ace6cda280c6daae3036752738ef13bf5ae05b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb4ad9a87a0bda0ddaf721403acb722c6f7c1dc2a9ebbb292c6e911d1d40dd83c4c047a562b1e95846cfca9819f532f73c93159c0d87a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cf5ffbf8cf1855f870d7798280cbafac85c46e6aa36708c8412cbe5601673104947346e4b2223374a549d9c3433c2450b53a313d31557;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1326fdc1a4e6c606931845c07520545970a64a6522af42b29aafd2829c6c470f4f19581d4b934c52329dbde87eb56e52ebace556907858b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4dfa2be7acdc9f9922051e77416222f9b77a0acbc5d034fe237ad3e4d46972e2c40621ffd9e99c805f99da50768235ba135a17c827b7b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd16a50ccb9f69aa827408df790d81113d70db1ca4e798b5c05dc41a5b6fead5af4617fc8c6c331914957546979b6ed803614b936926c81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17b54fa18cea2074e7373aae50cb7d7139078369845b5d78512178c5fb831ecee27813d44636aa9d8b7c68fa618de65992abde6ef087dfb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1074afb9ab8e3b66c1ee7880b43f63967ca26ac19c66586ba8a18fd553baaa6260c498a633d6e2f29c55c8108fd6f9de01afcffdce9376c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd0f059a19faa2cce1bb3dddbc3b527f11308f75f12440016daea2f19cc14960c1805a855dd940acfc2f748124c3888e8c966e8e9ed4f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f396f1dead25ffefe659aa658420f6529f08ff6b2d153f052b94c82769a4cc369c4b306e69f822c83e47251c603cc3e507a7bdafb9b61d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80e36cc978aefee23c22b14d3159e524a227ca9330d2c1641798b4c906d7531787dd8679b0f2051c29c6eb2bd4dbf46578ffd8b9156b87;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h105b49cc6e38eb2394b1db71b14765315aa3301ae1edd7ca15be5835f6b133c4a2d1f242997991805954c912ef107f9451ebb010eff675f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f4b0e16ca3f6d7a21be398769cd7b751c348c5e843ae35ff13bf089845c6fc6d90abe76af24a601f8f1fc561f5f5d4a77f304fce2ea94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd57301384590e09e92ee4a2175733b524c991574c81ac20415eac77f1579971a64f00284a41cb13690f2512670117a22d4d69453ff863f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee9373034e8856f5fb9fc601e1cf210ccaef88db37c3d781c6485cae9a0ea4a3cc8e1a748c6102dfa0eb7cd958f1ddd4c9fd2ba952f508;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd72eddb198aa33ec7c75f4162d4cfddb8fd26060ccee9bf1755bc3297865a79b7fbf340d0b4992f4e2e1964305877ef42d44b382c543;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h100701ea781b5c9d547c4595834139cef01097af53c39dcb42a252437dfdbcada93c86e4ac9995a340e94cc7803b1786694c33f128b19a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d0fea82e32fc5589571bc2df1027743e7570107214f4d644ecdd880d301f46670c75545bece57da37123d15b64318e08b7f4270bb9910;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h73f0f89d116f859cdbe8e57d5d24d378eabbdd0380caeaaf535c1a4807b3fa09363a5c6d5b0d79784d344c685d4a8818b4b80b6cf663be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9d159ab49992fba9d67990bd370ec8d834665005519cbff47da3b8c9e29a42ef7aae3973563db9dc10d177ab726f0cdb57a7cef3ff878;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a6d8a0c8a53cdc4df3cbc47eef4065ae5661903e80d4fe3fe42f1cc2c6ce837a01dc48410196adf4f6fdd173b9751a2e1de69533cd06c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14705eca48579c4bf2b15ad4298556d656d45db3a9ddac6d948e49a3ffb4c0a28dc5277a6514116aa0e898e175badb9beafbeb74156a8d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha034e443fda348f482d0d9c2af0a19f0772738547efbd8f51833deb5b76a6cd0900a8bce6b440f1e2744365977e91b717510b7281cd383;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c421d40ee3d3e5a1ff6f9795e8f695c324f20134ac985d6c650b1d07951679738f2a0062ac455c7d24004524b713f3d4adc56d8f766363;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69b5f9d77165aa7fff2abef89286844e38f702d962cb5e645aa0921e82959aeb919596d600c48e8e2be37f702dfe4faa373db4b4ff3775;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2bf644efd37a2a6c2989920ffd96d27c83a74cfd3759f967fff88d47c4b2677b01ea1a0be5109988a2c4d8ce64189df19c5f936e9f3db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a93dec240f9c5c9ddacf30e44bd960fdc216c254f190b44d2a8f499ffb90495bba2085d49a035a4637874fa76ef6eca20affa752089e07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e6bff14e1c00bb376fc0b2bbaa364fb109c74f57cbac42a77dc48a7f536f7258647436250f93a5305a24777664c8994c52cc7fca4b2116;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he945aca5377843ddaee147080ab5035d5521997d6912f6089db38e610d1b2d730828878a90b651356c3994a231bcf183d1da54d5be932a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5845ba50db946d801704c69810ef2d1b1219c22725ceee4e43ba0a6db4e4335ff4bd376ac7c25098edc05852966f1f4f3f89d6e66b56b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117a23ead5d78375cdcbd57fe0849924ae70ecf64569d1a591746564f679b0c98ced6068bb8ec7bb403ea6b59b7c95495126f19bd5cd62f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca354f8089f5d4f4de0006392422851c21b4aba61144c31250751334fd3a27ba4a30cb777386137f94426e767acf7f458170c0c6e791a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d5c2f5be8efb2444c4b464c12a8a2ffc4338d4450eb96e9f4bab51adfd60f7a8a782b631020e5afc40fc801990692a8e952f651fb5fde;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h113398e6d778097f8a9ae138ebd3455e2d986338fe2cd6696915149158972ca5047b1ef5feeb5b524754b47724017c7d064674a7e82f35a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe743ed64de4ff3e35fe4438e7eb4acad4608a7910985dc41eba7e1cc56f0bc11c1269a74ddaa1ee544d0c8229fc2e281cf05482e54024;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18de7ed59f834fd456d95378d67dc89bc75d76e8a224dec52b58a6009f853ccbe96f38d580ab2f9d3629bf8dc4ad444f33d6fe5d5d7445;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h21933371ab198e2c2bf4c3fcc6eceb97d95fd3b406ecc8c357ed7d5864cbb43d7890b30e1722c934eb5358d865dc1c7050f3172c511527;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb1fc682ea0484c52a17924ef1360957abe5f922607b776739ebda214b0fcadecec73d5364a9082561c12c56e91f8b739f4d8fd4a33d35;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198a1cba4c5752bdc9f6b2e8ed8dac4a61b50502a5eacd6b35ab8ec6742921c906fa590807247935d7857311bdec8442d463540b19aa520;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94a1b4e84e80bbb46b19b2f26b11010b7abc8c81a0e2d694460ec6f3018c14d9a0be08862c42b9f7f710d18a002a7d93072c7a92c086c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5b57cffb851028f41f96c51e06f0a806755db025f8853f4c6f5f8ebf99d0d33fd47bb83074e6afd02be72aaaf9495dadd4f7aa98a7482;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h169ad5bd6228320fb738cb9f4f62d7f30f401d38516011654414d6e67a86bf20ec6921c1c33c710ced97128ec0520262cc818bf7c981ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cec3bda610ff9cbd07df2235746ec2a335d45c3551b4247e6a930d86834c30ccd9f1066f62dad9e99de861946bb2d44b4dbf8b2b25be55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd963dc22a7635abaf0cdb023707cde0d50100d422d9501123a00e16a60acfab0fce4597c88665ac02b0577108af9a16fa5c229f3f0c49f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15ddebff681b2cac196901af50687d3aa8d767d495c444744e2e7fc9a93a2cd3a915a586d8654813988164edc11ef9971e682f488b5a982;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54c17448854ccaeaebffb96bf3456742b53870a7d5cb88aa0e5a81f8390a98bae13312e070b03bc2174d96c7ac3f8cdc3b5fd2f2d7e1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h163150966545a1be95ebd215ae80b1dc505b4080a564d5d47c8ab4419c4cc26f968a98ac846d893dadf5b3474d860da0e2f350bec0242a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f64bf731c8960b6c53371807b706fa3b9cd7cca6bd09ece460b970915db1c4157a5738066b6a914ca4a08f9b1aa24bee581fbfb97761;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h139cb64b697724dc0a9f0b7a373bc94cf4e2c415cda6c9e9b32176eaf43b101f2d4c6b3c9cbc409e381c599f679ae9bee36477beba1ec3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf4ae1c68e7a8ba306c4b8d1021ffec954d11b1640b1b25cb9a6b278e4d7afe1f3e4d1ccb3ec9a397a877de1113cc01078ab36699e98b2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1457341f1164f2a06d140643cfebffbda34ebf872a6dd7b05860a7effb520e71e35fa2294b2a5cfed8664a9b27ccfa942cf55e49210dcfc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b27ef351c0dbe58dcbae527594afae62e51e1af219a6994caacab21716fdbf02f5d541b32b2603268c9a5933f629f61f21c7c1c679a6f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h235a72f09ac8271bd7debc8505654cd3a95811732630065ea37e5cf94bcc2c994cf7747d1b0ba5a822e6389155ccee65ed47eb81eda07c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1776d788f455078a4fd1cee5cde79d8ce20dddf2ca171aa1b1f5bcad39888c618ebcb8a21edc0d077a868f4274ea277871f5a4bb641c45d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc8b090c8454d769ef328c568fd89e32d937cca9fcd09a94e34a9859c46c7e2791b58688ec1412b522289eb6a9a67b1847aa85f1cf4177;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cde4939ea38196fdd5dfd9b0ec1da45374d7aa6f642ec39bc36aacd891b4bb8950771c5e4874153dc4c9a9bc495e54682d4915572d73c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hca027a5e63c2f210f1a8544d2d365b117c365306ace49ed8cdabc9eedbe66d2c65315bd11534798e4bf5fa376e4b19328864dfbb9549bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5ebfd1aea8e1c975e82a4541e2beeeb2523a6315abeb67aae18f2f76abf4818e96bb95d00ab9c4c6c69beacb9d81eb7c29496d37ebe961;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h83042278260a99751fe4ecb4a7958f2a921edca66941e9e8254f627149e154230330341a2152086ed72e51f7fcef512a06452a89b1d1a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eca8c74d6debf2debcbb4d8a31fb3db10c4bf3f9b10dcd530a94fdc6f8ae8a210fec936fcc2b1ce28da8529fb4efb9ac686f69e9c7e09f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b8a588704013ede4db07395e806ee4f32e1722984f25fe6eb117cbaf8b4fea570ebf79f5fa1f04416d79058e57508082bc011e0c5fc47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a144c747fbf83ce163602d3bfb9a25d99a5bb11d449e8211818c4f68ebfa94bb65006bff59ef73d9d58ca6e7737f819413ff9edaecb17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h150e519728d4f4cb54e1002ab5feab8cc2fa0e8f65706683a9ac4057b1c2968a210f0463e26c9ebc271c2bf36c8e421486c742e01a847e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2f76a08aeb7b86e7373d7ae1b7eb3c376cbc02ace2bb8e3cd77c51fa6130066943ac5a20c65c27f7a9c39c7d49b7935f8822fb1d2033;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h41295cfdc5dc118a9d31c707d38ddafbdab92a31e73a471f1fc1ec3b7ca5464fa2830096bfb6569aae63bc6ee7e8834485360f5af77d56;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13baa5223983be3406540145c555068fe3b919a9a85aed6958ebc19ca69aa9a25cc814290bf2e78de756aa37ab19fabdbf511286e3d1687;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15bd523fd5e99a4adfccbfb25a9050a340f8868f15fb4f0a64ba1b4cbfab0463462b062d71176b47c4d9ab1015b582f6f40ee91b300f48c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfcad1c28d23f4f563682805ea40ffb8fc74f7001e3827ba9ae3f7aaded5768f68a5147d859cfb8935a56f5569987e856b180935a19e157;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7121b5b055003cf57055ef4d9a8e8e96a562c83383b6b82d3175cb64e872536c1247d67f8151115b10d3c2a9a0bf9eec6651e517dc8a81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h147d96c250113430d7c850b2c1db98f1df87302fcdf470769c1bb27f54495229d88803add9c66acf797464d83da0f3615a091400fe5b9d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c62e7e1a2d4aa3d6355d7f8f843f991bca27295ebad0db650679478a750b593df7bb682fd076b01ba2bd0009e52d1e4b4b68860ef7a67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc377cc26c337368587a71ec52ce6ab9fbc6f6bdb8147f0a69fce25a15bed89247d081abbc608d04499b3350cf44660accb7612228c2886;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5020b5b02e62e6d4339e3ac21591d7ed5730a4b6fca566e2ecc10b14ee701533c0282449fe063c1d48606f8e10eb0f6fa8b24445b6665e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1627b5f99cf714027de5730f8e7edacd17e90f3f5ce7e50325bdb0ce53cddc4cc6b473dbd86523d359408a10b514011f196ada24c710fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcdb836119ce50ae88bf2c62b7be6332898714286f47fcb713d6cc7832c77b3a3a825a2cbcbf38ffc29eb689ed07f82aa73e1de1831c7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140ff59833f0846b9f42fc8dff4dd39473b3ab2ad70034c1f3c88ca96bc91cb569e814a564ae12fe8678cdbac2472353488bc2d3187c25e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h109ca3b8d2af1ddbb8c6169d6682e1cc56c019954389ec46932eeb06ca6c208345d223da46a5f39f3585dd4d67456b027ab70d3705a97ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8227da14d8dcbad04f50f136d938b9390ca9443df38cfbedceb901051761729ae4fb465862909088f3166f80cb108fb3eee416c38a7f4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a837b2aeab5a6d1d48b54762a309a2750b1f8776d46b4d88b46d97b29bdf109f963fee7067f00d91838d4ef6fd717bc985e25416f8512;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11fd30ac7a929fa830e85536d5b2648cf0f564f847fe5879a8fa168c5aafaa504099e0e8bd2f11913f1c5192b4030b48493ef4da5796520;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h44a644b68ab842f64d6500f6343788407f655710d3a023cb89796dc149cd42a7bbfcebd103b02084ddfea5813418b25b522b2adbe509c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h591d550343a60d41ffb5716d36b23556ebb23f5ddd8ae47d940c743017da5dea90bd07d46b5d433903483947e9ed86d070694eedf61cdd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdcbcd78aef12bf170a64559c77431220de096d11889343d7637e78f28d744afd0755d87a4200d0d9c25bb314b0c5f656af05f2c710872e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5e77ce8ba42e5f3d882195efa35834714c87898076c49d1a486ddf0cc35c4baec082bc518eb2ec62ae2594adf95d79be745a4664628b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2aeb450ec71e3ed96f64af28ad2c57d0e50c484aa4d3cf8e56bcc66d30d40f603fe120b9a61a19487a0ac164723ad27f10142436f7d9c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c6bb289f1203239f5f57dc38bdb954edb9e6533aac267a7ed788448e563e79548ff1410ae6c9ce059b69defc3ccac4834ec054ec1d01b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10a102c84a9f15f2300396b498ccbee265194d0abb025fe8f8a4ab7d71a86116d3d03546f74efce56c5b0a857ba85fcce66960c0103bf35;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18f9208459247830817e6dcf41148437ed65d0beed1e12e4010608c134d987f84a370df764bc986efd9c2a8559f70656293c5049e1b0a5f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h137d869748bfe82db1312853821e23f35cbae02db4a7fe1f68dc4cee9ee17ba528d041a5078e9b07d4f69e36f89d204e9c95b1481d40a94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hffd7a22c4fd4a53ae2b949924174444415c744a704bce524c2bdd82c7f64abfdcda4d75592df15f9ff61fbe876b4261ee6d67c9edefda1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h20beccd63fc2ad632a1ff65e8c387c6b304544fa19d258d2aa785ce3b8854e85fc59d5c8c9d1f795efa2b8e4f39ecf6344f166c4b5afdf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1968c1f044e94edea22c619a6f7dfa1ceaf8150cc7dcac9fe00c6d76a90d54c9bcc0234645fcf39156aa28075afac3b1d2838e5efb6de54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19c71504632c99b73e926885f1607259f8340d9deb9e1718aac9d23c2c7dedd73468948933c69ba5c961f347f476601c93e4b5f2faabf01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3cb29536e5a1515d40006be01931555a271c1fa32312bf03aa9a2bc8aae811450a8e4f822d5f634a0e072d5eb80ee2f828a4e1763ab86c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d998fd8dfe616f3afecddfd6745eb4b1e158e9c43273338a5e0873ce764275f300d5556cb1650ebc4dc3b3f5b949fa063ec914703bfc2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f777f4e71d23785fa52f04536b66abb6b3605b108cec696cf3dfcba103d7c569f34cffe81748c0ca498daf098b4634df72107dc4f59a77;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc52e69967dda49d54125b460cc67e84ccbf9624c3958a21aca7d3a8fac9bf2626f390df759607b1ce652c29fac9321e34445538fd77d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h86a74338de0019d2232d5d633c86ae554e744cc416e3f811da155b237b4f742beae6eb5faccbc567dc2741fb968943808c114dd0a5a030;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf399b8c395a5f6f19fb9a58e4d3af368b10334988d7159843bc6a8d9d392ccc17b0e35027af5770f1174d99d245541d4a61af58ac9298e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5febd6ee7b9d857e1591fd363058f6eae845650d189704c50c2f5e847feffb7552a2fb219c3ce18b433f11b047cd78fa4d1872f80191ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1daca26a2243caf073f427201679242b8a016486ceb24c2506f802f2c634f07d0abdc934729565c7c5cc907c602be71373c9fafcdd5ae0f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad98e51b5c36d61e6aa7c47164cfde1eb7224ab04ef264d83144bd2f524b3d021b965d0acb9b9115b6eccdef33fb206d4611c108f5f03d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18438bbe387240a306fa0405324bb7a6852f3c627c2cd619badc06ecb56e60d43bbad5424dd6821701d8b13bd6ca99df3d98cbabaf75f98;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc86749606fbcb0ea4c80cf519654f1704be6ddfca903b32c1d9f5ede6f8b1d7ae30b10bd42b5d83363e86215ac90bf62aaa1a63b033fb6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb187372fe6754bb04c5a82b7898d36161cfbadf22b981d5159556638904c4d50f0d32245f5c83b5c6dedc618f08f08424e5203773faf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f02e0d0d22c8a40ec2776d0b79458835fdd33e633d902d5c493594d0e83c40793b1ce386c3937079029dc6e383dfcea5756e5720aca912;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff61bd239ec6426d5012c4db6e1ae545cbb9a48b36a4422696ba554d4f3a5a69b442d49a3255452e3ab340afc64ae613fc630db97fcdb3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1656fefda65a4cefc5942702e59d63bc382e91021b8347b3600b9ddf00926b6828b026748929a9c069ce00c635243ad0f39d881bc5b7432;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h136562751371d2e14483f8f870755cbd4632874d09becd64576b33a23e6e729fdc24d4b7c4660d8f18bcf91788f2be9ca619d6a0ed24eb1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181b42f578aee21e1f06e20e20fb1c6daf0652b1f708409675c20614c7daf641e7fd445f8d2fef90ed7b2254f20e96800961d2622b8aaf1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf675aafe2c1d72405a870aecc223db1611733da2e089bd70f001f739572d51281ae9ab79db35ebaa55d09f587f0d12a0e466bb80e4d4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h98eb0cb75289e6adf5f62f909877c74fa397f0ca2a8db29bd8d960c80a56391d16240bef174f2a2a26629cea936ab67587230fb5d5fac9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hddf5e35fb3ac3c457d13cafb559b4deb8457370d237a3a9e20732d93784bc2a9815dcbeec72522197a16f2d54e5e652124926b93c5e917;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h34696bcc68ca3fca96881ef84cfb90d313cf02374840c122df502a5bd5da2ef5a725ae650fdc30649656f90494ffca9064d2136d08e0a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a1c94c1f8d914ff1f0cb072e58b506fd89f243687827558887afa7ebcee3728ef3f780f4f177b4771c1f13262fa8f00648db10ff2d06;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a6a6cc1645001594a4f631b0942eeb21721d871da5a80506def1c218612ade4d71c30da365c09281f5aa039486ee740c52a0c0765d3a58;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h91221525b8da93606a5a78fd7802eaef1d8aa73928f50ac5e8cb954f1001f159303e90fb4ed89831db0aa374d98bd8e92b0f09768656b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h53f9b64a3a12744eb55d62db1013fbcd6dbfd3f0bacf3b39485963726144e5865d9ea21a33a41eb484c61164c7212a130768d18088fe90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7e5108c38a5a59e5353d15d1741cdf8afafa1dd1de79c637aa6d86e695624ceae3526ef6ade33b2cb2443251e5a10ecf7b60ccb6e1a533;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3494a7e86dd5a0235394f1a12f2b6c6ccec49db943f30b8d7b634b9d4e7b71aae4d4fdba77c24efa6f37cdf2d8f80d7bb058d422551e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16086b66654b49fc0b8da582087bb23c84cdcf85c900932b1fc6a0158cb3344b37ad3260713678798c82f332049f0eb6ae988a3759fe04f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14d52a54848c3138a86ee319a3f306422380a782d2f64ba9576e42982124472e8d62da0254af51b77acabcd87461b89643b83c7db9ee09d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1acefa16bb96aa2bc78ecdcab4fc42a08408e21bc777642079b92ba59db980e9673a31431fa7945cd861dd00585346be63f908da431f1e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf70f5c32d4b81fae8e8ec7cbcb959e5bca845609b3d49e2c58958d96574b7e7fa960b32b3066882f10c645ce81a23495aa01aa74211070;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1451d72014919032554cb1c7039146df393bcec73d9fd7c32bac9d5f7aa1f7f901e50e95c11c8eabecad4b32aa215791cdc9e93a695b753;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1326dcd4d1705d724ebfb9c65246efb6993096220a5ffa8bbe5ea2b40db22139ee7921b003d1b715d95d0c3217894f5b6b49a9db414a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb16df753f17e02907249ef6889f4c4f37215d67cb16b9542571fd78f3ee81cc15bbd61eb3cf93b83955524eb1988bff18e34037ec9d00e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d3096f12923d1bad9d3d7f16ff3c29b6b080c64a90420d152cdce7f850c3a4277b4ab226a192155f7788ca62ec886df860e7e263faeea4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c8b968947dd1e0a43370d50673f9d02e6d0a5167421eb11bbd299bc85e721941145a28856b2d7e0f18ccdc91c2ac322c6f33835006e8b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f13b2b7cb6bcf30b4e746b6e713840af98e1d9c23be6236530a209b4a4c2fe7970a4f99a474c50af6e23e8913264c60b3fbc7228d5abf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h171b6e746ada87b744e98e6825412e5602e7a7c593fd6ab3ad6922f051aeaf8f1a945c1f729011509857c8c6ddb3b4fffbb3158a897a9a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164ef7a9123c9bc155a1b96632fc6450edd7ecc5201a40b73e7a1fc011ba2a6e4acf8e97817ee435736960741b19a50bb054cfc229f1a7e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h168f42b2dd56a958f451c58dfb36a4076b86583bd860c9abefae93b712ebe50b55e36c6a88a7301697f632f23d5dcb044ec2f30a2609e05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d38204ff619b8d8bfdc482b4aa541cb5166e794299267f3afe96144ab28856e95ba5db714e7a3f51a66d2d2185278611108c55e5859a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130e87259a6a4d5e5a530ff6f9005859685190d7084661a7a622cd7e3efc0e451fe2975a4016a6500150085d237bc920c822cada2175994;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h42c32a556e16afe9db7895a3d0f152bf0f8ed465d4c68c0094b663beb53dd5d2731cbe1d64a972d2811d3a0fd672ccf0c7a723eb672a27;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4e5fc9973c03e1ec56cc038c08419aea3de3d4e1f2e429568f7b6c3b81adc0a7a614090d090da04ce57490f98c31b438596701211c2f8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164058b01f8b709a118c9763755160ee829d9a0cdffd3cf17c9ee6872ff5430d61c5bb9e6d46b7c8da7fee25d5850be8f6147a0439c45d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd589c33a5d480b80a858000ef18f14acfda6e38bb21f32e3e3cc8beaf1cc540bc7bb94058be0fd07bbc6bb34cface4829526c634df7bfe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a5b8944c43e894a6dd3c9e53745644b2c780c569eaa7161244a8044491a9272174d6f5a5106fad9f9bd07b115598dc5cbbdf20f88433dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h163ddfe01f52bb4569f489a786c2dd36112ccb2e12b9688a46d99099291ef30ad6c32ebdd7558800b735113b5e411e5f01cff7feba8ea3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4d4e7787d9aa0d107d7618f9d3f08b5a44534ee954efdaba4808d6516296a5428d5b6801931fee23314b7323dcbc871bb03b135286987;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h42965324b9a9eb4b1cad4e0f289ecc83540d577935ac9de477b5c73a5dde214627ef460257f90261b5f87ebcafdd0b929a7e2f54b1fd9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4a98f17f652f38168a0b98b362674582613388364a3c0a91ece99aafdab8ae6e1611368e11081d75807bf6136e8e6050aac973401549d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd818c192cafbb7c5d0273e666e457df49a1f6bd8a1d7736a90eb182543f794c31638817db9da3235cbe7a6a6c4b01e6154f52b0e5cb05e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h148933429b94a1e5b8596bf008c87b34a06954dc44fb3aec77f1bb25a23203d24714fdcf482517413f8d51c51c38ee3e40a8cea343a98cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h87760f728319e73964b74516873d26bb9ad2bf38578782864cbf7c1e4775c44a4b0a0a926cbf485ec3e44407830a5f061d2f4a57ff3e5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e39d37d4c3a0f16e09bf361a647b278b34acaf8d5f233372f97379e8a30968d7670a564f4ecdfc81c3ff9a11eb7172ba1f15a58d9f1e30;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfe922230aee4139c3566fade96f6f32e3f728020ed908e7a75fe8b058b11c810578c9c2c1bc656a6417955b7d808919e1800c461ef8a0a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h288c376c7c514b6385e4a45b5b23b7fd4d039c5a403bb22a60a02012f08d5f2e3b99f1005213861ebd37734d45422a291a14509b00df7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc4ecfe18318edc04bc1d7b3ebe8236c67eb4186aa803e35787be5ada5ad49af8d27b0d4890831b7e7dff760c006ca5e65ca7aa256918c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1748d9518d7b98d2f1065a8fa86f7e79935c996824c2c79aae48acb28cdccaa5b576fa3641074a823c0a717ce111c408925ca2dab554e64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb26bdd4c9378e13f2eaac1fab12fa8bf880a44c6add3631f1b49dd4ec84ec2cb1581d4ab69dd18ae4123a1d4d7910690f745c01127fd2a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cdbf34b11b61ba44ea6a5d13fcd7c32b61d430f55dc7276f19eb9d5a0022c0141c912482abd77b71f4322346391ce8e1394ab65aecf0ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b0f4a6f56c31de6ff67b2e6dc913828d9cb5f6fcb11c74d17fc7bcf20f8577b019ab05ebdd1a61f3da2ce5467b3399f6dfca92438e498;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h62a20ce46ac64afd38ce456f1a1e868afb4624484164853ec7d452ac6eb72d4ca9d44bc08516591734df5924af092b069284dff927b78f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1844ac18690b3a2d7588afdb974db27ef4ccdd2b75d04529deca46040b8ed0505d4b9d6c944b63988a5e44e82cf785f88dc30d89c6b83ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc7d8db441e9a38238f8c122f005c689fa369af6bf0fc5aa1c848a1e751c1e816314d96609ac9e5403ce60a7862e7f3e9a22029d79a0de7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce683336889e7eb8c592e851fc7d2c815a764db53a9b6bcffb306cbcf89ffb21ca6a7208efb320386a6719dc3951d5bcdd4b4a879537bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h125b90a7e5c96bc5db2a4778c39ada1d2fb754550a3695cc6b61fa56e37d23926a1f6e8d4d7cca3c597d5be540331afba97be20cd381c01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h473c64d67ee119759a375b21da61ea5742859e674a9f1c9301c1c56e16ecbc5300aa64f1b6b6d2e0980140935bce9e5f1e265cfd3322ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5ea257bd0cbb312df7ac83f840421e7d381885c6cfd175c9b0f0eca722091a252de7f4843b2e1db40187622903d5c5943043bdbfaa42be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d7a9bb047747287f2e633ee489f3226665277d2ae5d777f31c2ffa83131ff5ceca77309dca43d4822a0d5df602a2cfc81d88bd7567697a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de103624aea778da4d79ecaaf699459f3d43ede491c3bf76eb9406500d89ca76b036b18b816c80e8200535576d611e3f28567eca0c56ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h910ac69099f5a42137feeba0bf4b8c04dd5a4406f2491a781b2571e294938d51849ff8aad2fb83030b921e275cb73f02fa2f66872fbd0c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he6c47eb8c2402670fa140e202b31cc1c50bd153d71b89994e18276fb1cbf3af967feebe0ab59a5c8887b4163d7efc34af2f989651494ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1061b714d7870fbdebccb73e7f5e351e2f031cfdbdc23fe925d98c0163262fd665cd3ec82390aa28300f35ecc79251c1c64cdb7e3e39df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb4d5f2d166d0546b595312572713167dec692da610bf500371bb405b548af33299902e9e34beb15a4639a3e9150882127bb18cfd4382c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h52d5268c34ad216c194a0e103d71ffd170c97747ec72de792b1364b78fcf70dddc52a9313271d1419f630405bb33cb22be77ed592dc741;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8903df0f4ac6a9a27368da7c4f0cf055df6c3b9ec8b20fd0bd6a1c119202044e60aec8ffea956b54d6c1d5f6b5f219a1bdf274875d65b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16b814692a3bb54ca78dc7404026d34f5c5db08effbc4e634cf1fce76367149ff0c3d465b029fcba2074f046241bb550b94c0a18c85c599;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b61ec45f0a81ba768db218e8e04645c01279b217e28dc7ba308889bc837752925afe80c9818aef1f9a7eafc01e52e9be5e3a993bd71d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7696ba0519963307de3e1d734c0e5c663d7b5ad50a791e12c9fc4d891aecb7cf7c01c56b725d5da1d9697efd74720e697d4f37e12fbf77;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hce80fd76451910bbf171149ba9a09e52aa26eb9e8717c8e352e4261338cf68ae55f2f9a8bc6b99297b25b1a252520b8e4261dce56c8341;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h123955177e21a3c1bac4aeffa70bb1f5b2bbedba0a420bed445e927c6d8dbdcfc014b77e77f7af69f9b8e50d5e2c1b7c2934bd390cc28f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h135dd35e99a4160d1b0f5546da628cafad745fb19b38cf4c04d86e3fd3c53c6a17ca34ca76b8df09036613dd48fe33da6abd33d66752dff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h420f7e13d36989307e300ce643c8a588219ce2ccdfa20fd0bc50bda99eb1c653f1dad68f0cec79f12214f44808478d558077d9c4bc3036;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h693c07e351ad7e2210e0c00182705fc4102d4e1b855bc88d4bdabe8d10153cd8d962061dba8353260238e096d43f1746fd10f2a2618c78;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hac29b3862c706a483a42be1b72168e46fe770130235eb885d70a3ff56987ba0cf91b0df58a8319e6979d4f82f28601fe4130183a93fd35;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d1bc4fd6314420d4652f09b50c3777d6cbd6916c4d209050e7d1bb2424631ce862285d0a41d87ac977e5a981341f5cc793cdd2246f83c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h22b29643c6eb60d9a6f1d373a2b2a2a50ed1dc89965e3d4a9b039343c7ce553ac0368e615f485eb5dc4c2525ff131d58a58e4b1619afb2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d1d5090fe4f037ccc7e307f6a2db84e54d1eed4700877be8bf0a039d18ae44a93922564d20769026668ad78a875cdda72edd2cea1ebe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcaeaf8308b663acc06f3fea0d341a2c20fe3dfcdba3b5314d96f4a1d582bdda617ca3b3b47e7984aa1ad9639ee8bc23f2513ee37ecdc43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ebdcb9242466405df22b403b0ffa0843d40b4c8c5d39c60434f5603fa336911835eed61f4c92f1f78fc637e2e090e5baeeafc8cc6dbfa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc3a55e57b9039ed06e0cd2dfd86e62f579f9d5724245797a137fc26682ec1b014428b67bfee704e572fa84e80b514d47828ae6b21e4b02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77626012a4c78966f3ecbaf6ee0bb4966451d7d159a20fce7b09f2b52b9181fb64180294cd54c1a3e8fa4839ccd2f642ad6d8e2b4f26f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9fb3efa0b68704e80e180d3e6d561bf4a65c69d3456657814c87ab897017149011ece2d186f692c23875be4d033d3bc3c86398db7d906;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hafdb5f41a2366cba5a4f32eedfb3b72f47284024edf8bb9b90819cff4352052f3872a4bb260280fbf0a22110f603ad83883a4c7efc9ef2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6469f13b1d99f5bb0c7bdb813d1ec35203f9fb71705cc3e99b3bc377b2724b01ef02cdcb5edf5a3bce6492ca79dd2bb3aa86841e019a8c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h57b54fda661dd1a7febcee1670b0545be19ea31bbb948e4ea38e48b30ae9a2d59c3ba84cd150084a72e85cfa5425dc16c5df3ec5e376e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5423418b9b48bf347781ab6ad54cb7e3fe46a2c4fa231fc80d17e843e4f72e539329137e38e9cfab2d5cc93a79b9c503f8be9f5505c50f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cdd006b0d0e58960fb7503ed61d8ab4ef981156d41b7b42b1eb921ff06715544a59a230c73769354fef317ed2e848d71feea22879650e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h121a0f358f1985f38fa2cea973e97a7dd879b0e2dfb048f11738c55467c9dac22028cd848eecedbf6d07f5a154bfa05d8220ddc25ecc7c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1df27a06d9d52abbbc44b0835ad1a944db40e387e469fce42851f748298dddf4a2025cff0c4baaa56e52a521860be7e2ff79688fd40e4fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdce612e114acd638d3165e0ef73dc5d3f34a75c04c562c758cc3081bd06ca47d8c64ffa7527e6d5d88fb8e41de3e50554bba82795f4d98;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h132769deefc511d53599bdf85e3ebf0f8510e19febbb07373fd27e71cb7651b3c2d07f75d003e7a354eb7183184cb6adec7b32258e4d445;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d9a967a94dea617447e9ef71b2b9046a74d01fe8e70c4149b48b0e083f209bcac89dd34c08b046cae60221d97cdf9c1fc8b57f0aacce2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd4c401450293cc3f49bc1d20d8a1b743a0276b74a78e6c5d213d7559b261eebbb8a71f5752d3c62434b7af4c12f08302e81b7b43d7bde;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bca7bcbee6ce42ec6848b4fa1c249e8fb7313630c409cf43974bcfe21d48682e811eaebd5c215df49e2dff47388c8de6aed4376947dfff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1403e597432c4f357c879fe0e7fb42af0173b61c387863439336f24b2862a3ccae9ed79c45365492c309189ad1aab6bc2b36119ab4abaf8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a3d773ee8207541ee7601abf233ee3efbdfdc6ff9286c12c3227b01ff50e1cf446f5c775d1511052a206e635fa3d6938d3d046cfd3d405;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8da2ce3a06b287b95fcfa2e572b26d7a6b8898ee17ab4c0768de7b5efe86bf165d15802162bb835abb319058eda120e6c6d939ec93f76;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h37fb66d6f13dd3d94eb932eccb96d0f43324f2fe8c118dc6f1c92bba99f9672564c16437c2659a25d04b5b6060f21d49089e2a1a91c578;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heea7486ca76429ccdf91ec466906faf586284f8db4bc079cd4f43f46a8f4985cacedeb9c8792e62d8197a60b102ffbb0b09b8f0aea0ff2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf3b02905884c550aa9c589d1bec89968b645b5620bbf8c8a7ca9f8e6a32e77b3bf983dfac2f2cf311860a6eab22bdf9407877711190a54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he5a842bc1d6764ae92360937c3c1b5fc4a404f4f3551ba1714ebade77e133766244da19cd3bd4766cd5580a1c3a6aeed03a72ce2ad41e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h142dbf16436c1ae142ff438b490feed3b2dbefaa3e80dd437433f4451b74d4c2c9132199921fd43af669951fc6958c8a6595c90b3bfd341;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f8c642afc1e72c4904c78ad8a4207130062232b1b15c286320772fea1cdf9562ab2a5d546e7076d8f60110774b44031a1a123da18bba9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab6a0934e040741e483298f9505e4ccd4938edd18b05ca38dbd9c4158aff3c65e2570b2ecf58b72f71003a961fda96de7c211a205dfd52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18e804857d93b678e64fcd853b00adffabc66b564223020fb673df667ba1257e3e858a45f1d8fa6fc569abc1d8dbe9c461864ed833d16d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2882b1a79b69067beaf31ac34b9166c49ec7f40d0f96f21cde4f0fdb1d72808878db7e828eefcbee9b4757a193d48d5e25181d542f3466;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc0d212bbcf9ac38379e85698e493d7888b367d41e182be976aced7dd2a40106e202c97583e6c470dcd625774d192966fd8337cb8b4fbb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbd4eda7c96f5cd940aad5ea9d12a83bae905049b72207baa12b81225ded89fd843b99cbacc7f5935a6f8f3e103b77014dab8c74ecd1d02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8600658884fb3fa368dd836d56efc332869f8e69eaac8a08a8192f8f36817655b30e0ad126962532b9d942307b374dff60a68b3059a74b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha3359d4dfafff5c91c91b8c5c562ef2e551b46e07de92c664ba8f1f42f5364bdb2e9dfdbe6b1c5249f55b032496c020392b8c71ec557f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed1d8ae188de7f278aaff5534a3eb14262169b313f5d981cc1b727d61c213d141e4b4b82345b1c0fc4842fc78274d2692672c6d6afae31;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17cefec9fbbfef7f4b2e6511a5f4b4b8c24114eacb3072e3081c1cab6faf4fc70bc5e380a850e9364758ba2bd8628f75965154236bbcd90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bcd34baf5123d84806abd33dae0a07e2d20661a9569907a6cb2e651fa3586a79fcf7d71d8bc96239ca73ff655f2463c3c7e3af0a3e3605;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c866e46359cee6f621bc50341a0b8182718a978e6a4637fbedd2d7bf3e42c080aa4ab30c0a8ca951157fab6e9bc700dc66e123d7ab2f7f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1800f196599ad3885f63dba3509a1049db6e478181d5fd7f19da478404948f555fae0f59cbc88e7ae2337a5c2d63e99f547c2ce4cdeeae5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5a99f66d9819780a9cce11fc44eb147f57723a32fe89c373887255fb495c0f680e0ae0209d924b93345029201f45937c2c2880a2f57eab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c9f1b08c2efc0c7fc630a215fb8dd2b6fc6a5225770dd451c642e2911ae9eb500cf01a87cc385ec6371bd0393cb7e578c48d5cf19d25e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78a54a828f788be00e897612ccf693c5d8adac4b631a7013442dea7a52af023195df7a87824401c9e976c63f17ca85a734d7e32d0cf545;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e22bc1437238927b4cd803aeab94d5b91a0918614cd3bb268aa5fd75a82e2a379b13a8ec7cbc5e4d5403a3ebf8327b89b88474deed67e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7290ad1a4cbfb1da93f81d674d308f3bb7a64897fa8e283ee6e1f4e7b90853ccf1f187c9b4939c80b788ee53812fb92077e59c95e65ac6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb612a86428055d604cef6a299a54d2ced66c0fd98fdadb42cd113914787407d7d7a6b0681e3d5eaf49b7a9c252c26f0dc9efb97e14ffa6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc4b1e924e21e6264734753f65067ebeb1d11e761238976ad68275f378ef8e8a1e8e97fb5e98f277ea7e139e0883be938114cbe44e9ac3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43d9f10be9cceae9df1744f8342ca68931079cfdcbf3b627787719f884615ac8e71ed6e74df7dc9797c9a7b14e4d39f2cacf6a342e0ffa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6bed53711ac1d3b2b66b33fe22f1503bfa2d430957659a5b669a12b047ed7150112beb086f1041452089f615956bd4ae2c29d42599f57;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9d5e4f87f1434a26efcbb98b941a3ef72a25f40cb559a2253a385796ab3e1c5d449068bbcdfeb84fc94bfc70967bdc565c061fbde3870;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6f30a9ea7cc6aad69820a81ae902090aee1e3e64d7a539b386054015b088ea59215f0e1096a6e5d5aba87f47f87c29cc68a1f353365ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he38d8e567b2d13142461d400bfb2b7c7e38b317f1092c638932933a5024344e8b6ef662f0317d60a2f2682827b962f22cb09ecc885e008;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77373a5bd3b92c9bcb18ec267ef8190ee5263c12a50f9bc537c87df9955a15910d6a85b1081354bf09bcd132b8e1629a25df131b3c2294;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h117f3deb2fb667dbfcc532c9c20b3499aca606b70f38979768d1e99db04783020e856e481a9876c85c60db62c6df7baef55b47f15685fe6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4332f4cb00280c074a832771f5a43191b422928c473863ce72448fb243cabb46a75f9f8b0c4b2e6f98fd3d316412fd3b5202ddaa4d6021;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h65dbcf4fa36faec40253cee7be8ff1131a5eb91a023ac5b7d5fd06aa5dcdd974cc0e4b1887fb54e4d641a68e4e878a626af94533ce8848;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e767fde232fe33ee705b99cacf7a1b2f913a860f10cfe5bfcc48b11d29fd2a8d6934b52401f6e7a6a9e714f50979275dbeba85de9abe79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h23a9c954ed08bdd2bb0913fb763add0133b59b51238b47d248c52bdaf3b9a57eb245adfec1280f4062bdd3a11773d878832d1b7bcace0a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdd3c4d40fa53377ad43158c0f92a086dfc63a63690efd857cf184aa8e627b76250006394f1a51dfb67ca3195365393032a3c68644e60e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1daa71df71a4f14ec6260fe58f10b672cfad0b9538d8d723826feb18619e0e140c0682b3d4725d9507e7ab9fe62fcc2360c098f337a5b3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d2c03823a914f6ec1c893563d21efa7d54880487dac705819a12ddf273a0ef0bf8c6024185f248d95a13e8a9fcb5df5294d344421ff4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h55f3ba2b16158405ce514605bfe6ea959eca496273254d9a6c2e699c44c69e7df00b383bd2db408ff6736c9e243fe139f3794c6072cfcd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f95ec710276c58cd79af84a4832f330b0775b9fa66de5f93143a8bea62ce1042b0d82ee1d405c841b9058b0003cf75890272eb08b0b23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h32fa23258b9bb41fa0d99eabf8f1ffd14c533563a9e08ebf1307acfb9cd4beff0fd1df8e333759118db19749d09adcfe00b8f872235929;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c92a5f412a1333bb737829800c7fae486e47f540b2a08aa8ed7c84fcb1e3a6453e6ae7e63e3923efb147924a8c5026ddb9818669530f1c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf264961728e9a8ad92eaffb4f77adfb26e5e17c89c12a510e949797d28079a17a09949c6fe47c00e3dcd2e5688c29966326014cc67704c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ec62d4c5f70b8c7aafd933c2177ada091a418b6e839cfe9f62896549faf4960104082a030803a5326d10cefe6efe848a8ea93bc289cea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15edecd4905da4a4d8f2c3e4d1e0a814dab5414609687d6c9ac94bf5b79ec3e22a20337587b92e04fb926111f200d2f1cf4959dc8797613;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a7d9e5bda1b0a8a2efa242974c74d7a052252c05976f59e24b0c891bd77a5b8c29decf5921ba2076a6beed05a6b83c6f6f1658127e79e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dd17a45b02c02f0fb7c619749869dd104421c22f2f09cc50b66fed595b40c87e9707d980acf27dacea8196b892802413cad4a619961007;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6077fa1e5f80ae12d3ccb4ed6cefe418637ff8a86563c1cecdd4d885dc72f65b3cd2f1a2be07017ab7b9e69f46181ab44a1eeab4a1cbc5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11907c36c1a65daba6d41a9b4eef7deb4e3b407838c6618416e3a32566006bdc0c9edd3ccf877f73eb2fa7ad4c4ebad3a7142af8e0d76c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed9b54a6847ae64701d3f5ae3537038dcb800e7dc45ae37c8e6b8f8cfd837a6d5af1cde8bf797a632b3f84c96b7f598830143135f7f811;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149b33591ea338b52cd0b2177672d957ea49c7f1aa41b445855a942915b7346eeada348a7784d850625dc727ecaaec8fd0028cf1e8702ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h334d8c87045719ac529c60c226203314676626e4ee03c1e818ad0a7e12118b859c1d983da70a7c04b952c4ac3947e45c8958cb060575d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h62d01112148e049a629272bc7d6b903a485f0dd9b08541bfbb9344533cc32a7dff76e992cab6ce8a6298c87f6823c74e06b365f9e853d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1620ac550c2c140495af049837034d8b82885a74f78b4668ee3509074e29bdaf603ae7a16d516a4263057238033888806ffaa89f148c6ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1665a4f105b8b9aa1610c078e31f3f629efd40ef5ed69c9cbb584ec0c453ac3f6fbbdb44770107d892fc27b7bf853642cd8b48e527d6b5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hee9406d578336c7247edb6bc55afd363c2b86a6c982c15df6944e4b08f3c8699c1ac1a78d306638e166a415d0301cc9dc24a7d96bd2d46;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8441977608e1272fb845b9d6d0bf8b7382a382a8b1ec04e90bfed0fa869db918ab50cab3e465c750a1b7354c485112fe965b25f73d23ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc9b07714a83052e6b6b603364127d2a1b1f0ecb14cb39d2c44ad06b5d09300abcfc15ecca2daebf98ee8eb9c244167e1e1d40dc56adca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d896c8c13b6dd06cb895158282b89a05b66465e7b99d5a6906b018ab08849a6b98767ab44614d8488778a882e20765f6c4d3caafdbb95c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f0e7aff562c24986b12a5c1f64de6a617f0336bf499f124645a4adfcf77a04106a00137de00453d4c2a8ad0bab453302510e4c9d70521;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc972a3b67a8f983be4f13c9518bfa8ff9016ebce24afceb9e7f233e52e2dc69544c0e70826beda77e38cd7b49cd21af4ca474a52eaf232;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4088253a497771a3415a72092413a58410196edffe4928f5b376fde3ceeb1ede93099ceabb706593fd638c00eaa09b5299a0e081c8f788;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5de9431ad24ff913705c9095e15640c5114686d4810b367e6a94febdfbe70c9dfb686ff55e7c1f12530778c300b58437e3c862c789938;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17b37804ee2f0391986d5caabd97c2afa74b3c44eebb7be9fd6d8838bdd638fae5704eb14f275bf7fc755cae4f730016322bd90366f0619;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h52f712fb6db906772cb5d21c25068468eab3828be5b72fa772db1b25254eceb157bbfb0132a12abb0767206965dd70f19380566ecf6365;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14fa72304ce318ee387e979b25c857c2dcdcebaa82cfeccb878e4b39e118214fa25f12c8c82d2d2d76f7a1b8cc593214908240b91db8c2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a07579c11e615bdeff10cab91fff25b6408532649350717ab6e71e819c9000300eeb7e4c18785c2f82191b71f53798daff73d6b2971856;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e80cb178748a0a818f59e893f08a2bad74c39278889f31965081ccb4d12f63e1527cecb57ddb5c97ab6fddab2d7b68312197a6e3ec05e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h59fdc9972f84072a9be62ae2ed522f6e2d000b6b3ec1aec50b1377f025e06b71a39be04faddbb2f4041df1fa2bcfd41a3f06cdef0790f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa7ae01407f9d5bda68acec9820f3176354ffd5fcddb9a502f1277050836051055074714425b51328b7312ff6ee4b07e1f08aede85ee18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4a8f02491c1ee45c6decf8b6ed64e70b1bbd43e6ef88588d39ac5ef81c63dcaa492426ee1b9d762859adde951a8b21c76c941313f71149;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11350fc81cdd41b5383184bd6d0bd2016a79dfda3a397b1524fe60f57ad9cb5b3a369304414933779623ae127e5762482abaa9b2e3c7e3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c4b2e545b67863243370ed154d170ea2ca0222d23bda654978f4cafc1ba379ac1026990124aa70a8c45e0711f1c3d0dd0c77db6aaf6b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b38f4993fd10a33a01aefd51040972792f38e707e797ea25a6fa2617c34dff64da12342737f0dd69d61055329d811ec9be5caf4a811108;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8066bd1460782b67e6e382d892a287c3221bbaade8568f6a8f72f8082346437652d7a0eab2a84a10a1a08a2ec1a5a4815c72cd55f3c17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7ad3ae6781f0b24d6e49547036911b252d037c05ad3e4d9758ca254f2f6b337826c790bbc6d3c03fca88250723f50aee793dfcbdec01e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd8b7c68128327ecf1cdf7551f31b8def09425f4028cedddeb01f762d0e54e0282f092630f44956b621143bf202526438bc8e4b600abcd7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h381220b52d4a9b8fe12b72dca7c75d00a6feaf6629110d11512b13803248cf844159f8ef5b2ac3c7455c9c85fbbc6bb454a82d27fd6d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19b0540263c7c87208347af5c072ae0c870e2ece23919c6f7af42ed26d80055318e19ea566cad21163f2afe9ec2d2acf30e9be267661f64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f0f310b005415dba61a2df676f268486a4947522900b1eddc6a49263d15fe53d5a185c64edc2cde7cc3bb8f48826c572eea0090a53f535;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc413b0e634f0f998f3be9cb2638e45f4fb804a3a273af3b7fe1bf377670dd97b97bcc4c34be63037226b40ef3a669a0793f9cf6523ec8c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc9e10da04580d0061291b25bb69c4cab4d295df7c7ea248cef0c0e9db8298b0e76acf7d9c1a7ab3b1ba90b7fdf5e85b5cf45269d0df85;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14268dc5bcf62bd8f4b92ad41399956a4ca0bd5852372920482da860e249c923d4ce9e91fc220febc827f503a9af58c1bb7585480b6a267;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h956eb607c9c1fa6fb3c90213eab79d08d3b352ae13f4b17c94d21c6059e07687ca647a21cc2a9acc977ae05a6f3162d9fa6e7cdc33a653;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h884395577bce146250cf70171e04e4fb94ea92e5973d986beb0333b7d8c6fac5c83f385a2c9664d98da8df1f3e0c9b83e2b7245a8d813b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181d6919fdf9ce366c702d30d52513ad42d1ec0ba2ed664baa7a0a2b58857b0e35f4595a1d8527559e1294612812bfc521db95934d95da8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14075abff85aa3ab653f56ff79327d58763368bdf975af73197d0acad776ad9549303cb466f829502d8b8d47e143f9707f215c8bf2620e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1207eeb7538c9964c3c0a642cac6a2468ef9dfd6c878077f5e6127e5660a52af4601ade3f1bc719cbc08d4fb4cec14e7cab80a6e2fa82d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fd6358487a4ea62924b7b8ccf95b0500eccc1869c4560b7ca95649e9fde7859f8153fa01fa339523e0dd3c4046c1df16f9b5f8693ff7b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4180954fee42da6c4d2d61919e119ebb7f1faeea5a45b83035586a0971a69e736cf8300044f35f35894c4a1189f616cc6f70cce969075;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h56eeb884b49e3b067249e8ce5d4a362573e44e1cc94bf93d5dd1e819bc275ecae2d5bf1aa63c444d337386e4a08e4b2f88f8517b89aff6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1892c5da858485efdd007d38880cd164e3429977cc035ca9ebf754676c6e3133039c66f20268810ba76ae4aba87e07051d4f328b215df18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hafffb55b22017b49d682b1c54b9f35ab7f59e793875bfef62fbc85e308b2eba92653992250729c64cc3f5e743299f36f5987130cb800d5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hddcd02ead0f78282668bdc197d3a499b196a71d935e18bb4c0751274ef87c234a0b7e2bd152bfe63865b27494f1674a244b33506d40ea5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha1518a453ec5c5e1aca91f13fa58a32b8c2313f09832e9faca09f3ded139c7ced2a9756025565ec5747d90696226ad4629dc0f106be26f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c0efa54237d030f2c81706c2aa33c15f3a9667ad8f2a9bdcf7f9760e35a69aa114d2254ecc37384da6d700359e8f3e076cb2b8d707040;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc57492e73993954e27b22817d576edaab16e5afe18c9da243daa475ebbebea66a296227c67ab7013d63857fdf7a342414eefe6ae0ced41;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69be207d72547adbd4747349860eec9827b0723fe531ec5607fc3b6bf9d686f6bff80dab6a13f23361850e953196d160a574876bad3c98;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e71f8c9493f571517f669a103e6e7a26acaddcb0ee7f35b6aeaccc6d76cbfa0089a107e875e8a61a2bfa02c8604012aed85613afe0686f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181e770ff06d652d743ef3903ab3eac27a10cd3f10c126073f33d2aca087cb507f8e483e1a4ccc4d06956edc281ec1317ebdd95a8d554c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a740aafff5a1435d1b7ebc7543e16b583eee1a142f09abf0726cf9938bc01537ba200fa01f36084c26b9e87ec1bac0ec01c272e549f02;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb9af4e2f5405a6336c076040a768e001e380749d87b12a046e6d861ec2536c866825f70b13b750eaedec72b39bca51cc8a737fdc3a9235;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67d62bed5580ea0b8fb74bc01682bf7d64d8eb867d78d7b121808586432c4055b3f55e07cc1062fea788fc38c73e99183be2a75fb60b94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h29dde13fcca5241d21399c328a7df54f6bf879bef30359f16605ffc48ba64372fa691133c774d16941aeb519904ff677ca07876658bcfa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f3821d2bd863a9a62f343773f6d7d0999151df5e694252928384d84201da89df7c227726c0206c1b19f559d6b60d17876a3b7fd68e73c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf199a547863a1a93616ae09789e3576e1b1835fb9e74752213f87a0c5e731f95c99dc5e05311410b8d3c8b058b4d9eb604e0cecefee241;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aec557d6f28787668c9a598ae0fe6f70283335e89c419650b90786ae6417bd1c9251ed5439edac7995f707ccb74349411839b35c98c40e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194c6c27fe2a9d305402d0f15127b87d6e11b6dbb941bb75980ef6ee59674c0075ff1c2c5f90fd932f1c2f258ef1dc779a9712c25bed901;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b2a0f9a8efcb5c94f490b279a12267cae3b9834e0b7c1efa8b8544898548b5344b5f2af999ad1a3eb83837f999e7f5125adab5c4e3708;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h154379d342d092f717804af13e033bcaa30df7bc415ac69cb144750e5f9bae7898675f75aafbab1fe55c567a661668a70a8811d29c8dbbd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha23e9d5e266677df97d2b5803ca982a15e467f51a0f9aaba8330a5741b6c656174ad463490e8b57978af5a7ce30af15cfbfdc73e95f7f6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha3b68dd9d13a9e7d86ea8377bd5e44c3a60d40936ac69307f41282cd17853e2f724e8472c29ca916b1fe49104decc43e148d782f31fbc1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2cf606b876c8125d8de4eb49b304069fd77da4e9433b32e91c601440a0e148d31834e0666499fb079b374f353a890f53b446542c7ae63b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e7191c7c33f04191f5f39749d5a38f37750f76b5d844e45d459630d28dee4c6580260402bf5d833bc602080bb57cac075e4d6137f0d7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h22492f176d4bacf0cccca4c781fde820f0d82db82e557600338e128a20df1527b5f1c956122bfa8d4749e44877a21b19dfa7eab96aa26c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ef58639b83312cef399724d575551c6dbfbaae3025b1007d864de594e28f3f3a3a5cc8c8edbecdfeeb7f5bf52c9f34e828b22a0398d15;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd89cee1486695713064e2fa00009a8f4ed5523462c71ab0b31d4ba4a858ac85a09444df377b24d77773cb8430787f521e4acf56f83132f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13257d0cdb500657bf561d4c10a1961c30d429a5fe4d029fa081569f6918a86ecfc05ed57ec0ea96c6c78c325698581cd6178562e4a37f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12d7ebf937f17ed0062ca1589a40e5dfab57f8dfd69937bc83ead6d99c6d7e12d60410f6d85959b70f4c529e657941b5b8992626ce23f28;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13a0865c30610bdf396ebb1f3fc4c98b084f868d7af820ffcd5d86cddf26b3be7fae4450cbb0f5b3d493306ffec69e2feb95e595fd2d6d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h126167838a79bfb81e86c001277aaaeb0f2ec4a41f955aff128580311a6b2e148333b8efe99f476d2b22822b40556dd2f590f1996cc7424;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bbbb68e3914d1d1ede6ed3a09f25c11924d88b27472a3c4f6e4a50a6da31364d808e9465f5d35b0744a80a85154aea6c630f9194d97b0f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h65e7176b8c7e51f371927f43b9d5d2be77951dc0f668c4df232d17a448b086e61787a880b7d0b344a5b19c16a5f1b4266ef91fc30dd0ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he86f7669198ebddc71629ed4f039be011f5429b3c4e8f10edd02fc18707553ba85db92c17d49aa37ed64e43d09c0b6bb81aed2c6c27744;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h273dc9471c038c3173ea1016aee2ee7e1c53d058c78f88e1af53bcc06fdf22e8cd484716d7540dd50266650a97a54f64c620d66597f4c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a80854ae06161b7a686caa04ab07900aa077ebcd23816ad39de8ec0503d771f3a2be8e3da8ebf7c535deae13f6ce4e2a3ff06173b1dd0e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h74180d4668e4cc5e49719cf1a00b78f457d1eb12b8baab48a9dd66f9d3c926ac00c6c850385c3fadb61360da374863c0521acd56084ee9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfb7edc78a784ac6f5d94da36d1119584af26922af3bfd18ee92c64b8a2a863d002566b73b11eff333449c04fdee1c05c96a19b917b04a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h788725809b5202b4d69a1db86629663124a2983fe5399ad14728682f6d6dc7a384109b631836a4a914608c12d108fd06a67fbfd3e7d37f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e315e5f175d330b6f14e8948f28c1dae30d6f9cac673f955c738901b74c5f6135ecebaf717f72ed2031bb90ebe7395ea5e086c6831c0b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e2602b3cf812026c6ec859242b9be4acf1b003bd2335a0b2b796cad56cea19c0803e2158d4face0aeb288658c9669925e18dd5526df752;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b339a2ca589f801d8389d42f776d76a8007b8fed725e9764cd9c036aa53dcae79a987b2f54f62d203f6bf8a57fa3d234f8d56f31900ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf65d4c5ea6d8c5ede2f8bc592e03b028169a43a3aefe83d657a00e376497d9deddcb006c2f8d84936af792d29445331ff47e4b11b14925;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h183d3a9f2d24eaee89395159bad81f72f21eb1c502e8f4399f3bf2d5d3348641188289a115c2d8824f17b73cd56c77898a7f02d54ce3f3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ac494ad6a257078362698528c8869561834e47fec588c72b8d426f31113c67334a3cd853d80686c9df16c6bb19e2ea2e04dcff17e0c67;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ae52e97260b8647b7dd91ab7134ad9a6307a4887ce21d4bad7d9e977fd2cd92779234a3b3c28dcd2b7e072a23b760bf8aa61770cb0072;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e9506ed1ef19c5fea75b929da2d86fd87804c84a741510c274d2ca9ec37d0a582880a760e10e8fe2fe0ce06de9b122e6245c7bdb620195;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10b870c85d48a34bd598d6dc2ab03b030f4c17f90ea7aac98778443f825fa324aad1506952e5524c771f165399be9b3b04941a171079c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa455eccc0fe846948c3a6dd6c8c8a781bfb8cdc211c7e08895665791a50d5fccb3ad2a58680527c2bb9ec219da50f3372d42862c11dda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'habf408881084de930aecb64145315ee3ef631e07292b0f4310bbbdfecb3296894a77aa39384c49f61275da49199e4887ff03c3e1ab7103;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc3e7d160086622ea87866a11a2ecf2cd1ee0798cc27ddd2243b39c4eb1a3752fd1d69aa6fa0137235b6965611951e435d2534e179ebb06;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h190f5299ba9fb54eacefeca6fcbcead22526b1cd16abd53bfc51aa9e539d3b437eafcf80c22fae4acb4860ddf6882ced4fb3f0e2f6bec9c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc35dd8c297619c96789de186ff98df09c7cbd94b33d8b7bc2aa109e2ef4484ee5572a0880e8da7c89a8adde06383270f585a4312a6e24b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h96ddf75e9a45972c072c276593496531bf81b8c4af38d827890d947e17932bed70572c7dc6b6205bfd87ac0330d878332a43e180e5fbb3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he1ea31ed81d19d302153c1911318a569c4f38c842481ea691c66a4c5bd9429f940d3e2fe5cb7676fb209f7b8f73fd957d3321f5a4d407d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ef8ca44c39c27ccb34b71407defac55e8f2859d3f79def9c0a41ecd2c1c365d46c969d047cdd5afb7eabda379437ce51bed0e252609c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2aac4e4e03a595a43b0f1d90e7da571f047eb1f600196d6a25b5989ca44e90d09621ec356fcec0925504c00a98ff5ceda5cdfe2eb42c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h108fb4c14c0b260123b3525c464a3344512fe026e18eb625f66269fff6e34cefa09ca86db5d4716e01ea3a5fb9b0cc6562c1ac92d26f772;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f01624a95495d82ef0d727db5207f6daed93bf973e95746ad9c8ba3929a9ca0d70fd0fb3d14da834dcb08c81b7fc721173157af0ad4044;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5cbd3e15cab22ff0a531790b72b26a065fcb1e6faa76d15d405491f4932b52ee4902701bbcea20772e1a2cab69ce47ad9b0358ce51cb70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c012eb7fed7ca275d2d21130c86bbc283d6a91bb89d4148779fda67790384cfe93bc2a4694e9a59a628551c9d667df68702f2067b37d4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f16ea40ea67353a6e0c110f6e20bc36a83ae7f40c4e7904a26c8e6b4872ec55dc71ec0edab6573740fcfa4f2e07d3660ab5e3c7236c4a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc2d574e8d0ac91e06785c2fe53327875426abb9df85a1b3d0ae219f7e5d8e35782f044c60929b1514b5f88e7fd6b85fdc8e7aba5d16433;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h105389464083d293812ca21418c42f3e04faf671e5e2c428beafa6501c081e35a8ca7d049969efb53091247553f0eff529fe8ffb4762e95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b4aebce1a5e42998e2bd45cb9f3e9c96fbab6d4e94f03496ac4b7c294a488f01298b4355d6a76bd20715de115a86539bb05c3d7e4dd548;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19a427f05ccff10803218415fdc0a8ae639b76b3352e16cd7dce78e0747cadc6ddb3efe72aa31a55a47bedb72c15111d019dd154513b333;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130f4aa1606993fb5344a08e162f4fe6a8cbcddc584753eb40e9faf238fece1fb35665ca1ae724871071628f4119678a6f06ed6dbbd709a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb4e03e15c417893c2281e47b716bb4ac27c1c5b5bbd78ef79448384c7d0540df0b820d5ca9b2f97bdcf03e498dcc6e59a698efda6f5ded;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e4af328369526e4e28ccb2e7d883f19521cfcf506dc780124277508729700f69eaa4ba7a2f7c4efcaa8b66714a91a47d77887dbf1cbfdc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1585fd7a0ca16ad2577316c4000ebc2af7d3e6c0a0c440ff4d05f1ecfaeeb49a2025ed38d941b2f7174a34d956d7a44a256ca29348a51d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h30cf9e775b900c883eea1b1d4fd50c39945ab0f4fe3f41c9539370d46835f88ccd945535f0ef831d041625122d74684ab0c266ac1ed20e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1201f4f8ad1e268c0275968a8c4ee3ae60310cb0bbdc4d6a1d3a23eb93a76239f3df4aa6fca8e0607d7d52c25adc7da95bf2a76830258ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd57a582dd5714978cc30108d0d30056ec650e1e37f00b4c645ca6530c1129e44b6e8c44e89f41672614fdd26c77ca87202bc134fe532a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd9bf01d473eb42716d6dc8bb857bbc9174a42d542de3eba9d8e055461cfa4b8643e9573be516b729c4021a2dc76fc54098c580ad63f498;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199de0049243be30536846eac364edb454c58c195d7aca42e623a13e55abef5b81734a630bf62a08c4724648609b75dbf809d2a4e577669;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4840db6e4f35378bef863ca97ac36b8f2b04ea650018c2052a64cc66ccd91439c409099dd249dbfc466304df2c7d1e5555d9ebae2536e3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151eb91587375c51f3aafbc88680f905914a2845e4cd61c06a8860a771aec34a2b3286fc6666343f5e6a86da2ad0b2e681a50a4e6d72a38;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17dd99fc36a24cc51753072c79603d432597dcc76255bd6bb9b6e5e630d604f04ec121d1ad22e00afad35d3afe2b889979c4aabd6298126;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9b2a8ab18f8b38c7daf8b0d25f9376085254aedc72b4c767acedf646a278dc31e5938db4fc0bd8efc12ed006b082bab735bf0142dbcd6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12cec4dc7d7ca6709c54643fcfda4a421981ed8d81d2144a729176997e77bf0dce006804d428c8d78da7a7eb3900783c67b18460a425ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h700ec226ed6c650abf6b5ac4d4a61d80988c8cff3b6db4f481715bf2663bb3d66927f43186d827f1fbf7c10c122a0d4aac15686b86fd61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9c0703b0c7e6484d2598fbfe66cb719947eb870dfb17a2d765e3cd2a188ee69fded76cba34a34a58ebd8d5d44e9564d44bb8cc90716d91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2401ae52e6e72003449193dbeeb3ee9c7039e2a58f1fc564667cc4fcc1ef8e585f0253e41a5cec0f592943a51c147d37d0236b1d49171a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb9c6d7fc289e7c8c2a16ab2b95e8323d583eb84a7cd20410396db32ebbbaf5d8b5c67f55b7f5ce30e464a1800bffba359143898e0895c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea6fa69269dac401332b90f7725ffa266456c7fbc8b1c1f1896906452c8af1c1f30728fa9f0a7149733b090c8bbfc03955a41eed7507d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12884f59ae20b7a83474357ddab2b516e79619e406df259c13119a080aa5becec7879a3f8930ce3076d3f76d3a40557593b0373a3152d0e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd6444152176adfdd746560553e06c314d4c07616cf36d7c13cbf560cd6505307a36eafc840f7d1a1dd118dea3063cb6953648fb9fe99d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f26cd0a6750b7d3ed97175b55cf0a1a1ef326ee19b38bead7e9dc1c758bf3b829fb95cdd82236fcd457f58d917e46020cfd355db9b27b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16a262f4f6212787693f79e8af6f9048900e18df0669aa05f7e3483aff1ee714a0d8d0c9d233fdb4efe29bbcf021737e386a94ce2a83c79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1096c2ed2a87f390a517a4a0800f12b01f079ad796ec933847915a7057d7bb52710a032001e226cf6dc89f4a660a08cbc98b8c9ab96a482;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7ae316ab7f3107bc9c090e7f93c0c506e43c87e29e891d6df65e438279d6fccdff27962131dec5ed0808e4f6a72ba13f40051915437bd1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9ca0d284307646a480abd240c0cf434c05c855b6bc4cd8cfbb149f43c65c69dcfe2d3eee9b784321cc0bbf1e74126723ff56ac79654a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110d3d30b1530095edf9cd5015bd303da1750a4f273255041f36b52420fe94676a39f7f29eb5e3191e27599c1fa0455e72f82e12c87bdfd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5bc0116b56d3ba27be42ce6dbf6d2785f6c8204560e6e50df9a5a31700d26b66cd3ca488cc459e955899b701e97292f55ef1731ea740e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19cc2857655ebbf3f1b21221f847b5436860d46b18bc3e4cbd42b86eb1de07aa7156c5a11f8427dd63196f6450388024aa9fe2665290af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1609d1de055802f964f5ef5f662b197135bb75d42e71a2e729784fd147c72eb8653cb52b1709e83fd24cfc7965b542feb021c5db56a17db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d3c77c321a10da93c3f0ed83cd465cd4e1aef15ec8b55a7645ecd6ddcfba3b1cbe384a7b71362d81836ac7f515ac843672be00b3c12c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h360c14718baf5e2e752119dbd3bacfa5d632d33b2202bb68622b2cc4179ef1034c761009d07cc62ec8a81985a1f99b00f4f50b6f7a491a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11325a5c1f3720446402c98aa87c3d1c8e83a00cfe17fd896c33c3065077568d56f426a2361d113a83efecc4f76d1aeead0d6c2e51a135f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha66e125f7447c4688ec5546d7bc21225936ffa05e9ddd282dac36894cfe124cf2a5a68dbbfd5c4a9273ee81678c793cb469dbfbddefcb0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h223b15d9089021305a3b30e3d3170aaa64d96580209d2c9e046f6994b88df950f81cd9522474384d53e2147176381f49df2f8b3d820448;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f7971d34cebf98d8abfca61fd7bafefa0fec04fb56be5923be0e055980e36ffd78d375d3392ce3ffa518caf0b05889579ab02a825aa97;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e3e80cc84e80d916c3b3bc0ee502bd41b4c2d87214d24b39ee4d8683546e54f09adf4b92c820d1560dea3d9f4ca2d72b47e0c45ba3e8a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0dd4014fd26e075497f3d4bd1c1c5ac9ca6262895dbd30b37900f9812aee39cfafa89812b8f817963db511e91eb62d8be9ee124a92070;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1461f76c13614a7ccd0bf97055426468be1dea56af9df712610d158e6dd1adaa6fa9c39ec21cbdf32729d0c9822bd246d549c24fcd12eab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1837e7513c353ecfa73b3d6c041c34ba776488871de7b1a0b9ccc86508761fcfe0ae98b439da26cde58e4df798ca575a78214732e68a266;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cbd955aae77f74d250a7db26e1a886c14818f296c341fca0e31be736e9d3c0eafbee78563849e180c9308217b458f54a613c33b924004b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h113304f5bc184fe9242a98078e4d78645eb4b64f1b7b1960dd4837a4885da7f6c0d538e5cad8b84e375180759a756aa2786b2d3a1c7193c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1482c8581212c97a55579c7612d1395f85a6901500312c74edf2f26641cd4a994aeed8c2c4fb8960025a0918870a7d9fb0511c28741289d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b602eed35aecf662a8df74e551eaf0cb6dc19a16dfd123a49e877dc06d576b5abcc3d1a678bdb62587774adc0ee828c453350b09ab5ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cc4ecc14bfe8d6d1565febea5ec578bc1b0c2be3c43439cc4fbc001f222c7f80ad38a4db3ed9c3423310cf25aef1c87794b3689d811c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110218afc9b3c91cad2ddb8d9fd8239a9fc2cf04bffb28df2d5cb2c56fe2cb475c7105707f442ebe6a5ee2d84dd451c4b1fee40f091df5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4a500ba502cefefadc81da8fa1cf97f34af94e55bd904451b17abf5615bbcfb99303ffcd8c9e85ea398fb7436f458f0d1a1d03eb670605;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcfc62004c4566d8774aa76e0a552f74ade4733f9d87413882dbfddbeac60274cbe12405f810ac2c456a8b4bdc1c66d7747e58fbd046da4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb6c7ea26d20f4f36f2eda1a10cf6b22a3b91baf9ef1dbb2607238ecd923dac7bec587407f91156552f16439efcb227104fd1cd6480719;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h874552db8ca10cdaaa6ad508b52f46337f94254c227387b5165ac8dbac4d8011e90382980fd6f67d5d8eb58654ab2964da1c4075b290;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he83d3a31b767a1e1526e5e65498dce981ae5b2352d563d4864da936cdec8c81e5508cbcab951adeff617e538a76e081134a3a12204fbc3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h150adb13b941d73bc044c8fd0a1a03209208ceedcdf4ca34454f9500f9d0a7f25700126912f9f680813ca0540c995242e71cb88bfdd8b9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18214d8828508de63ad627df3e79c2c8fd240f70bb78ca89322ae25e45e784940eca8e69fc8aa82de9a32d09bb05e11a01982a37fc69fa4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0307834d1d5112e635da0df67a12d88223f7195aa9257eeed5325c74e94a1e74435eaf77b62653ef12874417f9c34c1db29ff3f6e292e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h93a850a402b3f9ff32929ca994b757beca7033127d71b31472d0e44bd75ff784a642419cc719f85b58db498c66691b4696769074a6af21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1329149cb89fe58e99aaae15ad76ec844ebffac1566a0c4dc77c98477edaebe8e82ff87ceb822083744be5341c39c212426f0455130a66e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c3c406fb15112b0d652d5866e3e33a8a910d48aa2fd77752a4d7cabfb1e33d90ed290d2eead2df648520388e503f8bfbd95ab013000cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h175913cb4110a6e41ef2a3541742b4962ff933c6bf195829d99fd3d61273bce2f8470002d7f6d5839c103cddf5ae4bd45bc1bef5a015daa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9745c7a009979c5926d4c559e1169a303e457928a3f8bbe4030667086813657f4dceb69abad1ebad4e764827d0a5d0955d835af885430;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f9a07f8b4b2a80288cf269a131d471a1dd9ed2bbce740f28eee4c3c19803102c11af98a6b845ee105c3b2f954738b9fdf1c993d3360a27;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f7f00ef28a911f10172dfd1d4d6dd28596ef1e5af47b205da2b92fefccedf8e60c1ae939731e95f0d488366a0308ba1c64e9c0055fcae5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fca5edb8e782f48247e95d2b69209b9792fcf681a0cf87e3885c1a018ebd0850af393c37be6ef522d4d9b30eec245300395b2f9728e2da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a4f4100fa19ce24ab4622f3855cc7331793b6ea3a04d4a3442644aecbbf5fe03aa2d463602c26736954c6ef16098f3647b78085c683e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58e4c796e416e0aec0e9053d08f41cb389c98e7a5c9237ec537dbc149f39fa5f4cd976bb3326c4932446fc4725a1a0d43b3084264d16b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb3abb76f273abab7f887e6a43bedae8d6da7ac19516a7156e8709ae7703baf621574a14e93450d66699627c38c26db44f1a4f5e8269a4f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b65843345661224de14a9a7f1de3355a89d5403f9866b17db03bc22c23408c293de508fe9aaf9d5eb66071c4846d8769619d37ed92de3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he9c2e9eec3ac7599ef8e2d1cedf19865bef03e402a47f3d167682c4bb59fe5a8ffb99533de69d5dbd06738d1fcff513e0ebbceeff678c0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd499130f1dbfa8f3c0bbfa8882523c257dd052c9b4d1bfd621d684a3b9ca1a5a16ed9b86fd9c11af15c3c2f8b871c37ec0cde5acc33e3e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1966f834460a5fe5381403a11f79fe811d7e8748ca30d378f45b123577f2ddb42436e86c9b99b81d7d0b414a6fed77439574c5df6209000;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fae35fa7c6b7c81c34f3ca2c4f7f94fed216123aa547df6fe4c9639c541b20cbc816cf6cfc64bd18d5cd624d85f204a7bf3ae6700144f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5b2c87c393acaefb34e7b9834381b049e642488d877f064545ad8cf9f2cc58f4d241667cd04d189b4776748bf54a33ab1fd4b0670c4060;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dacd9917731901b83e30c2e39bcc3b2d2195211bfb76874ef66e3fbd21de3fac350a9120682039eeaa0677f2997ee85700dacef6601ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1794a5bc6e2e9481749192cda679c511abe11a13b84be8cd166a09006076a9ed61769414f49d59be20cde0796da14f219dd19e034632408;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h47248fc6e20dcef4dbb77c47f8d6b4abf14ac4e972199f18174d4d4286a18339dab2421747888259a2a3df260070fa2101f0b25e7b8ca3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ef080c09456551576bf82e0029db81d67cbbee840f02c5192f1117d213fadb3da0e82aaf36045a650262f3031979a92da984ca9d6f3a3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1590054c64a35b134d11cf08bad87227b6b89f980eb8fd14677d47cbde71015dd2fed798945fe10351e22bf49b467c0bf174aa12d6f5d4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h36ee5595be95d6847d4de90fd2c3f76558de23be4f5f1e3606e92b345c645bc2d698c30a004ff38518f026bd21ccc7a528b34c98e0bad4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194a2fc2ebd33c03085f1502084fe17c3b99db43c7b4a4be097928ccdad0c0c94ee5f855fff8216fe13455c9ff901d452a58e19867db069;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c4334c005cb3c0ea936dce00962e6e650c813baf135b62de221ce85019cc236eb2f2da9d9706d2063845bb0d89055d7e1b0a11e85798d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54a68fd7f787050974dae3437423718698030c6a985d4183cb5c90f0cf391f0d363d8486350fa59c2ebc2abe93470e30df7d687274cdc1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h52020b776f857fa25324d131c3a3eef4ac3ce78a7e0244e36277607ef534f09c46aadd492132484a93d73fe2f8bda64be77581d6d0874f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1116e13988b109e033015449f3063329cdee8dc325c7d713fbc832fda13e5d2c1bacb009e64998f5dfc51f752fc55c5e2378d1d37b995cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6b9fa7e0a5a88b37926e03fd43070ebd4befdd3c73f49e5d35ffdc90b140c8827c666c3ccdcb3fbff2a0cf4dee6cea51defbb31016bb92;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h634762ede9f3a6457fcffb22e4c7f88f0c130aff9e920f1e6d7788f3b05b8060d93c9fe717e36ce0d9d4f396e0d84a1e56f8c8fcaef5da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h489350739dc1ee764af7e47b164e6e993cb027859a91790b078e12d73dbdb5a38431334db9a4fa781ed9b8d65d20a063f1fe77a300d7bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d72c459b59cf459cdd2be2c932b49432d06bca15ae19eb5b80d751ee5acc5eea960f316878f58df92dafd1f0e42af6d9f76dda4e9685d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h900d93392542f1c91424ef69c3af01adfa1b6fea4c335699df3b45ea8beda456370176e7694e45fdc955caa65e8d0063b3476224cc987f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h47aded6b38e3c997062a98a1a16d564695142625feda6f6f12ef0fab24fb7cd64962935c1521644df1debfe7ecb4e7ce53e12b1fa0a474;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11cb1e94fe4722332db586c4ff4a28a1d3c4fbc275df10babbba23c0b4ff82fe7b11ec90ce39753db2c80ba86480d91fa621e05826e8723;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ddb1378e0ed121c0fe329f9a2df4b185db4b642f4b1c244519f0cf8c491d4a55009d493836867cc01e164e1b49d44728373f653597f589;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcb86f014d0366b00d76c84ec9a3ed03f04a01112f5ac04aada3fee2e38cf7ab1363f4c7f43a57cbe94b1506deb363bd60986e4bd8f4975;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b04b343ad616683e632fda911aa80cfef7f0b8545b81be0a38cb74e935893d66e21e400ec6e9114a838a72dc6a1e727bf830e2c9abdb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12853118540e3044f067797c4841bc190e4236377d0ecb9680b6296f4f7e7fc931eb32f3c37aeaeda40f33db695235e378f280c1bbac610;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8a74e74fed507d43ba7576f37d0bf32b0cc32daf5883e6cfe7e108e982a9dcb658ab6637613b94963edbea7d5889693b22f2ac0b2a4a2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6fa343d8d47b3faa990be2765b3db024c6d2fbc88cb3682cbef14e8d66f0324b7ec8885687b7d36e1506ffcaf9dbd7d4e5e8d9f974dec2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b3c0c5c513b5374e00d88dd38e5c56829cfb5e860ed9451c029ef4fc6edca22d8c94c73d5b261d6f05f689fb8f34435a1cb1dc026c3295;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19ffdd6a8d401e587766aafb645efb0bdc8a29245c42f9454f8fe10f5eb59940f4474b3c25387047ea091df118db4810c9496a45399d5d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c58a4b675ef96ca36a76c6bef47898facf926f7e930aba028be984380e3a90f31f75943da2a13d094576a36074ffa887a467876eabb99;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15c158048b21d23973c2fd3186af53ed73f6cc1383bbf51cb54c73d57929588a229dd07fcf58de98fc4f9d39c5fe7e8214ca8a34745fc3a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h145e20a3855f831e48592e7d4d54ee5c94241e5e50ec52a64d05dc55bb9cad9fd83098715429bbb1cb7d3717b8e417bfccf5cc718b3ca31;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12c16cdaa6685f7d2d879b44da7716d4b582a26e35ebab440c3aec2416e18252b8882a3c76dfc97c83abd2339a9e785eb07b9e60aca1084;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e4de3cbd111ea0d989d19df771b3cf1c3d44496a370f37d3ae640524316e7ad9c25932c6e3f7ae42342ae73a18b09edb46faa4044e838;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9078c8b9262deb4e1b320f0e60f5e1c56c71ee4843e4edec025581f8105a19f7ee14324db1ef52ce26a9dad17e31e450811fae9da167b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he3772aa202a9ee38155c6b545fe66b63774ab3f406c3a067fde232176c7fdf56d0f5aaead0a8a7cf66e1a1593d86111208772b35344cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e8727bf3aa075ada9b59c81b57b03b807a15e57657b24237ced0cc4c074cd8ce0404223dde3947b99e23b20069e4ea229f7d6f42ef499;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81fc6908158165d136f46d56045f41a198cc7251d20fc2fd6b06772007888516e433b81a401fa50140dd54458764767b130c4814b88ff3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5409a5805995eb6d49dcf8b654869e686d0e3f78ea6e94b6ea10bc8aaa84ec8660098ddee60671c1cc8a0e149071d1b7b8588e6a4753b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h146cb0602fe039e1fbb06ca754f990d309684da16102b4cfdefdced42fb7d00bfe51f835f41ad3c082faec25355a7ec51b6a06fd5fb0455;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c4e75d4bd17f43592060a71cb6e6a474b39bcda61483127cb26097a6bb0001efadb473190bbfee4163d9b454a5f2ae6c53a1763296caf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf332438423d8449905147c6056a9a6cabdcf89de538a187c8c9609f3e53839fdb34b6da36a7f6dac5c527e248107bbb85d551776f2e06c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1abb7309813b4ca2dbecc0950f657f49543a6b2ec42ff4b76af4ef8f1b1c3f45dae72d64dce23a420839b913fb7af8e894a63a209c4ac21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f6d0715611e49d8d13ffc8410268a430663271a156d773f5dcf395a97799852401e987eeabded96153d93452fa6af0366f71767657960;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha27cfdf21b17fb22621d9bb4615e36f816f6c496f9c3d46b0e3acdb9deec44621635ae02592a4196f9c5fbadf0d6b51cec35d3e18c6630;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ecf2ed72fef99fec1fcf6a07f81f9d9180b7559a9bf31bbb3acc22c3bd5f65ccb59bebb8ee9748cbd0b7fba1075b0c49e91e59b59894f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h567f54d2b5dfb687c83777fb742d2365e665c7fc739ed2389520301c1b3cd17fc34503ceb850c71ce8d432d8b693d4e75996f1d081fdaa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd60b36a00c709e1c7f3db6c2b18ef29ff794d05b89a0d0dd5a98e87ebfcb6cf3dfcd789edc1c6b8dda4c36dc925ab8c06249d8a035067f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb33ffc746a1994a7e63bf7d68c47f8afd1cbabd88600f406eef40575dbfb84ad5a6bfd49792314cb09c6a149eb23fbc8696966c5407a95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd012945af117c7c5f75edaf7194c311ae7528a0f9277f01f6121f84e8552ec234ff5a36d11cd3890c8156180d576443302b0f9497723f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d8ed5b961839504332ebcd09ad07dbc23d78e92ac498c6667fd911f8df57b8b2586e5339dfbc570fb33faced4afea442c879f62028938b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d219f119cd04eb3b0880df5f28a9cf76199337435956594a1c1db7b8ded2e168baa5a880b7ea9428ac0025bb20c12887409204e3081a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b455864cdc85a5216eda46e2840d128da32374b7a219efe7f3ef551cd12f9111b873c9318878295a4d71f55228df435499dff0eb4eddc4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78c997edd17e17b85605c6c9dd150d861fba090ef96d2c5e219d99109c6f106a92342b4bb34a1175440c93f78314c346aecb6b98f5255f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he713e3f15589b28c73c78d471d80c6eac8f8683b5854345f06637c1e37618ee539bf02d414f29293eae46229f105c66719b05f6f4c91f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h418270b98be4a435c613778ab27642bd12212b8e8173d36b8e2198b99ffd45485c9c5ef07a97ff896e07826dfb5a27f53a958d9981e3f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc7ba1d5fe71c771920eb588168d45ac1d98f6898bb1827064dc7ec64387bdb21ae6095a2aaea3465778b29c636c5ccc79c4a026957adf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha07e1e1fac241145ea27d01f65b3af70f1d8a57f265ea1d1626cec2de0c45fe0d6149d32aafc30613a9f778db634b986719a06706f63b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5acfc8e63690298737990f5cfd985fe9474678d877b5025259c134358cea96accd4229b72fb4b677f80a60aa0ae1d3fc780b5fb892769f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b176e91b8f25017501c69726767dd7d18d4b78c6c5fc0cfede49426435dc6a3a1c488e3ab1eab33a2ff37dd4e32494529a3a0d8a8547e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfd59048e49547a7348d5c0145f7e887d1c149d5f9e8fb89e3b25be392e0e8a5047c027df68a9c04cede23851ad80f8e4db32a77111c174;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8d6f7cd7e38b376b133ed54f54bf7ded34406bccb5d272a3678617e681133ac7a1f9f274be36fc7e49b9141e8327a7b6626e839faa8d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157069a73e3d8d2fa7c1da12a23338844f6ae4a14a0444180a18c1463d35c9cbe95807a145edcc7e1650cef3660879e7b8ca08cff28952d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d4e48ed2d00a533a77f8c28feaba77aa15dff1706d77a1f0d4c294621a754f3c72df294d4bf1cab1589c9b9c5f83e78cc7755a3ca5bb8e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc1691bc328075ae935c763afd02647534d0e618455abbc7cbdf649fa900c592d74b77de22f0116366afd684842e179d0cc93407f62fb4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151ff53740cfb99106870c2c78c7e9c0d6b3b8d4decff61d1081ea00753d4d11774e48e8faa3b4aa2d99393876fa53e3e139269ca750fb5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1adab7707c13a6ba8bbe78dac5b20d7578e53040161bada67f27ba672b695013bf24f852a063a9735eca1b77f9c54fc0444838c17b7810d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d351769085a5d4371c93b49f22e5d2034eeaef64ee809f2cbce6f0e1ed535c83a417ff39e5af2ca7326e91695207ce1e946b826b87d1d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cbf3da86442ed798f5ff8aef2a4095a0692599a8e07487a9fe6196bf98cfb6cac3168eb306f6f5824533423622f45bd8b178b88d81be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5f0e2d849ecf9626469597a0f77164f54622eb1238b51a04e147ebe55a49188589498c38dbfbb42ee033b3ac7a7ee0ceecda8fbc7778f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h157ee86124f1d35999dc8c0e8d4c1d2c3246303778817ded808f9514d037b0983c53a8d5b6be71157dd743b792514ddf2c772b6fdb5a00b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcfd275f92d2ac0e8c008855dfb2e5b94f551aafd2f3d033767941b77cdf790aad7531a554e21296334c6f1e2bf2635bfe15e73212225d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1711bf4ac150c9c02d772205833928f78224501cac8972e4037188aa3fbb38e9d8d0051ee4a22e2221492cbfe9f903530b650f4e9835e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c446872da3dce16a1531fedea164774d991f5ac2c01ebf3a2cc21738e79b81c75470a9535629fd1185866b89cc9b89ea54cbf29458d53;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h171800d6e3ea8a9e98142c6b537c19bddd031faf632deeffd130e20d961de0525151908b8db931f9ae4aa55e47e201ff3755e7e43368186;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3dcbd04e186d2187c64858c9ee0b1c701eb8574e202f226a329ca5c52c56e01c2cd24c27c1a6ae6fcb2fcf79d035cf07c9b29492039781;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1566a43031a455c2c9e5049eea6bd4e8b733487ca81cf2b6bc1f3f3c3e8c34c07bc88afea27f5233f062c285ada51227471d4768014a7e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h132d77def36c68a5d2ce78b51e20b417b2290361d6496fd154086f96d14a35a2311c9cf145efa7a1b134b3a88c27093802eb7ba31f410fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h659f781ca317c6315bcde3578f2beb26fb6e360487c29bbf78ff4377bf5a0eb498b0fcfa4a4ce6701ca7d24be5418afa2b5417b314933b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13a927e1fab863883a55ab0e8527db323304d2606763c3d9bf2aef0a25adb480ca7a4ec1d025100db17ac3ee55febedb77595a2f5853bd3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5dc1b3bb93247202d08dd1acbfe392913c3b9338ce95dec11ea91a3bdb2e10fb0fcc7756048cdc1cb0b8b69f8d20ce1eccf31cf0460b5d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a7ad39d8d5860a3fcd5ea0a87a19b7d6ab42cc978d0911f86a16cde7933c5a6e023c6f6beed49b0a48f01349ec80d295359356d8eb5f4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f45261acd6dd79417a80392395572507e4b1663fef3bc76edcf9692aa51563fd61d0a5666d21a4523d0cd9fd7160393a67f29fa3dabf8d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c1df1d3ab29cf77c720920f09953761bedf5a71ac242f8c6f085c6257afce621b14ccad46f962b0ed8026383e3ed0edbde738df46c3552;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc4f57d6c39dce7f03e5cd9774654fc9955770b2a95086bffa6f5496131104050fbe2d358bbebdbf6e876dab169690f1b1c94007801add;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8eca1589efbb45a3c7c6854addedad89875d870e46070bf1665f905a164f26112352268d3dab13d28ac69fc7035f3fcd6c2cb06eb9af2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4fdaae2754fc088fe8a7e8923a6e9ef762a8b135c3179c18220e6a453043e8aeb2deb70222f17802a88039f5e0616bc4ac23c7375e6a0e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de5854526566594bc2d535454bda0a5889fbe537bcdde524e50b28e60d5168d3524e9225302cc752480cce3d5a04b569c2d8977c75f3fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h151e323d26897ab9f431b14ed93537350555cde8bc091749badb44ab1a7c1e5f658f4ce5982bad8d1dd1f39a998df52b80018c9ff67450;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a244ac82f1887d89bd19cb0fa89e43b3d4af5d692262836b2e12e974dfe568bdf66f5788d903d5d6930e687ae72604aff2b98925ce88f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12c6f51e5816a24957eab4306870a334e39cbbb9ef46e5868cb681d91e469237e81821eb22f7f4f84ed39e10cea0e16084b8eb61e7e1315;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf4453808099e07f9901a287c6eecca5e50184960cc5941a3cdf2b94bd5f38f37860c7f431a2a8613383e04a89b01a3a664a45f63dd15be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h112c8542a2229886c190da57be6207ce4580b8ebe22e8a92fe3f4c4920336401a7f66b11086ca1c3230d871eb9d8604ec1ca9da33369bf8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc69eeca976b04a52acae5007a0eabba9f2a402bd64bf7f30cf8d235683a33881ba03060ee4ca7ed6d61224e53f3481157ab609f9ced8e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d625558b77efec2459347a8b70bc90e56879247f93eac3a65fa8e226c4ccba6e137233951b0deaabff6e5a7e415c25394bd4a146f5c641;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1488630e4f85fe2932932ed8be228007b15861b51ef5c7abeee4df7c089d93bcc15a55c7e3aae906010916e9deef03d892f270d067e73eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h193f517a3c755db91b61b861ace2056f68bade86b31eed275936ebf33ccde781b6af75da0ee0c2746b5b7ae46e86ec507f4133d0d3ca0c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he504fa6a904881a009c9134f9c8463745eb46249eb9d51c492799d60237395da92a5cf6499aecde4f072a5df4aa4d45ad64fd58d73ef8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161e35be55f64478e59ad4b92029f382900b70c0b13298061fa0e5449223c6016c17b1859ef0ac630459526a68b85da5196d6055a88f196;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31eaba2927bd1aa14bed5320ea1c5fa2180c49d5ed70170fdb9b83a9a8c91247f13063869dade74deadd2271663dd2cf69dcb30f3ba3c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14e83aecffed1ae252cfaf04c393821d43ecf1799ef69cbbf100b2fb6af064a55498169dc5722d9cb3b7accb194fef86c06157152586a11;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d73933408a9c29cdfab45d6e9d3f91f56b4aaa81eb1f85d7572835326846d825ce2bac46b48ad328a4dfc5a3683251a1040ab0ca47860;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc0e7e684dca659ee00a24f6462f2504201c015b154eae6228cab52a6e1b1b430a6a04e2868fe6b0dd5d0ceadecdcb63afaa8c306447df5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd390a9d48b2161750c5c04cd89a8473d85ac29e065068d4eabc08faab4e799c9d828a546fb16f56c736149c01828815a646593f1452614;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d553bdb18794cd6ca0225fddae6131ffff44ed2bfd8879d16c53ef94dd8cd3587f622727d342a6b21cca79273c9bfea5268b76514cd1ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6617dcdf07957216c0bcc28e709c334a3f2eefc320c3d6d0efa75ae7ee9aeedc96ef0018269e66e286fc40955e1ca2b056c6a5493b7195;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha06050cd9124b40cbbf0e831b2af642987adca86d7387e6d3af4f750e3e148861918a0702cdf1b30fcb7574a702665560c5824b59984ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b44f679e25251b460f97cc58f5d0a3b2e0fc90e69c12f1e58979510f94757abeb6215f50794be5dd5bb65a42fd2f5b089954df602398c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11536e2ac59bb67d6b251bbb7264d32a317fce6f98c441688cb959f54f4a2565c7c9786e0c3a8bdc3838b668d2c9a4adf398db340d20d1d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17bc53674a99dc4994380ea1505ba482cba24462edf5c01a84348f45a0bed1ccae0da8c2e4b38bd97e581383de47b30aa9ddb95747196f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c68bffdeb5f1807887a193763c52b46f426eb627a5a93a388a08a3998dd1e03a9c9e461a2b9f2ca2ae483ef3cbc0856da94938fdb3026;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f4f82ac708314f661c8988749df0e2a78c780b4330361d70b0139a4f2dd3568086bccccf9049f3cb0156839e28455ea63c617639426ee5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10350c56db402f2daf8e9a85798b7040ad33bd1b5f208e42db54ac3ada5c5a457f66b50d91d77d1cc57fedd2741f1ad39ade779a82cf531;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129da72ac5af8a95e5a874c9a4a087bbcfc87ce40ff9fe81a0350b1bbd1330421e0aa6f933afc6b269e55abed9043b39c8ef5d180b840bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1503226986d6062cb9b87bc03a8e1d0ce20c007ff84ee9fd57417157c6fe590bf74254472c6f333ddc1547b4d2b89a6e23d9ff49ef9cade;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1259ec5288bcb9e19bbe808491d6dc05532274715daa929d39f78c20881cbb6d6db3dab05055c2aae553c8066e200068a9b1db0a5f7c5a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h972f77232fd01d0c354e20ed9b2d599b12a671b7536cfb54ac5372174c2f997e8e90e6060dcb99ea5e472aa277f00197fb7ea19d0a47e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ad4581a100e1cf01400539da433adabced99ca5c4872066e1ef7e682abbf6c2a1fcf38d142cecc02478c9e3b0f3501c18ad12f5e0a1e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd2fbd9e08deb728c00d2fe7e3cc9f0cd8438c1b119506327ab232a67d5561f4c6735775dc3ecf1c995edf2d6cf551108aedad8e73cbc6a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6134f61ac35107a3e5314334199a633765a7a85104f0b2985553c7e81f30267b7fdf2d65b763f280bc57586d366e951f0e033271c56763;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1883e9748db110c38e9e4da569a0919eb81f8ad4f9b0a6bf73c981e24e99c53f247702f3261cc9493e3068c9e6d5ab7335573652d307877;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5ae43dc88ea514ab709b21ad2a57aca77d489f1fdd05bea6af0cb55b6bb98af0b6e47b32fd4a2c544858e4198fb4a0c91ef4b375d90636;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63e445840b63435c69b52bfd906340a11e9a5f3b11072d07fc4c8e1c80f34958a9d9d06995137def33f7f77367ba6dfd066c0dac62cd1d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h122927746c9921c0ec97cb986eccb71831a45921a3361e73ad24d2ec2f55b46fcd28c2b5f85fd243493f181503376e094ec7a6e3cfd3a55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfb7905d69fcaa0f72f00960b3c6428f1e46a7be504ad3d8fa443d0b59d92f9fdcc86ce12c32d78905042cd895bfc33985fe3fe91dc4ee3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h111cb18c3a173e783d9d8bc95c9ccf88d627d8f5a54b079835f82de94bd6b5ec12d2ea401ec279225622af15326be33299c3327424e4ae6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc20547c5db2eb38de1304141c114b005c36ccd37be3e164e50ed9259e9c12d97e34cc2e8e3d31b03d5d4747524d0138dccad3f47f3afd8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7bf6b9fc7736bc88ebaba5ea18b715b9f961b0b9638ce0183d166bc9277109adbc91d0d35ae2713ae374e66a95db77080a5d610ae5c5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13483370213b1f64c943e6a322b8e5e0356be5c71d2a91f1e6d36a865ae10be2731c928d02ef757fa37c9e15fabe0bf1a2b6fecf7ee351a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2a5f5cc8370d6eed3b68ac3336f2304c1b9476cb1e2dc289bbc43ade5031df09c19ed726cf1756d7b62acc2fbda975abd408879a8e349;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1866e085fb24961137687b9a8038dbd0c369e09f0cf98869bb540c97054834f31cf24dab5f903998fa58641f3f989d828b08e603bc3a711;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf61861c330b2d76e310ca35f0b736d6a51f301db20b9a8b0d63d04ef4d3c0d554ff2a851c7c717f28a93026a715692eb28a5e061450ece;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h83e34272e8ce78b66c50b03579c04e21e3355b300b5355407801bd57df8f9c9b4f0a9bf2bdf3b280a3a6bde961617a89a89dde5ed9652e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19fcf7bba521eee4796727311b2a9bb67e933d6ff7ce6889a0d5ac93f896873c22b201e05d633b0afec834b8e620df2db40468cee86423b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f297cebee85b56c369e06ea90a0d4623a0e33e37ea5b3d6e0862be2c680de358580816300f27b1a01421d1ff832afd0ca3c29b264a3b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17728fbab6a4690efc7c8abf4126cbd6f3e180a0d08327f810073d86e2c5eacc641a6414798f3b53bc70b6b99cab72b94f977ab70480a0d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63f69cef99a90b52246e209dcab0e9c61b700f7d0a30c6b10c1a58c0fcc5d8a1ac797d5ec77c08d1a9b52cd428e53939503510d2a53b65;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10a509d99f57e1511cdd79e8df0b90054139b558ae3cbc246f2be17ac9281730e86782771e41b95483112f1a614a8de48906a5b85e17957;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15471293308432bfff00194b78d5fa7658b8ee6487bbff40f0f6728b102b32a28a966e759a95df0364cd7e434b77a09752870466b05dba9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h688442583c5c83ba25658f4b54e19ce36dadb6c56b23294d870791ded272efe6c81b07f27ac234d2c355c83400b85b356f48cbb20bf4c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca0c15b809945d11ebebd6393c33ee7bc16f3e20180ed560ee2f20f43a237c36ce20b6672309ea37515428f18dfe7893ab0c5f090c677d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13719b7c18f4da5a84c34fc9c41335015d3adac3f4ad16708667edca4885e1bf23aa8940d50c54803e1fd6fc7e94568f25f592038a072c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h66a01dd179f9f194a252af457c3229d0dff79d84d5c35a62d3da6bdb796016b551b5ec982b15e71d4826eee5a8f02672ba5d6bd289b981;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc255183b5f68f444c02f582d9741e374a82463a2b119071c3280b1fd50c887141cfac6c3b2e5d34c9ffab6d9da3b3e76ce2fad0ada201f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9d5042f4f1fa96caf52912ff033c4ea0d1820a59740f3de15bfa3cbd28902101a73005e4df0984106965a69fb59498d6e18a4e4a0e5859;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdabd9c28dab1c1cd19e7006adc7f652edd0726ef04f0b6af44d175d09a8643e75220a1cfcd35f4edc90596b3eb73a247f8cfdbed7f5d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c08e00e1273955154e858a4c984c11bfa95d517333515a55de68c9a90c16b19913967b202db241297444018ffb949a4c877c0b8ef75540;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc21829ee13fc00e465923f0969e71761c08df264f83c5f594d0bcce1a73d64515da091b3b7609e9c46e2e893ac768d1c6d2c44946c536;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfa0fb155f1a0ea9fb3746a0deed2c4c783d017efa86bc04cf7a493dec25514faa653360f1082d20d3d929a18bd2c9c3ec4a1e436f7d6d5;
        #1
        $finish();
    end
endmodule
