module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [27:0] src29;
    reg [26:0] src30;
    reg [25:0] src31;
    reg [24:0] src32;
    reg [23:0] src33;
    reg [22:0] src34;
    reg [21:0] src35;
    reg [20:0] src36;
    reg [19:0] src37;
    reg [18:0] src38;
    reg [17:0] src39;
    reg [16:0] src40;
    reg [15:0] src41;
    reg [14:0] src42;
    reg [13:0] src43;
    reg [12:0] src44;
    reg [11:0] src45;
    reg [10:0] src46;
    reg [9:0] src47;
    reg [8:0] src48;
    reg [7:0] src49;
    reg [6:0] src50;
    reg [5:0] src51;
    reg [4:0] src52;
    reg [3:0] src53;
    reg [2:0] src54;
    reg [1:0] src55;
    reg [0:0] src56;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [57:0] srcsum;
    wire [57:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3])<<53) + ((src54[0] + src54[1] + src54[2])<<54) + ((src55[0] + src55[1])<<55) + ((src56[0])<<56);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b9342a999ea95de97a43a71bf5f5a849ae3c362e6f894c3ad016bfc18273b4cc402bd508f514c6bd165fc1af808ebd5b30c07e26cd6b7d4d15b47bd095544028f412cae4305b139e2b011c8d2383bdb49b8be452f05b7f664e9045490cafb777bcf29daa281e96262;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8613b2b48af0159c1eacdba7462df731baa002d18b4ba810aa8c74f949f939ca66f37b1c0d282c439461f3cc86ad22ea3c109310ee78ac6167aee664c872caa492aff95df750e26959174466fba5bfb4ea8e54dffc29333a33f4a7d128b96f536a11d00790bdf505b5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ef35673adf9fcb3b2b8424d91f35e401ccb5dcce223d01093bf2952151d2fb31cf6e626eebd5af5b4b1ddaed25a0c031f0172576890c21b8e11fd3b9dcd73872a735ea117044ec5d501e14fc84355fd1a8e0c67d2ffd6f65447cb76c74b793ad7183b687234f9bce2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b3189f880a76bfa48c478afd88c951eb41db508dff75242b751cb3698479777039ea8f349c30644d36ee9c3bc07acce76970ac89d2d1715bf850490a93faaed3728579ec415383b23b35c802ae95deabaaa0fdf75a0cc3ffd619017bb89fe341e75b225b44f2476ef1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10173c7b0215a1fafa55c5f7ee1e8dbf236ac6da49b85658b5707772c81148f58fbc17491a39f085adba7273a9181f556683b97cb46b4e57bb84998e8f85b825f602cf681351489edc96391a3f3e8fd6864a4d848cb18b269d88ca53bae5da8209c160538b3dfee1c96;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c9d6eed3e74481f61bbca5c983ca74e9bd9c4d4a34065bbc3c2592d243305b48448389d331f5657a3c0d7a862081488c5fa89e9be0b015323dac3516c521d3b76898e34699c66139e79d4965f33c103f239db31e4a8681d31169c63e15c9598d564888939e48cf4a9f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8973777213a2a7e6f55d15ea0290efeb2f5010369d5f8281d6de313737dbc81d3a09cdbe2d1fe876f6f5628f514dda4f2c0c4421807817ec4538948fb09a37db55b7cdbf773fd7d25240ff659bd4a4789ff021fe4965b19f6577c32077f746717db2fb928ee7aa2335;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h132e14843a33b03eda8f6984ef96fdb8f45fb30f6e833b2428266783419c59c4a94ff9109e11a58ff2b4f453cf8c0c66a8d930a2d76e0fb938991a1d8cdaac36b37d2736ab8fd244e69c63c4e7040992ab3e68cbda995340c78cc7024ddd6285c05a70031eeb9efe7a4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3263cff3ca2adbcb8bca4098453e85bcaf09ad8e95944a9f484e58b7bab4c135bd8991538124576c4942b7d034fc70621cac87ac4ae716e969d68f637b84ae564ba86854a7236b657be517340cd23d5f2c13a8d2095003e633e57e409245048b36ae702be5bd10cba3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dba5ee62d9e29075663f934a856d5537885e0143c8d0b97577bce9a31d1c378a8e7407c047a2331fa1d55b7cdd31a137144ecab4aee37a34bcd0ef4579a08d848a894b25eec18b072f7f80f500b570d5b62d0596c8d33445f208928a30981566a68e722dd6af1f095b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1245c9ab3c4f1b840430b4e4f719d5780a98612f117f15711ff76317f3107c685ef15f24461019c2bbaca2eff71d76a532904966493f4432335a76ee45a3ae361f89600e337b2e5f7352364a786bf08fb64e2cf09588beedbcb66a6d6594a09a60b15813de6f676262e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h55e67ec05644d2b8faf408eabd24a3bf4a87d268f29b9562fa5e58d715dee7ba48b1455aa9760471e508b843cef97fe0841517ad0aa4bb3ba5dab229e2914ef2e4aa094fe2abf26eb3560da5fd26a2b18bb2503a6a328323c3426d426b78f5c8206f13aa6c93609cd6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d59c6acf704faa422ab979f07978e44768c9689114219a0a4d6545c192921f82b6992cf3e430c85bf8c7a3483d45cf0fc66e84346132cc3022714697187cfd55fb90fff067f10f7a1c63276c0faff30029824a6d75485706e8a6f7af1a5e633a8db40fa5ce6eba832a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hffe85fbaac70018fc463a55d6123ec2b21a52e2fcf493d0744130cfb436fbd1f151065793a50d4f746eb71e2a60169c7b44a46bffdda099726e4c9ee77ca884d67dbc98c1d4d2b06cb105c08ecb0ace7b45c21dc1e099e46706324639ecd2a2a48e91b1cdb78c81262;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e9a906be0253a158b46a65dfd2e6c0583d5877ff774f90aea4ef39ba81e70684def0806a75d4c19e662bd951eb38a29348c55ded2a64bb13e90b2357f74bd975cf392c0c8dde67cf515b8474e2c00cdfa40b2f0cb8ee4d86f0ff35dea07be0bc8acb2794bfc842303;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db8f1baed5b413c73774deee8220331f8a9584131e41e53f070a2b3cb01b313550107f6fdd470bfdcff1f819c862f1ad03dbc5a4e11b62c0d1983c55b690b29fa50675840d68145751298ddd86a9ff6905de27a0f4021bdb19739e24f313b4d903bf7c49c3b4607a93;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha7a6d93087787bd62e8f23b32394aed59855b6c278196fa6d4b84d7668078acf981c6110887048ed296a3ad6e74fd9512b75faf220dabe03fa1964af3a324225ab0c9ad4e61ce757b755ae186d903cb4d00ed6138381a20a3e25d61c95c6b63232185fde8e88e7d1f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcf592e879dc644bcdb05e028e55862dbcac289f6fba1b64c98a28ea553bb5df6de0efa512fea794dd4fbceea4f09446dd6b12c04d4189a040730457cd7919eea3b82ef736d3d67ba7d011d8aab2e56c0c19aecff005b75bb5a572a94c53e9d29d39c4328b9bd4d1eee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h68f94bf0fd1cfd735b636286d7d50974259e8791990b47eed8234a5abdbf7249c42535119c30dfb5f402f88963f9357302b55a4f21f21dc24e44fd01f010f832091b0b646d52d770022bda2a9090adda7d781304112aacdccfdb44a64b6be9bf45860eb0ee60f3de7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123c4c91978fb7d4a7153b0f373303d17219ebbb4b48e5deb03fe7e55a4dee9e55d4eb9baa2217debc573664fe0679e49a07b226d06ab32966486af1f285c5c9b46225a08a2d55fb82e19b911f7c324bec72cfed5ea7b8ba1a7d500aaf12fd5052381c5a794b99a6c46;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4961c1b222894da246ddea8800bb05b87a623454be7d80a01c63d1ec482d00c86305e0282beeca43b47088a35828e721e69a03943ee2165153b163970932635594a9f09e4926b5c86c00b2c670d5cb79253b4438ee0cc67ef5d7c56924b88b0adfb2e4cb18a84add2e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h127d3f28b840843935dd62c256ca9d881e6b3432d7b90dd924a1ee7755983b299c99659d2850d38729c55cbb433d99fa55f5c19c8c46d416bafc6dbf2ad75069768d7513ef9f3d06072ede12ece1f7df55b667e4944e94ec47ccfd7235368bcde196f6d9a8d4db21007;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e70687ee877bb465557913954892596ec8f1e4bf82d7d0518cbe706ec5c51d405e40f22a922c863ccaa053397f294ba9a6f50a7a7996fc0f8ef8f031478ab27c16466ea8ceefc99f1826f37a1c83426415f10a4bbf0c2699a5e2c4dec8c2fd701830142898b2bd0200;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59ff2f5e8db932768b47371be07815f74b9531de9f220e384737091a7a8d99c98d44c193a009eea77f884d5ebd22f72edbc27a5ceab23b2e0db55ae734ad28962b703e5c342619dbcce253467062944af6e26948cbd6d643eaeed8c3e58943a537ad8e51a680c43893;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1452ce16589b098ec0f613735128b567c5896070399d4f57c5bc930745472d5223acffc1bb908f8dcecda47f38cf6d2425beb98aafd521383778eb8e241dec34fdf9a889b203424805ae30e29588ae9694e605e154e7c1f381e5c6947eed28da65da4870d88db35940e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a31977874d109ae702dfb08cee86007734bdb8a96da39201a1093ffc2db99ff152cd867409e35d3a9c7fc4a22a0c012acbe447120edd3f28637b659d18abca924214376345dd7a0c6a5d1956182409069044ddba5630a106ebd8998be27c7788cec79747cdb5f6fbee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heebe374d2f1cd01c601f682ae7dc00e9b7e9389e9b9b02f311f6d162f1715f9980cbf1fde02dbe8338f39ab87c697df1cc8bd9f87927b9ba7a7e1498f3f398e176a5eb612cd8e9e44925bf6af1f1bf0803d717649da5023557870ef3c1cd060a7252b1102a6023a951;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1251aace093b79d932ff542af90707d9054c86b2afda716db12f16c5a6e90ea64cf3820f00130c8b63df84cea8f275a67a9a877abd83b32f031da4dbe141359cf67a420d00ba29d9ace1fc73b4957f8a0ed07810941a330384e1d603151df24083be559356c54c8b56a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1660bbf9cd3f7e792e8a01b4c439f0d2c13ed8705da54b28129346e9060de28f157986012b740fc5f303a4631c9d47026acb6a7cacba8c3c654fb1b3acd446fd23c26e0571c4acfb974c07e077cccd232c829cc9344fa80d7a332d331034621c6c61d19fd67932cbb4b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5621195c1e77e437d824ddc2f14199980cc32e7b35f5af74dc3004c12a236af4a590f8c411a7435d89c924fa9f57ba3997161f6e8bbba5ecd5a9b8dc40efa926ec56d333cbb777f4bf54d9cf135fad303ab8456e0f4ea9a225c1070aacd30a85bb363bbe54fbb00936;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he192618aa688b98ac0444a075f5fa0664abcd75d0d790ce69c174bac74040150b890ab8a9325b7611f458a455ad7bebb79ee376609552a00591b136a7fcd9b434a8ecbcf978633440830ae73953a7f054b2c40f9fc52c480ef9088f18d00c5e24aa4e4b3a71ddc68af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17ee5df6107adb5bbf61383771033f39078d93731682b92d61d5575e7fb3735a43808cff2fc5710d1cf87d7ac59906b6447fa0e4bb9add6806e2df77376d425cec445c7bc5f06be8935d38063f7c07e404a8e21518cfc008d7363ad0855bd0a83853992788fd1d6b695;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a19644709be37cdc66b6d083d6785c9b5bced4c9060e2c2474a5cc4d7bb09986170b6deb8d65d415bf8e9f5869e9c0bef28201433008b689396f99523321aefad6d42303452d8e9e687fe359678a4b1bef2476003c44ee803bb7089b636b2cbef8c94c9c61c11b36c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c00727a2fbe81e613b28513603a9deaf4f23a9d42bf7c60e58730b91fbb625f43e8ff8d46581b3345ff02737feb068ab9d9707b03168a73c7ce1c084d12ce9ff29d03fd6f809d191fe680985259033a4a3cc7e762367d6d9b6541cf19bbedef37b37d8c80d23e2ef6f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1946aab8109e1ea04874818f7781869b118b2eae5272a0c2427280d80753ac7e0c59ba6c4d8a68e85998e444a9e8f32ebd271680fbe7be43b96c4cc4574b916cdb0fa8dadb2380e79876c9690a5ab76c057da5861174b79e0fc228fc8b84b0973fd21da2133c9911f37;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aa2eb11f413a6af47d906826f2b972e4454a7cac41420e48f25b312798d9b82003c69ae5e152dad07a7c8ece369a4d768f1e8734ec78d9c740e833f3ac60a9e1cda8cd1d750377900bc6edf8355dd38f049241d043cdd1b1534c5d29af0230d391b5558ddd234ce5f0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h94f3a17e6d1faa13ae5815d862f85b29f45e1bedc6dfe34667572a75ac39e2d2a7e4b3a44cfdc09ac36ebf03ea01875f10e10ccfb087dabf920e7f3fdca7c65a71ad08b116e0643fc5b3044425bdf64e82e420224085a81d3f1db427607509d86c8f7a6a3832dcf218;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb806f86d461d871d69fd5de15ae560fe93ea5078a5d4d87b15eb23ea02a0d57225d8dbac45801fa849a6b73826585b1dd34c63f692830962ec11dd7c1182c719f44512ff1366f947d4bd3aa23756c93c29a726218c0595cda0d0add578682e2adce0f4a550a8d426b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1863306c2b163fef9ee47863f54959509a5f204ab36214357cf96d86eeeba7ed6f3c306ac8bb38fa1e0469eb8c7d0988829b6a36711c368f9f8024b2bb9df3fd5beecafca98eeb66ae12827a6e0f697ace6a857d00fb2ba868bdf40ba82bde8e87292f23c642cc821ad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1313ca1eeeb3c204332568c87fce9f22dd6029e2167abe390da1289b06edf5a0a4ae504c15bcedf601e3206dce84139ade024b5563a0b89270a50a6f551b1524da315a536af0370db2496630258234ba68a50c30a85acc7a13c2e46dd57d5aa8e5cb02104ad8714ab7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he801ef3fb4de233fb7dbccddf888fadf6870df2d2ecca24601efa142d7e7bcabb3d7b8799bf4a55dbbeab794cfd9c6814ce41b4f76623b31ce4af570b1f7973886348067d09571af73c53f0ce4355bd498498d068af7c7826dc4b3407c49354a1372a3b6006b11ab8a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a3ad3d4d644a73a5763060b95705a68d44d6c3fd42a1e3d207ab40c4280c2915bd08bc88e97298e8e769c845660b2221cea6bfa1478b35dba0d846d60548836fdab0f23be888540553e4e1065ddfd51bdf2e4c3a9609aeca99402d591a9c4133257b87c8b41a2271e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c8c29c1136e946cbb991740fb625fa931aa2ee30aa5114b505f0e210da8fc6e399ebfe089f1301d1c45d61324b11aa81c148f4768688ae884acd920433ecf622636f997a67046056f35746cece06ad2aac992cf65edc21445f9bcdcf92fd20d6a38e84b7a49ba7935;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17a674b6c8a3d4e77587c7763f4fd615ce495a836f511c3d5ef59f512d43800ab826282abed2390446475675df81fedcf8e2834f237282b3170b02470093daf0f99c4e96d94f203f45a51854d495cf0286d198e1ff4e2f0601a4d17ffbb96b8f2054499ca577af27af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h405bf8d934c1645a577f6087c63a99f469433147da2690944ce4b5ee4b6de7ff77255f9ed49d89e2f30c3c8d24c4f77fd2920212625e7f36ab781dc995fbe31c7205c74e34405f7285244ff5d6e717e664ff6a6b150a6f7199d4420b86a0220ad834ed71b682e5287c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb378175b6ddeffa960a90745abba3bdde51587adff367c3642bba0f85765954acd4e66075e7008cdfe087bfe0b66f87c66d580ba3a3befebb87faa9b06ab2cfcf7e182535d05e620a79a9311665b3f2b11ea39244c78867645b591c5b2a84082474d8b7ce5a0ecbe95;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6bcebfabadaad8128ecfd13b3a87c07daed7693d4b6d5c9b9d7b991cd8a7019bbfe5a560a9667cb9b0654ad63c4f1809e12e1258390bb584ff0bf4cb32eb7c1fe00dd537e667f29f52a94689293e24f642020b32f984fe22b621246ec545ee117102909872ea4c69bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c465cd9bba263e51b27b48d68e95944c8f327235eea175f4c4ee3e352852609ba2c0ccbdff0230ddaff1cacf9f60bf91ecb4c9b78e9d926dc086bd1b48de7478dfcf2734c3edcd55efb75b6d54cbdf2e53a100a5cd772736be71821b408cace5ba97699d21034c1ad5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15e74fc279a652325ea13be02cf767dfb1908e1d5c30b1e2e8ce7ac696bd4368cc54045b896464b28d4d2745a27120a96161fc641dcb8a0cb4bdcdfa184c94393771af78ccee655417edafc7a515bfaadb76f9e03f0f708a2a73225d29601be8861417e51447071c056;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2751048d9b5654fdc6dd3ef2e62cce91439a5d3971113efa80fea1256a546233bb7f8fd35feafaea2ea3c94a3befc6e19e5766b8d321188e1993deea7c2eb0c4de17c37f5800453d077f5986e6882efc857a0a0ec67a6cc0a47446f480d248d7cc3bfe9579b583d61e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f4caebe7ceb4e2d8e5c5f2b175efaa182a0c0e5790d7516471370c0081167b00a7c35e10e5223c4533258e76bfe1ea72e7868609b7c434b1ea71c7fb44a500711881117e5174dbeec174d28b532edd848e4549abe57127d15944f82aa4fb9e7dc0e41de3e70c61c50a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac1b1f803cd50f9362dee415803852dc450aef1c25d8d3788ea4ba283e6e2c8915082e1c12f614afac501841d6a1d679ad700f92e647ab8a231b73fd0d0d537f083707ace615a4ec64b73b0e8d9a54b6d09a05af14287561a29617e335b1a9bb8d8b80ce0c07899c86;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h61a68bc5702f0323a4c15e5cf7d05ab8bd34ed4da2727e05e1f1b9dde58c86454d0be324a4922e5662254c95ba308c5504c5d490fd4c2a0038f05d5e5bd1791ab1e2597b9ba61812b973d5af02e0f94722a77c2c106d632e0a83c088444fc8e9c0b52fba8d24aaf744;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc138f8694bc65c81e5bb948a00581d541957171c5111ff318b486bf73b47582dd87933434130b5dc3cda167e75b7bed831a90eb0a155a678ed106f09b1c7e8f5b0144add86940c6416c144a987e5a73860aa6bbf6296c1144e4802a4809f762997a2d4674fb5c1287;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8ce822b5758a0e422696e503bef7e601275b310cd929317fdb10ffebd1c4fcbb163945c14acd4b1b768de12aec3067f47cc3461a1539e9027b95d535950b26560b188fe5a91dc6e1cfeb1ca7859c34976a6f7534a3579c2571230180a07747457a2b82cc199211700;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b667138a6ada7e91ac04b7616d49e81318bfcd957561574695459959d6aa736192bbe81339282e27cb6ddcda91a91da9e5a41f1dd72210fb055a3115d595d93a11f69b1413cde3ca04a86508df92a8ded83630faf67b059e678d276a4c94d0d54c795a26a3f0940c7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67755e1721dee955d829f3c4eae311b0e4e5a4688d7dc4603898b1763c72afb251af49268e9dc44386e04ae74d684d14fc66a9d4143d8fee451b37c463cef5634f9133491991e3b1a6c762817893f1dc958c309817692d1d35b3c301a4bd2415abbfc4eccd0691b706;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h131b467adea58561085028275af814c15f38e3f345c1dfdc1da07918565d527002a6cce4a36e0af04300b480bbfac2fb5ecdfafec5e67137bb5d56f5ccdea7135e8e1b19d020e257af6c07247d976a0dd78a179403478cbb94f447bec76f7dbb3d2eb02f45c74606e4e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e6147995f7713faf33fb5732daca18428ed084811dfdb8663bd6adcb624d01cc1fadb62aabd66891a85ddf04f60141cee2d9f302f54236284f8357cc1763e76a15730572e36a5e88ad47be63e96d9a781d50aa5872f7aeb40f6c5f756fb18f9f34ac576585b5b3892;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbacd4c45ea760794ecbba8ae79d124080d48de922653820f6bd24a5f26a4db4749f0151e602a128670a36ab0a7fefd72c494d776b8c363c8b0d8f3a5c031aa3cd9924cb18caf708ee218247d3be62ca106416c284f3beafe854ed8cbd803bfc630c6c468174915c910;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcdc749b8d1d74897ef767df548e00ec050b205868cac3990c3b027653f088a0385556d9c77fa0642fa43e51de0971671b4e624d09d70c77bf07aac7ce1801df52169e572eca10fc4f4d05bd48bfa0abe301b637df31604a01f7bd8310e9bbb1a0bc7bc7e7c9b1893a8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h61d37a0d69b9124864ec3433077e2d03d3c4e71e9f8ce4d85d3124c22695d64248ae6e220d794dd27a3569e6bf530596cb873f4f528cf3ecfb51b65633083464d09d19cbeed849986ba00b287400682048bd79af1689a221402096feff7e0a1908d4da06c9116f256a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h80f809d193964be164a16e281e8cb50819086f97b4f0e190647a7597c93844529bd7837230cd55e294067ab6bba1d611d91ce240b38774df80f0df05c134fab83bc177e021697807e738fdf491544ba1721b68d99a7541dd5ce4b3a5ea5ae1b0b3ce55051c2a257377;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1178d16c4029f667a3a4bbf94558e4af753bb4877fc2e3d147063c04bee2225e8f0f97d29e3ae802af0947319327862c0dd2696ffe32b8babb88927c7592e6d7953780481bdaf2b1077d178de65d5ee2d6fbeafd4f377ab08a5686afd8db566016914b2bccdca9eccf0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d755d8f735513609fdaaed0d4c3454bdfdca683048cb3a35533efacf58a4830acae39b3eb42423e055aea3e0aa69fdba962a646b6ebd22c91d4c92712214decdf3b2f809aef12fcdbe12a5d18ffd0bf3fed31ceb6e9bbf61e74bd6f093787dd7f67a062fbb12c2a617;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h808c9104c030c246879d5e76ab15d82cb79c7ceed98112ed14230f73d7af51ba28e6488254af14e552e5e3bcef36064c2795390c46ca464b7750638ace19acb2a6b02fb7a35ba3c5e05091ee66f98706711fd16b85af6a855786f2e677b909a13ebcc8bd6c27498d41;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd7605372d2d0131f94bd2a9a8835ee59c18a2f09983676c279b2e090e6aa43fc684266ebdc36b992363b5ed272ea4836d8dd08ce6e489383ea97d1e619414ca7a8f1cb6439bcfefb24cde9e9e88b4a91338051210307ec9112f802da540cdaca64d910bb960f6fe48;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd64d78f3ac232a960c785a9d9ed4e05f48b72d431dee80da56039dc4b3e07c1dcf3a459a8b70faec716598c74f2cf5beb93a421d450aa80ac39cd58dbd61b31ecd9d0b61518db4a692545c2beaec4cce04a3775fb88638d0bcd76c6527782ea50b2a617fe5da6947c5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h119ca30beae248b998799d8be52e4761f8d3ac97d5bcf0707487e3ecc7a7d1ba342f7cf066ce91dd93d3bd04a897eb86bdab47b4bccd239f90d0cd39a2a0f81c1d377a3b5289fd612ce1e150d7f6d400e08df4211b3c7c9979c8a42e6d2e21fe015fac1669523337b62;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d6635691ed709175fb620d894d0c9080b08b7af72dbff5552f759d5a94be6e0a232d9c5040f31bf6ed76b214479a2231682d6c7f7e85afda3d91d9e9dada7d4f6a590ce089112e925b37ea09eac9ac3b0e5b391a7a8dd0eded809fe410b7a84f5166eae00565e282b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c45c5781e2f39ecb5b4b0d876b1fd41ae0647d2bcfbb0e27b405254c3e613b6d060cfa4885695ca8583cc013ed8cc269fafc3b6c07aeea575ce3b64f104ccbcee03b6074ee584ca4646ba404e5e18dc413d31783f65f386579e30ead801bc92a48c80df875f8998d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he5b6b9062aff40b366a66eb4aa616ca267a1d1290aa39adfbcef894de3917f3af6378afbb72d25c6a7246f51436038dcf61c83ee66493b2b964e519b0f735249b95f5eca2585086ec2562ba59f477c820b4cccb8e69409b93840083b273b5d02651fdd6fb2c03bc94f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c5d90618a5472e95b353875d7a281eda65eab4ce29813b76432db745d23ac3d148f5a13600c74bae86f2439248790e629e69224d982097e2df628de24e414672f61ceebe2268f107f76a71a16fe8137009b0a5f3157d189593e98bedc53ec119bbf7e58a28889a1a65;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cd7709848a7791e2c4623efbed1377c20ef463709f1d941345bc1c115c2878f192f692ec3fc0969dbebd8383007567e6a49dafbba6f4bf2deaa501feb3f64abed8f1f80bbbdc4d037a90151443260ba7ce69ed575424aa9c48080087dc099d9465198a356f6c70363;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8cf35a7fd6278b7a91ed81fa62463f52aec6aa09c77e396d33eef734b90671bc6b83bd2993cdb7e5e4fdd11f71c9a2ab6a31fc1f320fc2e3b76c546810e2e2fa5fdeef507973b09eb04bb06a94aba9cfb1eca6965fa9c5e84139d142d9b2424473f583aab1cd8283f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba185b66ad680077d64c219d93bdb1971f7724246c7bb5cc3866504afb60445c69920e9d8fdb7de222bad0dc5feb6f9ca4d8fbc776fa5af8e6495cbb78bae53889e1a1f197c0efa05c1687cc0e00cc2c248dfe5668735d36a9706420c3da3f46a53972ccaf92d9888b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167d6184297e69dc20e298e9477489369edbecf186ce68b24e01b70b340ee3ac836db6ddf13a9dfb3c7516b4b0c57c9f82132f5a70b2efdb6f0bac7eee85cd8b813a334767b35199eeb942b99028be11bf725dc6d9d17a23b4188666c8b2af29851f04154c9112c1f1a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b76be2890c682694e6765971664fdefa7bd3bfc024eb6a80574189bbcb0402a69c50c2ce105ef6cd99fb77b2459379a8631df828b0432358df6b12436ff8b2817c720a2b0aae4c0232e06cd17599357d8bdca31862456baab56d704f640d123c4aa53b0380e8e7127a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1783e27cb03c378bd045062e44734227ca5fe9d98d12e43216cfbf7ee4e47cc7723290d81dc8b4586669e9964fca3baf34085db8d25ea1ec8c00995ef65084277ce034ae037f33afb02ee2d15adb03feebdff1b9041dc9449088da9938da16c4357045782ff69b0544;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14e88c5d054992ff39f8c9e7d4b37f795827e74ea52600d513cabff6eb93be0d52087e88250a124e634be9e7fefc78dae3395a7d8ac14c8f47807045a253a7cbc79193796722fade7611e35e5162d76b67fbad5c4585e6b7afebe5990b84c1adea74c0ebfbb47905ec1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1acd368ae26c49e2759196720224bc2845e84b5ab439bc558e59418279bd34cf365d603ef3ca03b61e1703ea526a0e2609ee6c174e326499d056d6f4cdf172423c756502fc3209ce9d7068a0bc803ad48698a8e88b8921dcd0a73e24b1570ed60d7dbeb235976c6003;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ab5009b654212f1a1379e12f98b67ced81f79267ef96bbe8b36574d21a1a9473a71e0e77d70d30b3e1fa7b23bb1102703b5bb44533238957ae03dd6eb34cedaa2517817ad539cdf9e9614472a0fda28311a1c54ceae128380f08809eb5649b135de1c8aef7a993040;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15e332fa65f1a508be0540c6a426c871fca57c7d8c1004fd69985e8c50d463769bc6c569012bb7a3a54fcc9d8f72bdc7c24c0d8cce8c9cb73104cceb1936406f4dda6de4be385f6633b3b6b8b80ad6b9d12fe73bf05a4204179b48e3faad1e27c0bf95e3c10ed1f5823;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183ac7f3047d97487fe30e67e558b682d83de142e1eabb8869718a932f9815023debfa7eb82e0f4848365d837417a20a670f57b99ef01b62764764ed4f5ab333eae56c2c4ee52c6fdb81213e52bb51cdfa9965c3a6564a64055c83549aac965a29588a64fe6142ecfd5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h33ffd92275e815b3c1cb162bea94f237f22aa78d4f57d1fd7209af01dd99286692797d81643d5eb3e1dd40e2b9b98eb1db750351f96ef5f484588954b28091e3dddc60346a56cf8ce1fd2b2060a7c2d7c92e3205710ad802bf234112a2f4716512e397a979720597ce;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8eac84a44342a796ec6aa6de8784d875582acaac73ac97f434d2cf6bcf11ecc85d96994bb5f9fc323cb38b019a9cf86c359b11255a99c027fb774008ecc289ac48fa13f6486750ddab6cb747dee5901d0fea6600afda54d5d4896afb3dbbc01394d10d1412ae600b9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h126694fb12c3a86ecfc4f7de0add178e040bacb3c67dbcc66b94aa495f9cc6b3d021d641aca3acccf0fa505db3c143980501a8a9117b5cddf6b6cc47baaee6f858e028b14b6ee1ccfec26eabe7b3fed869f960b1cda43c40d0eb6bd723b26bc0ccf35e2398e8090487;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c56df320c8d1fbf1bc2ab0cc55656d79b4b9e394bf2c42d7a76e5a51d58f582037276145888ee9fe0eb1c0ea994af24a29aaa620a65669f0d83d3e8f1099201f765a05fdc825a898d8fd8664dd8560df9539c8f4368c6c28caf1a4c2c59dd836663a9e27a54ee89df;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcbcb2c30b3142d72d599a8ce135e9fb2112f5bf93b4b5af0ac5b0c48a77c2d642ba6f4adbbf801d575346952ef545fb212d0c9e932f4d34dfc520dc24232e314c11d63b37ccc8c5b7d0879ee5a86a1cb18301aac9401f7a1129e47312e45626f9abc83a9bcd1038d9f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b7bdc585ecca5ff1fa4cda0f57444fdd912402704a070a1205eb96405a51545bb18260dd330e51d6b7000e81cc8627ebb5f1b147b98a29b30f23d1a507ed75b4c5e51d25647403f47553c5533743fe8a6cae3ebb8b815353b767fa4c4268515f3a4a87526e4994e1b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he49cd9cde1772053bad7c1a6f44c313113a70bb3eb7d44fa2b2364548f6e0dad48d11b5a35e412cf1f186c430daea9405fc1ac040bf051941ad646511505c346b3a9fe6a9c244af44c56fc442da54cbe98fe8320bead929e9703665e709eb0c70d05bee9128b86b27;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb69de78beaf8c116ab3f2a9d9ca3e141e01d92e03c0c29f1b04592b5ee0c711199d5c770c6c93792c25b6632d7712de663713278ae13ec7eb8a03246c5c45bbfdd1199f3602cb277a63b72a5afd10a5b0c8049bd8a172c801ce1940131dbf871e1c0ee99157b7a8514;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ffbbae5ebb937d1601e4fa3ad6f4e2a3c19de697c815815ca9c1820ed512f4b676701053daaaf07d1b5dc69e7ef54c50d11c229413521cdc4dc22a01925a17b12c1f29803298006dba2254e0ccc8de364f5f9162fbe79bb28ea34f196194d9e5273ccd756466b35df;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18fdaccdc8fc026a283830fdce7ea88c4641a71326d712ae26b7419a964da096070f019f234b6b3b31dad93b50a86c312dad48cc098c6dac8e9ae04267443032b75fbb038e396bc00a928e0ac476257ec9f3d4a130125f8c9fd91206b01d26a2cc6cf6e26182fbe98c3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h440efdd05a6c951b917b265b01bc93089ab451e4b70504f2626a0cfd9fa002763070af92a23f30a2af9c47e5f1567c9d3e5290c68473ccba3e1cd6f878e000afc1ca57087af4230ef5b23108d87eaa3a57a23f90c616a8e90aedbfb6f6d41ae0d5b3b3316f52a90b49;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h644eefc64d0b151df3050900cbd83aaed50cd7bb4030278967a0b705d5d2ac89668be90b877edf6ea266d846246944537a2145fdf41d7c91c00d5905f21e88e309f19031c0e66a0183214433c75058e3ac99f44ae769645aec22aad86857083db635ee6db5a270fdf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heb5e501e584e5e882524cc319cba2984cbef9184b2f31ecb8dbdf461bdbca6d83697e43e57b6ceb0468f90f6ede30740114e79761ae4aa5d4cc3404265616f808a44eb486f5e7b055b9af4ecdc711db52e0f642dca87324461cfaa768df122d4b5e93ac124bc2c47f7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8297ef71b825c64772a297d9d6407dbfbe29543617ec508e58e52b3f72eef28eb7a2e89d54dc060fc8a27a2d99ce9c8ea5ee0a9e230f08d5677d433603a426e99be202209c97e0e394ded96e340c28d048633c006a974e66281d77ffe2ce3c14ccc1d543f52c4a0e21;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c2f352d6a415648cf4db6b58f7437163c13e9c001bdaf04552b8b2ee4fde8a468a4da13180b69ef3532e5ea67e8fe7e05975cbec907c767d3f30e57670b47276965688ad826c190b2ac870014e1da724a4edce76aa2b4eeda00ecbbe0145bec629240d3fe0a5aa2c3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h151d624d87f5318fe01a3d1e103d0e2cbff69bdb4bc7578e694837c6536dadeb471138dc6e3cf66a84c9200b775497cd15302e5856bdae79686be4ab801766dc4e67804e661e7f62d62722e2fd838fcd0bd9497806dc94161f60bd0ce118e70c1091e34febadae57ed5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eabbb1222b42700d99bc978c72b733ab207af59535376992598eb01a6656c879ee1945c8abd08520ea9bc06211bb5a5e0dcf3192f54b0e0d605acb4b02234de9550b394b22ef307cd989eaa7b60c67c97aee9b092cd3427f297679ed7bababfe355744390d21be6b0d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2906ed165000fcfb071abffb0e185a9c6ed2c18a25c992fe3eb6c6a7d53fec5876f233a30b2aa86cd1a10ebfff0be4cf4ae2af7e978a5089c00c5035973595bfe5d5ff9b9c00072ea5e828e8f8823213e18c0eab07cd232d6ceb74e6a5a7fbde61c920ab009c0ee04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ff00538e3e9eddf50ce6ccf5c7e03a904408d515c55192c628944e29bf6f3b05a96b14bb70ca3118ba0385f040041d800039f20eab8a630b36f2a5d8726273e1f2d61fbaf22b1a6c7a032f4de41e881bd10af1340ffd8e63ad32c1016b938aa3e5c6c39adf568e787;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f5dd728a904ba7bb93aa6b317d8f5898538f833d60e3e56133822d21f66010bba434f5c4bb0fb67cb88b17bc00816b342aabde7f3b034cfd91a49984e7d5fb46857dd7d4007779f687e571c4766dbf782a8829ed875e6fe9ccecd5e8263f82b42a04e553b294c8102;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d3a279b7cf1ea5c1b6317dfb6612adaf0cfd4c80a615c501f5fed1494f5d4b3925263ede71a1c661890b171ea6388699a5e650dd3f218d68306cde33159c113b0653b8ce7960a3ea330b106b6edecebd44e19a04c2906156879ff326fdb497843b2d518ac3a4814ef7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187e355e2ccdfa002ee19e6559d71caf511dcf35a2912bc99148dd4864b71a3f2eb297f05c69c4ec94ec7740d21c7fb76ef185a883fe45fa551c7d3b5c5b5c750f5dc1b749f2d1a12fbef4200604dd7824fbac833dc45c570df77e374cc7c07d8982b8f19e65fed1dbf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59111556c55a2584098d26668d67fa4dc6cf3db65682a88cf4d5e549436cca944cac9e2befd4f6cdc1bac8354db5aa8c8b4bc5377b3823064f4bde090d0803912c9283e2e168e8e50996108bb3d658d95a5929ac999513a4c57d378c2764bbd4b36019cbd0983a5a61;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18df528cef9e4037dcda67a1994dc4fc13f45775a829a64b9b5e00bd6d8dcb644af94044686303e0179b0b3b7901c836c38087b6f2d5b380797975484973d22d5d74f7361884cff9332250606ffe7dbf60154e261145c4011fcffc0741efb5fedd7cf5bb2cdd0f3e645;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1403621025e3ecd2568ac974737b2c83fe91194ac387a9b13d75f805ed80143ea2625b4cda247a7587fb3354a1adf25766cec48376155ac2d4e15032e2a9877f6355ba0d1719d1f9bc36ebddfdf439b03d8190c01391d8408fbc206e5800efbca8f2c0076f8bbe7914e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8445ac5f6db4b56af45ed13d3335cb3995a160ccb5e257e5d43024c7b9bd92a71a2ebb1ae2cfd3a19021913e48d54cb82e98038d7538c89dff3030aae6056bd963a67613ed07b7cb94b1f777a9294b9ee9ca92baf1149a4eb2ec9949fe9ed0e908da39dab801ef147;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af5bc300d1906635a066b78b4a784d44cdc4dec3af509a6dfa9b371c07e874d8c02e3bf9f74f73c5fa8a4059aeb67626bb4be7e04000c782b414f4d33e0e8eeecfc6e8b7e324c9f60ce8571d77d9693589ac286560ef148969e11b977d79b25e429d8458f85c42fe47;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183703cce2cd7d976e6453716f4633561a3fe3b4aecadc529c6d609548fe2323fb890deff7a6cfa9add326ebc1e4a46a4a0bc21264867dddc5b065c6297dbcdbdc2b141c6f0688e122ba7c5ee91b333b8a711cefed8211a055ba49044454eab21e2f7ff818e1c05656e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haee59b7c3adbc5204b8627144dee058dd673f1cfca9a6d8d7549194d09fb1656dda4a8b5277f8a5a4a48a17182ad2b211269b0a4c6edf66a077b83911ec7ee85354e738a3ab06c47ea89bdbfcbf6e6837249999667d2fac8ff6b5c0ff981e4f0e1baa08a0e3983051c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12b5e5a918d35d3e5a1a84b5d9973eef9daeb8823afb86baa9b65a15ca1686d507193aa54cfd48314a5bd3f581ad5481b81ebfb78b2fc880755d51e7e8df75f27286de8f11a3d867a60a8fa26cb52bbbb5e5ae1e7074da535366cfabe7319769066b7d17345f04edb41;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec4803a193848258637c6d56fe4be2700ba94fdbd187ce8947cb7ccea6e79a04635b837ee11bae2bacbe2fbe6a7acdc9f4cdb7628ba2bda07f779c52a7417af24b4ed76d4c82a7a0e20c705f981ccef35377f416cf59ac1b41f63802d9885091021bdcd5d081e30153;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5891f87f7cca6c41310671caad510c9a2b2851e6ab793c79e39c7be19574f956afe00f31ad168b676523ebeca78e640ab8bd4f63807faf5eaf5db9e58763863c2e2a31adc81ca2caf82240b4a842ada8941f69e39bab8f47c74943329f39271f63684dd3f706afccb8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72d246f85707432d0207b11ab9de8fd3f37a31bf36d918e5a648f60c75ebadfa071995acc94edc48005b5b94b3fee40734e427a6fa036b538f9453cd1f6a390f71979b41fe1ee503f2b3ebc72efabc656eb753c9fe5982c4bb7716eb7a4693bcc374eec8125d2e331b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h153caaacac338445d953b53b3999b5fbb5f20d74a1f9f5e4078f92bc6b3b0baad4fc08563382767d5425db5dad33e36b0ac4bc115dcc5e0f72acca0c038735bae7c213b2aa7d9089c8619c18853edca18b25f0bbbdc5c8833b9dffcaf1af7ec68aab1a04249e37f584c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138b3cc317fd2001059b859a5dc0e33d2c17aa94f9edda4589473103ec08f30d783bec855b4c78c3c761f5b476e697a6eb060d2a128481621a2c5df6fbe2eb0c6e1b54c9d66a717c5657b6d982a1df84cd28006fca682a4ff9976a43472291186fd3912da0922672289;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8ddfc1987ab1b993e82c3dccc7661d7d88c62aa7d8a6bb94d52ac2224da123004733aee4ebb53cc1bea21db7e65c81820ccba187f609ed4b096dd1d04e947237eea01cc82c258f3e83fd1fe1433069f730d88e73c839529c7aeff9b42ed9aefc866d47d049ac216a74;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8161d0faf5a47808fbb060f8880c960e76fc4b9260518dbfa60008402ba8a79a7ca0b91eff25f2a4cff7003c4e7dd80fceb7dc849b93ebd6820b60a7128a836551fa2c0c75c743d91da5736d34633b9fd316057bb247549fa4f8d86282989174d3f84f91425c1c79a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h102ba795be82569f28b81ae81cf0860eeadbfdd876b2c5298fc039238bdf94b223c8fc37fed4db9d05d63f37631470fc457e1bb1aba90451775412b97561d47590dde11d6b80daebc36e3ca36d542575bb82c366a28f753b1e5c9d84cbf3c28aa69a83d36a84b9444f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8079171d5a1dce623c91e723790ddf15d6fdc14ec0f2339ae952342caf469d38afbc16e4be96d161bf1ea128c53ec8db0b5b75f4bbedc0ac47b17b18d4a79c199f732b4229f87226c088cd42a5ed43724d898a09de623230505e89fa1aecfb3e2df35e63f62a17cebc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8769e7d24cacb83c66d68ff546a0f081eb044dda7a3afcfb5d0b755da5f843f41ebec824967289cb10f5ffc37f7c23139464836593b61174b39685e57cced6d268c6f8bdb361db62ed14d26aa17e3b431504e55a9a878044ef40ae8da2c0fbf3662c33740543a0b3c5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h128e9daf96b5ac4d9c484f5f18bb5b9d30f4e98c01d0b3a10ab239dead60abdf14590649a3bb63dc7cd6df7f42f2a1c677d081211e9f0345f2a9a9a98cd29e4cabf40ff250577e88b4606234b3db9f17d342420ed5d2054e17fba23fb2257fc8f52d4d23bc0fdfe6a67;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3cd6b3507f3b6cde6fb467345aa9b7aaaded1d020cc56b05472e0d5b2c3dbfdc5074ec56523eb6e3e2fd405f43fa11568230032811936cb342f28d5c1462e3f555e1d7053812bd30359c0719541f3fc3fbcd538e2c73638f5af056ed330e5e7a85b27e5bcdd8d14f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ab3021850abf8dd52478ebeda055bef53e23bb4bcdfb943c89cc124b479f1e1587355399afbce9a0b732ce7c774b13af18af057120badcad0106f594864aa601ceffcaf974b41d96b85e2fe9eb0d66e3ca76419dc9ef18cd224f92fe1dbb294ab4bb69d8fd357587df;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h107dc4e6da496e787107b851dce6c8dffc553122888f6a5475df938f4558cd4445708e4cf73fa8ec368963499d17d6de98ac2476533ae4d6592eaf2060c4aa3f297221b1f2b643ae8fc1a690d101e8d64d95147646f806456f8b197f59556aa9c4b02a765d976c0a3c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h185e2281b38648f78a7bdf7c663bec0c030c2772d46af8e26fab19035f07d1c4feb0d97e4235ff8d7f74e91f77848fdf7e0771ca50f792fef076a02be2e380d6285b552b65f70cff52f9d8e8499af9d81b226f32156838514680004f06d24ae18722b82466818c49f3d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ccc4f4d23711e633f4bdb135f622f33ea7b59a7e16451a97258c251bd7aff03dd5a871872c46deccf32befb2aaad5ac8fabeabe6ad49234cfbce1b6a6563d3354ff3e10266ecc4434ce356720efd311533126192e227800098aef0bf7e502821eca7e88800bdd55ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha59bbb290d717048d53dde01cb84cc1ff2600f0b801ec9f4984a55aff5fdf666e72cc89748b9e9fd0a474400e09dd83fdd57fd69306dce8ee439180238c4d69b7b85ffdaf7bcf1aa3f4ae3043351a07237c8f1aad288c240b9e0819fa76b68c5055c45beaf5c20a983;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8f5a4f3f125dc84141eca9c6a0eb57d9cef87fccf68c8cef5062039caf22a7f26306e53f697a0a3d01b931764eb2cfcb526e1394cc8e6b5b72fc4ef59a480f68a20eecc1f161e7af50222e29a2acee417424e593e563a0be9f9da435b5aee88f4d9e322ba0f4cf49a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h179a1d80e1a43cad6301fee089ff6f12e6de878e8b2e9bb4f21e323a1038cb41ac0699452b9a92420fbe0f6e8094cc1b01c28b5292e8b28966a6548999cf34105cc9669935b0bc134949739aa750a39e4a7149dda5f10478a8db96bdce8ac4e3a7f9af9a9a1f4f03cb0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28767a486880ed9303af65f7982b589090ced9ccc1f4fd63f36c7005695b8c1eb2ba2c7ada613eef8a8b1e495576949cbc7184edcad9114386b6f96774fa9d9d8960537ba4280fb1ef6e34450315a81e2ba31efbcd506257e18bac249a1f5b8b22e6ebfdaa0a4ef0b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he766ac93f3f5039a49300fbe8befb2f7ce0fd0ef4e03e5b755f01c1a9f701fbe58c8625a38a7cf2124cbd53b66fdf16427581b6d161da7c86d9261c6149381a546a38a5a52bc075765c77cad40f7942f1126494d0d363cbab3571447961b02e49f3bcd3e59ed795adc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h78f701dbd6d51a97610a2ac9056838d584682245ddc6688f8a4331c9ceb4e33ee82f7cff6418b64f47168f2bfc350ee3d99409161acec011edddc7438fbdceb6a15a9b478ffa45b7e2476a7ed7de7c20d10a177e0651e9a2c674a012205f7251752ef80543044864e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc1d39088e3b814c114088cad8e8f8ce953d26fd6783ff6d235850fac8a0c3ea6ed25028c66f023d563c4a1b08024175d7d1f036c25e4c8f5b428ea3a8b3224c4c6b0093a62bad0054b87074e739d6cc2f35a3d54db05f3bdca53e4638a5a7599410f0d47776ec1404a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb28cfdc96bc4ee88a2957a30776430994c3e76e7f1a1ba8ec10b35d88a6fa8c731ed463b82c8f504c498a0fd701b3afd3bcf4d7f126da0bc01ffbda661bdeec64927e5d9b778c699a6414cca0d0042daf356618cc67c2e7e28bc856652ecc50a2ec3bb399ad52ed332;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h139ffdb984ede32656869dc9fa3a8c2cd0ee55b5461d4460b8295bf330d03a3ddfd9066fc6c25a8d63a8d13e6895e8ae798df61c1ad8a435ae4dda7641ad1f9695d84ba77bccf008de9c1f8964c595e3092779de4e2bcbfc9db2f73813849af221bf6b160ce9e5b2a1f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f703852e0cd989d9aaec7b245832504d2235fd26ae39836e05a8969b1699bc7ea19c9158f7e598b6ad47a4b03ef612334a16c8d99691d7332fafb79f2fd255195ca397e012312e922c9a28a04e0c4c6860f9aca82fe953f1c589ec7af88077132476cb78ced44039e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c561dfd5422e42a62554cded0dd4f1b5b25edac2d5d65f92c5f762e5f335fcd366c6f9e8d870c027c3ddc53c76b3281d0e2531e2ed3a9d02a234b8c29e6c6ab7ffb42e159e33c38781dd2adcd2daae17711eaa4e9e90177cdadb2a17f7cc8a01c0e28dead31ff0bcdc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h826701b51e830fc2f2ad9a309598af23480314fb24098ad12b81a5fa8ccba4c49f653ee43451e0eae10176e0ab506c046f90d83da81ded78e4b821881cd90bc7b51a5f48fa7a0c6bbeb4a2b004bf6ac8af587788369f219ae611be186f1009a91340b05b09882bf780;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8f7d2ce798725b5da3ccd14bca0748a76089a71ed1885c9f340e6786c2ba8505470c51f8f4de9ffa7f9eb1c958aae782769aca4edace28dc15a8570f9cddb93d6ced6bdc1ab7f73e9597aba32a7f72bb4ec77713b7f1ad73313bc39b3c1957eb30d1d58915367afde;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18bc4545e6348faf17ed9a07a3b0b33d352d9aed3e2f9c89618c826a8169dcee53253f785743d7c0bb4138278373e3189a8757f5e5ae72a3234ae538edd3496687df3752c676b3bba2fa728d6cbf20e2f9fa32627ad31a1869159151e50f2d280fe55005e18e27bc05e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1327a4cfcfa23afba7e95e5029fda9852d233cab106bca4f39ebdcefdb51a222d0f9d77c3362fb24b2c74c3277a4324a212fb0bbb547c75edd073996a89d8583a89c7527d3457644d90ec0cbe0b9cae621fb8fa74eeecb46bcd531f13080b89b579ca09bb83ec0f980c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a98780c730fe1657279eb5e269987a06f5e8febc6f98e15230e2188287e039cf4fa92426320f2d575cf0a7bf3133dcf534e998fa20f9729cf5241c8fd8872534ce9974227823c1819b08407112085639683d199cec414781b1376b4dfe8175d8450cad78dff25e03b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b6e21bf071ae408f75d7e7da331a48c56dd1788f1c58f62af7f9e4e53fbf41729e503c41e9a610a0ea3e5fbf0d218c71839d7468c6ebfd124859be61d31bef16222f31bfe3be4cd607a9a3d2113882f92c931886368172ef91f21afc8aaa5fece258d953999149d280;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40403b9533911c9e32546aab68834744bef7a2ad3bacff927f47230f32c669aea2f135541955f72ce5e93bcc4c43905000579b304c1a955b963377f5f5b296b027164be221aafceb6df53f797f8a2827ce5c3617a184f5cc9e56d4316198397ae6855c2005dd2d2726;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha75edf9286f80850c21f80fb3f115469b3994fb97df32cfbe1ab6ff6a1ff71543533b6fa7fca431cdd012196d2d5a9939f6409aea9bb20b4d152216d07daae53b3fe78b478755189bc02e695ec4abd33d3672c1eb5a58bd614e853dafd6f3ede097fa0377212d92018;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e2d9aeebce4e82874d7a3d855d46f31f1880c28b75a4111c848150fabd4657bda09ac532d41e376db44aa7f0b9a97a182d09db45f216c91d73ab70b1015dbc2ce0a94a3c4d92d36ad504fa5c75fef517459a711ff5fcf1d84f05a7ecefeb1ddac071c3d3fbcbc1ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e38536b6aa96de94e3f6b4ebcc539992a55cc6af53df1121d98f77396900c14c044a28180daacb0e4243241c1eada668705622d891de6ae3a9ba86f30590c816e981ddeb576f975cefabd4c6f84ebe56aec4d1c3f1cbc9ea7dd72f02ee149e42a373cbe2d082d81d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he7c0fe8adcc1ee199f8d87e420ac471556a45455ed4c580511be9e1fc26c46504852a58e6d8895ef442b3e2d17339bbd6a8b80c5a77c503ab4dadc2c3a89518b99b58543d3427d10fc5dcd2005cfe2f72fc3b8663d239339717d5c699ad16cec12cbfb2e617f43846f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2a052543169cf37fbc0cd0ac74292e998c32556137d16bf5e254cd1b34872d0042a5759f586c286a0b2316eaef7a4a0dcdf9982645e2b393f2d141b2dea18d8c5e08bc0a49d8b9d71e735b60b088f177932d51ce8613b16921c6639b33627705d360cbbeaf0d107314;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd2e60bcd212e8337e0dc27b6bd998e6f81becba7902a6394c2d6ca244c15a0a3fc297508df2d37ecfcb40c36530f59a111a723addd2e107e33c0666ae7230dc226ea1d6a9d237618d1afd41c909eecf25d6e0e57190a99df49a81eb67a68f756037e25dc861a09d3ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a1c757019f406e56fb4fae5827742e099f32ced157a127d3c4d990e614a0da88b0fa562d2dd8aec8d4fbe508b9fcd47c119f03b9ac8bb22c30d2a9a9f449247f34a2a17dc59e0eea70b9434a0d1e9a18fa1e26fbd4d8aa5d061f48f048b8589471617f6fcb41b5115;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba5c7fb05c0955666caa763a8a9551715442f8cca52eecab53b556ccf091f9e60a7c62bac3f858016d8ed9551ec8599b9469850b327775416932c57e5ff911cf27e4ffb4bdf53d5d631bc80b17a9178a836b7539d2bcf1d540d21b3626c268107df48614c00f5b2614;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed3fb50a440f8637bea53b97472d8c54677b4aaa538d8fd074a4ff0b9a86c9bf2a5aa8eca9333544a9ed751ad4cacdb1998e04459609dad95f333278e820e72f64cc6fba8611c4f9ebccfd961fa707c1faf2155964de2775592e88de9d276e681e47c0c096656ff44d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h190764ddcb483e6433c9e9de1cffce4e8a128fc92550e01143c3659b3f8e89d16b003c86eff53362f3c59f06123464173fbb14335c8a296eed071ad578194d4febdc386dbf6700c1c74c70017fb634d7f6719491ee24d9f82c5577c279b7941f256d023ae0f16966a0f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e844450792390a3e11ff1f904242a5e94c06662bdaa39aec636f7de557abf064e8e756a3262d29a4998ab313407b5aa68eb2983c9465dfdc81dc9adf152e57fafe42a334fdbc98c27060e8a1096a565f700af4657af08344884c602a2e4e1721d71088f4c7199a2e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e2135782cba8199a054db01735b76ecce56d57cae75adbde54a53d18a71863b3890077108bd960b176ec93fe4d5e2e2309cf1a2ac0446c154900136d6dfd079382280e7b006d872f7c2644383f0b1ad42981a97d99227be4d10fd1af4f2d5fba300dd8aea540290f4b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d09c0aa5c6407a25197b7b80fd5c223e7e85cf7cbb7dd9caded645920e7331266a9fffec5371bfbff743e8c993aa0eadc73503ba2bff12b78b36def8827846abbe8f8bf40943f0a3fbdaa0192d0db50ee225b59e644e593bba1ba97dce68fda57d76462ad3a9291da0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf966da5102587abd31e8f5b93962fcf493642b8b0ca478f84e6b25c0300a32f0c0724f44d09bd827c1f95e91babea28eba78e505b91666c51918951872d6372f4e9f7840b98185931dea2897c0064ac50b12e0bd1c805199ffbb2ec4b292667db5ef41d3e837af6755;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da1bb8b3e4c162ce3a6c2d2647d4f7eb06da60f9e30e68100658d0c9f0cf3a6b8fecab65c170881d8db2a96465286017612d2c1de38629179bebb14bdef63c823014f9d65a5346bfc8f1eb0273a9de14d2ee2bec47749954632a942475f99d6421c2c1267fdee8f1fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c966e729fe39adfe85fb40f584a4b3996a0255e73e727d08af8deca53604fcef7a72b687d46fa547a9f45bcfb92ceda0e443ac7f7a29e7d91b36e8448ee0e52194b9c2eba5e87e34c6843c2737d5a65ccb91f6f1fad30d19ae03751c265c214679889690a8e3f013a4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h543ba807eb89d81211f7709bb063012ec8ac41ca5cad58346eada6f8a70db2da506107b7c5e57c1d031252b670b340acb05e47bfb71881d5d18c77e2a5cc1575361b4669ee2cf33b5b58a02c5f44cc78ba84a39e28cc3fb2c7f32403c7f68d750b97564d28537b03dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142cf7d43d393d06b6d5fee0a7e833796e0482c7a58dae6748e6239e9d5b1c33e1b397ca06d3385aebad29b2e591661dbfdad752cd33018350457c26c1863c16a2fd11a7c0592f1e6010c8aaf40355a1a6143b4718648f92700ed44958a619449df92ad090b0c7997ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h119cfaa2c1eb8b3af96a92a6cdd117b311c0e76ebe312f28e6faf05123d2105d6246919e45b6a316d12091528bb22808b952f9a7a843e829114df5fb4538393ff9aa4cc941d4721e971e2a0f8b401875e65d8e9568fdf10244677e38aaab724acb876bfbc51811be969;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c25933867700412d26e3ba695b2c47e3a302084eb4d97c8a05a100880ac53b2b34de3cdb2a05728c97586560c6a0ac57a18270c2232e9edeadaa02035682b575f014f959f51f1e4c9be29bb936d53d597b1c19ab38bc9c1f62749672c5959b03a87b6e86613a09ae8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12aed19d63039c31a4b567c11c8449d72d082accd3d9ef866ce9f37d5763a5c965f8a1af9818f359ac59833dc4bd76d53f07464406e6c352c267154acd48eec4a76be8489d946d94d36438d1206799b1dd70e68338e9563bfe97fca4bb91254dccbf74bf5a137eb3623;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c4000a87c23719bdc3855ef9be174e48b70ab73714a2f897056178d27bec238cf60bbf12f3065bc2f9b3a989f39e054de99b748cb273325e2621f9d78720265db55c9980d2b23bea3e53a449d4b7cfaf5a2ba630d73c8dc434ce9bb6ac5268d6f7ce58029ecd182ab7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed3d7c2b93965120737dfdaa9a9402000ae56cb2b9d3f9e7f064892a981f8b070a64ee999755a92a5c8d49fdd39138c18308e5792004411016c88cbc68c2f88353f111b4418d4a3916c77840e0d95c5d8617e123868a323b9e41377ce53b9b1ad3cba6cc9b5c8b5a00;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155c956bb1894a16711b655eb26ebc9ecb3be1f4f8682bbfc9bf7fd5684f2eabed940b1dd3867d6cc43445442488b7e643524eb05a31a8e24439a48b26b0e492381d64aa9b377977b6905492275edd44a2cc90a0549bba6ceea3c9dffb5f35a5bfe1ea93ca3d348f7d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8212b70db5a6c9a96a6104d7749329abebd6baecaff939032df4355d1ae1bc524061183f014a3b3a02ae112b9dcefd63d7a1dbd693de06567b2f21dd072a9fd9092ae60eb2fe379dc68f2b85ae6c69cb6886ef35d966ec29211704518cf158bd94d51b23f4a78af94b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1342ffd87f4189aed3c0753cd8c29b4dbf0a50b9ca519b40840255cb300bd3910f4762dafe12a37b3fb15ecb8f49cd2f4ac13f56c59a711c9450f49783f15f1321cae9f3897686df069b2134fb25e7141ac8df4905d75aefab77517a8544206fdf4d5cd6abdb3c98567;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he4f5e51a6f99bfc52871e685fd156ccf05c3602b65b6d94b377820ad5bdff11573d685e0ed4b151a03d119c580867d4df28d729bd3aafd134820eb0ea33df35009967321ab8f0d52a0ae99d48ab2126c23892222e42d9d543dfa9d2423c6e6da10b77e90e1f503ab95;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b48b2e73f911f538b25d5804b0df62939754ccbcde23efdcd42c6208d94f94d0e8f84dd2e46165b3610b383c179c9c9398e386e3954642da19ec4993333ae320174da7120ca0ec9102ddaac10f44e0e3aeb38a9aff500e992872039e991dac30e1dcba2499f036303;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d456a5288d8a4b39c589b699de43c6fb1bc076a6aaffdb834c09c12b9418cc32153e208729b0bf4fcf4da9bd070ea0160fcc661a7dca615a18808ff3ee5a10c81b3d0880de5768dbd32723a75374535802774fce736762f40b28381d5de626b4162722dc9ecfd794f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1586a8894979c36d5f1998d9751a21797ab71903cd2298101fc82f2ed38d7f345af6951e97a0834789f92e2838e171c2fb7326149f8968a6d555b0390ccbf24f010cd7d45bd776127c657a8a7188cc98bcb78742cd3bf8d03fe4c31269f08cdfa43e113bdc5e8182357;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d9f0c0030b86c3b024f7ee15545f9f11d7f7cde6f9c895c807436197e847d37219cd7bae09d96a209f072d12d623104c438775916c639c47d2b3cf90947cb58b892aafec9cc12f7cab77d6c0260eba03e39ded5f41851ae9a678d7ce2eabf4ae6b89dadac262f9ee0f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf05b400e89ae4eecae510afb2959d103f036fbcbd0ad205c494857ee78045d664c7c6d3c39aba552388dc3c5947273caa42e045394bb57017c5dc5e2178c47f33f5d7281e5fdad918ce12f82c7f00861531e9a44286fce58abff1c99b2f51aa2e0c8fb89721fbcdfcc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db916c94eda1035398be92dec71fc7911e7d01bbbc6708632cea8e28d5a45b834dc26cf53271b451c681e7099f62bae9c86a3bae13bb5a2870eb46cf81125b2f9184b8fea402d32c0e3a74d6c749124a48074ac9688732de12a88823a30690b81f350621f2cb1fdca8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122eeab55013b2d2760409a5e7096fd301d6c8410f911398b1637062f38c82cdb9e49adca2fe4d5565205fcd2e94664981b97b063d25316eaedd6299aec407a1f44f8ca2449c9b4721f7c0ae5cf00fdfc6625442e8ddb19ec864da95f391034f557561fae48d826bbab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63292930ec6f35dfb3c6a955b46ff3a90f4a126a2abd0b75d8cbf168da599054ebe8ea062ccf7dcc10304d1c38c05c19b02a799103ddd8ded0b7b5858334a6bbd1c5ee8bc9d23e569cc41d3bdca075a6ba4959a31d4801a03848adfe0f6f3bad5ee997e559d94fc7b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0c692dd4c17c88687054f6bf3093f3473ea68f6807cfff077145ddd33e10985957a271f3687c5798a3d1dce135d7c4d134bad0e38138b0b6719b46d57ff8561e00e3dc4e79025f971402c96a8e533baf45850c49ea2377c72e02742fd8c1741a943a99dbb82e03f3a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e6217e339069d1aeae5ad330d70800f01099369e16d25d814ae91b034c1da5d6a639931ef10b3a9eb404409fd5df087c9da5175887c1766a84ab4de07bd4fc6325c74c5766a99fc6b7722b55be0db117f59ef1e3afbd4799588b9acd31400024fd54a56780c229b76;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h630bbdf3c55f07ef2a8744b011698a6c7b1746cb1e8156d08d2408e8918a643034e6fb7706319c9ff61d4767300b866e3b5194d048a678e3e389241ce940b6431b70b0508172b015257fdf2a4d3f024a88d4a9fa5736ac7cbf439409bdd4b00efd5b47c62ee5fe6111;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h562ad284f252142debfa0b7f5f09a26c3f80fcd8ca2705dbaf160187ccd26623957289a819fce7cda7dd6da4138bdf2ef14c86dd20d7c8357277de414c88e2a3ff79e5c97e0deafc8a1ce41e5103de6cedd6466ccc616e8b672934e751c97cad7e8721365ea15e31f7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h286fd88c4b0004f0d01036f476e68101a478144f71b5d8761992e046629ced641ea29c68708fdd48a095b5b3a2dc7d92ca61bef7d5aa2bf696e7127c3d69cc26fd79d139c2bcc7fbdc6556aa8aefe12a5c49170a2f048eec0c6977d9f2a23f3224e1c32af093c51035;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfdee1c414819b3577c17cb2b54d47df0278fa761c03640b56cabeeceaecbc30e129a19f4f4ea205c22d41f3a269ab8befad65d901fc49c0054b5fe4f8c36d8cafe79c26b3ce500d629f467b01fe16eaa363f64b727d76391667d759a248a879a071234627d1506306;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125064c850fbf24a20da21a2fd27fcd49c73f4a5ae04b70c1f3213caf66b14727d466ee9d4433fe50810b5171828c08715959b347e501cd2576d60ffd31eee84370de6c2725e1a185cebce7ef10d0de5bfb070e1fb923b73b7443453ab7d91de9f4b680e1d4bf156580;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13fe803dfc503ecc0f48a93a61603cb0c7301cf931235d2f9c108beb048a6b5e0c78cd2fcca052555516850d552980fda4e6b178b9cd162c35212446f74ead90b7c7a8c3a65c2225a11849ecff83cd397b58f116c11f8eb0792db80132d06abde17ce543b5f8a197834;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25bdb5387370d050ff6b0e3e482d4d75f090b7dceb8cc512438600e49da0fd452da37be08a22737b8ad10683537a4532ebd62f10d3292f4dc93240277053f53eb8fee9487e6adbfc782045ebc3d4ebe5a13f151d14be05dc3bda36fda8fdda7c54ebc3c78cd7b66d7c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c787caa06343a24a4dfcb3fd751446d2bb5ad42d88e50d54dfd87dd906ed7d54be341a9b0ec24c0eb27e40164f429cf662ace0e6de9f4cdb7e1b1d95627646a8de6bcd2405127ef5cd444878289b73fbc51e88215e63552a831200044c8d7c4cbbd1fa7a0062bebf58;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d96a61a2da89f542df34b77c3421b56d4c82cf46ec13161e8cdf1a8d093bdd724370f5341e9ce61cd076aff1d5acbeaa5a17bc2dfe741f399c27e836acffe47857cf614e9efe520085447ab9c30cec5e42ef6532b05353f6f994fb340cf043b506d48060f78f8cab87;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16335c49381e7b42077105ad4ff59506ef2d872985705fed94637b13f42b0350dbc6a7605c923ec69213a73219dd5d6aab6f9ac239b896e4cea46fad4b99a1ae83942dc7b4cc3069af8020d65f6036d983a7a38f4c97886631d8636cff1455116a0adeb26aaf774f09e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9193fbabeb5962be8e960b1d77bdbd2a0bf8da2b9f82871ee427bf88757f5e030794d978a47bf810f289ef8f81a2c44c1584ac5ebaec1d0567d0e6ed93a4ba91044f3e21fc75e120eaa3820093ff1434050e932c7ba29d6f0536bc65c4a10e925a965efdeff6151420;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2eb144fb8b71be9781fc2c33371f37656e56073e2cbb881b7b4af0759a703e3ccea4d6047ed99de006bda91db606cffc048a428930c02bb29a8c5a55e13bfa520e9f37d41ef06f242c0fd73b293a53dc0ab473cb39a12b7f1c97f82dd9e748ff6e25c5071787772455;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9d5a1b5fc9155a959d2d0cc7f66b231e6fd2b4e3da86d7d93ad2c02d2a29854775599f70e4f3695562b457d2099b6b1790fac8b55e212aae3b63d1b24eaa963eafaf0430f19bd40ec258a8a7eab135fa127cbebe13d83849194e5b8d64025ca5d031e7855cc2271f27;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h644e7e4fdb517aa1caba65665e44c984f4daeaba99b4b2ca406ead782ccc4016eb32378f3d88be0f1d26e9d0079530c01079a69320c1d08c1732e1df42cc931853ca2d43b502172456c4bcb4e387a390272439e89a43c1a80b47f17371e4fc77fda64cf0205e2eb81c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h783f47a4cc8e26fb7ac1c501b1888b548279cbac1fe7370e9c77428f111ff70c9ea131c3b013ac2a6a2e42b442ac07d0e4ca893cc77844c9dbac340b5a9400196b85fb39430741b2c931734ba027f9b7a538bb6cee3cf76a8fcf4cb784b1aad5969968993622ccfd5f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h185fa3ae042bfe924b37a8f1330080273a935aa93a7d8922e66442ef2ee163a2e4e9af8a152bd9d0195e461e846ba2fa24adbe5148936503c424e864a9cf64ac9a6271cf76e8cb97fe57f24f49f077b24e44a5586445b8a99bac20fc8b5ede7f7b4d40c09eca4fa4ab1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174b4aa15d6ccc9bf7c6a681261f4680bc0d6d3c16b9487a8af1d00622235b0257415229dd1279ae63c2675ea86764332f88dbf38131bee8b0881a470459cb657b8ecd6fdf7881fc66bc28be0194ed5ee526cad9fac68a1c21d688369f4860f6f629cc3b8c6e7c4fde9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdf4f3858ab63890812be3031917bdb04beb9ac5dcf6c521c36d864d2c87f504da2de59c64bbe2ac20db5f2c18b4f49af489037b984117f436d5039294d46c8aa31947471b80b7c9e3fa7cea9e6a29097d43d2cb099c02771125639c9e0e7b31797e44d7d2cbc9a80b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h645aaa78a3303090bc55c344e1ec5db09b05949aca678e18e477912af94b90024087bd01ec3970de18498b777615dbb0694c48ad9a9c56e942ec183f51606efa7f30d8621bca00e15e399d5b10bd63b10b661f3d84ac015afbf729be62074a11502d4e29a10d812a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h143e63b939155bf691a9b34b73ac4cb3304a93f20bde87dd10268098078835670d649a32eda0b01159483e3a234af7dd9758fda09edbb06dbae39850efc2308b43e1636327be2f6891b75f0e7d4e3deb240071ef5cdac4744a44fad7c14f6371bf4e62d4fe751f5255c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e9845b72aaac7ba5e774e53121d1caaecab37e75c709cec26ab207d25bb86f3cfb949693baa4fb378c741005ac03df9ea8126423c4f4086a3e8d76afc34a1fc0988878fbc36f5aa4d6a07306e0ec743a8708406d95acdd44282149429a4eea90de6c8f320f0fce573;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b25f9dce4ac9a3045f4efac4c239a73ef6b1ec0fa56830d309b86f363dafa9f482551c072ca72abaa696f62a27ed64ef002759658285dad04951b10e08ff4d934167adbcd38d90b5f6eee53c313c6f2965285853186046ea7fa707be7d8f7d9675e03bb61f45c07aa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h154e0b8a58f3944e05847605e3c68f0511768e40ac86104135d9fd65cdebca07e2f65d9584a0220f399e67f92a0f49decec35f86a9f1f0fa41bd19fca7cbeac4f7ee7932dc3c391e4c94f716cdd2ee7a65e2450488355fe85ea1d33c06c5876e063120d51a7b8d468da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4eebf10ae0d8590ba14d0b5a1893a826e8ed7e3d99db97d563cf698f4420580992ed4b7afc481d4b3666e9b0f87d9c61f9c453865228c1eef1769438be2a8b434176ea7390ce85b2cf3c08de19ac3dbb264f25e565778c273048e0f764d535683571973fe0fdcfbcbc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2e8af20617fa873e8905a310f55152f79e8b60ab8dd8028ae12693dc2989b1ec7efbe4f788f19a6370018d1c1cdc747ebd9efe0a028775a84b9086b7407b59b2b627e88da072eeeeaf309505006ac607fd6e31f600360574c45c35981468998d7f9bbf08ce1565883;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c809e8447fafc4cda0549c395b880fde4d8c72f1676ad5a1069cbc18b0e256db14761483846f8f891ac465264ec52d195b0c3bad8a93042a73165f9d772f3e0ed42b3f6e96e821a1b3a5f76cdd62e073f6ec50d2579bf421da68da9f25289d724767272dd02bdaa6fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h52e1a51463c24be213baa5147dfb654fffd8388b73ce231306b3ed4e762e7f98febb400ca4814d30c5ea72c47be98e42db137203391540ebf32ce9221bc5652530dd7abe6b0d49f382d80ddbf1a5ff545ce6fa6a7e879c18157c827f0796d43773e48d38c64b579463;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e07695718260a7e11fac54416a0690e3d5ff6dcf2c8837770d27a67b8d44027effbbf2da651f40e2bc96af77c8a2fa7a76924a8cf1be5ddc7fcaf5018a394a7826689148afa229213914302a939784db99fb9e22dccb737e3c660241e7edb9ab8704e7a1acdd98ac1c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hccff7ecb7f0263c887e4a0d1ce737b16877debd54ed79caaed8ee616ccb3921c2886acd642aab51d0333dbd33de722a76b0e1608465a90c4283536842ad89d3c0dcc72b2f1a76b2c10f199e14dcb56e3d7b0b73f842e9c547667ef9ff08e822707a86798d147414898;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14c62a66ae194b5e33473ec2dcf5649f716ac4ed60edfc6561021d7e47f5382062d12f56046d1d187fd8d7381ac12ef968d12b3ee39e56b091b103026ad3fc4ff328d43e63e4e84b0420096d3795a328c8df6b86c0143c5bfc693bf43a717c83db55dd09a34e4be8f44;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5bad4d6af68440054ff8d9897ec1dbeaaa68178943b4d9f3698a0c9e0e5f6f48a5bdef29f956ae8cf04f0aa0e1f36fe1705338fb401aaedcc20e7beab73e465b8c6bc24c94ae06aaa9d803805fb58aa6630b3c8d4216711b745312128c65369bca6caff6a1b67078d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb32f2d62b3c500e119f5a9172bb84e9fb0799f4bf8441bc44b48ef5d137d76ff6b26b1046ca63885d88cb4d8faa8101ae3e349520cc5185152e1f03fb293abbf3b2c6f4b11435c679abf1d72cb3de474cf73c6491f0d847e58bd9cba99244d4ee20bb2717c4d07f55;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ce7f094c8ff840bd740649e733b8dbb59e360e6ced3f1cc8288587b8d0bf836e34ad1afbfd9f7dd27bd082ac8f22a539efd243cc34e4abfb9c22c75728c931beb8d43b5f0f7d33a7460e729abfd0c9b3c633b8fda28aed6c51f0fa596e8554391a48215c21d8de5670;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16ca87bb33e8e5eb229093d122afc1757c79c8ffc89d3cbd81c57eb61ccdb82fdad2d3e296ea52ea7a077703e2510140108a9fe5bff8c78c32e839f479323ba39fde7f782ea6d90df0cc8f9d732e17ebb90fb1a8d95a831204180217926265a832c3c672760ead1fe3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haf3d327d2ded962d8180630ccf49fd312aaf52d289d032bd60218e48a69a2bf16ecd07cae762ad64767134bb5a80b560ecb17aafbbfca9ccd896e052761d642a7690835ce1a50d60696d269a3f85ac5bac906f72968f9ff1f09bc8296aef0ec6f0ba653e2b13f6ba82;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc7b1609c491f80bcb6a653ee3ca502f4810336212e87e28c85100f3a1cde8f78d05e62c62670172b6bf03f579021bdfc2ed85134f6a7d86909c0b7c9d5297973560e51b9f9eb66d10d4d5ddfc3f8c00c459cde45fbcd9917d80e62e9d1113661569d5e3d91c09f580;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfd7632c018c6923da88326f469bb618bf9a111e491bb1f65f1630db7de037ac3a27839a55ae142876c4de0ab888f68ce261150167a0b05d19f3213ff619396add7f01cae33289dea98f727f5a0a333fdf1325166c54bdb72f8a66731eb8909aeb57d6a66831870a53f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123fae65bd4fe7a7864499f356bc1979f81cb7eae9b839dea85898b865c18899491e9f3fd300cb64e75ed30cdce5b51400e25ea6386b5a6c96b752df933344266139a7064b9c5b43b0f9a23ebdd448dee2c0f6606c248fad3038f1727cce03fe0e9469365898f427192;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43083f1ab35a867668d743ebc2868e9c8bebc2998b6969deb9abf1108159d8ea81f4d2898c27b740f9faa2d79a911699fad876e48400fb70369a8dd9920fbb35d162330bd548f4809b06e8483f4ba71a520698169693d0f0f9d88c9ba7fbfc1b696cc61531caad7bd6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e036eb70795842721387e50b929952c6e121d3e2155bbedfc7e37e8d8a680f9aed5b0ba1841ee2e999da44a6c2417fc89fd7a405d261f8afc8771fa05933ec3c1edb3060c16b0865609ae61b3ad0575433d7680f0fa336f90283cea14d81b68390625eb48e1351ce1f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b9a14e4311e4e901f53555e8b5321ab3797d1cc124f05f8dcc0d936531a192c2d2761afeac644f44edcfa4afda0bd628891e68c69215577e712392f1e6be529cc13a32c21c3209547e4f805bc6d710054f9124008772e6373002c8f0dd835bcdd2812900c29ffb759e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18fee28253d829f7c01bc2276b0d1ce307f4ef9d913778a63105e5eaf1583174cbea746b80bc184f0539127e3e41dbec0dbc6e281dc672d2422e62c3b216bf1e843f1feac3833939524d674333acedc6552faf94d53c1a2f28ba669ce3835dd0df4abfb4bb2f70dc373;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a6d496b26b80a2f2b1e6ff4ba265c049196f27d948683f732bafde90b89e45eb35dd5f088f1362b7b800ea7a150ee2fb41b900743a4a6f243d404822e8eb9093636505dd928d3708ac82dd95efaab26ef236791af94595e8289d3871b78b03a561bd2e61abe0471ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19dc9553d62d39d0e1a1ec3d7c5aaa9e2f279bd7b5c52534783ab7c0e734dae61740a9869ee9db6973e838b712682c304fd6f353e98df76dfdad30ea06a832273c6f89c65e63a56ffd12bd51fc17c8614e1041e2e17aeb76b08b5a66b108ec01c689e939a89f25b4ccf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1004baa80fc1a2830ab87c6f208102430a56d49478913e5888a1d23023c5cfeb62e85911954f42ea613b0447c3fde7509e7a9d6604f46aa564c88b5e9a7ecc16f96566288389f17f32d1579318d9cf76670d6eb68222e8997d13af5ef4e2d254574247a64b7ab1c73;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h127f5e7175f38d3877eb29faa615589e9ae81e075eec5185c2d5da78d05b2f861121cba6a12967cad9be8b3f6378df29b10ecfd2d92bf04edacc2e75a0532ed00f0febfb3741e33dd75eb08390f3bd9a4ff83ad796b38d82fb055642f5807a980e77765042fd64cb339;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed94e508d9399039d6692095406eb25c2cc5c5ce64b151dc0fae209c16eb41e35e2efa963beecd7ad15bc49e999350f0f0ed2b985725d4dadbee4654d19bc2fa269d3768fe017e55404f512c5d39dbad005542a9c99ca3069495e610e0846e753c6353df87d07e206e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16d2f26261481d468a678859d35268b8d5119ede44cd1258d8ef2edceeb7b6e5d8e809b3a9fa1ef15d6956be4997ecf6a70ceb8ab031677eb70dd7667bd7f3c73934b802d61df61fa6297fc8b825129975906af9ac8712e50404a91c21abe87da4b5c3aa8da54db1ff0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h181f7db7d8095dc84c372fb71ec54bf9b385e9526792dfe44585bce0baeda17a94d588d85169292bd3b43e0089d4739fee6f892ef465b0502ec83c03dabab73ce1b9c9b319d58ebd27dff8934e3be5f96f7982e4e7d6def717d8fc79970edcc857c34e3cbb468ff835a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1315c386e400b40a591ec50ff110dcd41e4620c3d65dd7ea84f5c3660ed659573f1bdb0f18bfedf62cc6e88a3e7732946874601b5a15d244cb212cb56dc7e46b831c5e6d83476ab6c7c32b3ddfd0f543f2129d0a752b92f7025f604a6ffc9f1f5b6fe8e1c3e293b49;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdfa01a7d40acac6ad33b00415337a0d20bc591a168f7a8a473a1aef7bb8d6fb4a71c774d0040295085768049c1f6709a14e633cab8f3b8290dacffcfa9b874eda805520fed5d6f13b2b458e8e4dda506e2f9c6408fc83ada60648437f3ff8b1e82220a35361c4bcc76;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h39cbd2e12a069271c0b7c9dc48f8e3daf05098e6172c0aec8e6591d013aee4f46a49022eaaf8bc1c05fc6896d4a0c2cb24c39fbd86e59c22a46abfe53c1aa1b7f296c54f89d96e0a26b97752f3aa47dab4075819ac118b6f03595a94e47c9f44a8829adae69a567a56;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he598c6860206b6dd2836adfd0259dc1e2f426fa2fa317a77b1a3bca98f0d56f1316c3ad1f386c224ab84a466420f4a2d22659aee1ef7f5600a5ab0f4edc2949669b1a47d870c5a6f3b54ca663e2b63f1d8bbbb8ac350690cfb4720aee2bbfe8f84e4b6299a524806cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a0720c95c8dfac8b585276281300809cd66dabb135cc22a9f36f632cfe2e64a1adccf355ae3242f7dee1a41c6fdce1639c115aedbc0f0871a3ccf8ec0d8f33d1e6330b7903bc7811f39051522bc524357c96616a944f168f53099408763a7b1dcb09f42aadc94b8641;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a6fef2a26cb9aa19dc1a04bec3d28b77668866af949649db85d32ca6dfa631b3bdb2417ed73cfd13f0c1dff239432babd89933a4e73fc62bcf7f027f1c36552afc8bb6d07f84d42a33d8e20eb15d3c8d0a90b06420586f7ddf30f7351479855784eba6487951dc33e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95d7e9f9238f32367f561570d552136ddf2e7b03f52335e6c77bbe035117dbaabcad1f307c1e82c95094d80de6542cdc3e38d7006a5b49308f4de986ba1a439c8c5050e9b2b1161b635b5dd4326863e4708c25eb6e9dec05359212cef08c22175fd9eaf61c745d36c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1020e6a7df59e8334c4ea3a314b22c2c5c2c2ec188d01367feb74523dce75a8cefbe65c343896a174acd18e9f54ab26891bac34a943b6f8b4e6e76e069f6e6c75623db0eb1acbf47e28c56e6c9cd740aa7f86697a4ea6ac94ca8dfdbb84061d09971e653ae5306c9d23;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he5fd3988e458e931f4ef22f4f723f223c4afee6c7cad7158a53111d1a14a9f9bf36e453363374270ab9e329871498ebdf289dd4b80a67c3998baea9bf0f1b6f2c6a394ca740708430d44e3c1ecd4483dc408559f7218b716106e8934fbb1a523361cc50785b498182f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h91949a65b5da83c7c74b2a60ccf8b0aa889693815add33805080fa0b0df34388bd8998da3606ade8453500961578b3824cd310959af8d830e069ed7d931ddbdf6657e98cc02e9433a9eaaf798b41d30c5a0b52dd4752c4f34bc03e534d8aa316d06f6c19d354e05317;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h942a8deb4e4b6f3f3b3d0d70c8386e4715d91acf31e954c58eb60306e44622c2c339ff6b45a3c6083f46d257b74c8d9341796b24659c5749418301f79a8e5a3f170dca6a4e0ba901b1bda799ffddaacb077f77afd83c5c1acf5f5ea1843847f02f999fdad00f5def39;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7df19f37a8498a3360e1b3cf42eac0e071d1f7551ecc57eb468f62e04b8f01160bd9a4f2756806b1367384e95760fbbb260316e2bc96ea25762c9072b77c80724f9376cbebbe9c3d56af53a6b723b57b08e77e05a218bb6b6359cfa28420ff729f9a1f1b915e46639;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1503fd09aae3e08dbc0f98f5d17ce946746608dce11c08941c51185a594693bd9009120ab78f106e66cbbeca32800184823e49ccf56d1726fb63bd3d1f4c62fa644444c884e25282f288fe980470b62fcae8f339d094110f48bfab8497ec3f714e63cde176b14c72d44;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4919d83b6f93ac04cf2470e943be3444339bd453879fb725cd4b2002aaa2b97b0f2b11093a9016e775016cc29df8ba81cdaa9ca0b8cfb70271cc030e5c7fb6258d0bf894d74892655f9c951be70ebfc9b604733b22b56a0007d04199e9201fc1794f44fe6150151c80;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf6673745b3abc784328caad419cdbb5fb6529297819f5ccfb10529ef252b2157c6a347996228c5a8d6d25e35f25fe9f3869be7b82d2fd945b5f20dc12a069d68d970755cf8d210339f88f1421624bb6d358076e95e8ab5ce7f539b0d511217fc7f14217c677f9d5e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h30802adff051e4635f5df71e02ab8d965ce00e432530e1d1b9830bcf0978c37297e6e1e235420fd3efdfd3a88a29d26fe2d3cbf61cd7e243f1aad73fc8b9752382cf096eb3bdd1a1c5cb2044a2c2223c99a476b0ce80e2237f7ead7f145aaff4a33fa36736cdf32ef8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b3f0d0f7e4c5428ffb22a5d0709fef0cafa88580dc68d418780f58ca4eaa3a3901a5bb60b2f508c301033ef927727aaa96e901d11d5ffd25a07e6b7ef5bb2d092845bf175ca20f7ad34d36ceef5fd64a5b25b6f9a05c7e81b929358ffe1afb43073fd5658b96a8da8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd8dda98d443b4aa5e5083a84ec2470b265d0da8a51f9e000bbafabcb2e399acb4f6aa44f1c95bc6603e3f67a0543996a86632755ed6cd69ab43e86f8198555c2abbb0d595ce3d3ada7f7fef8cdb4c8771cb1fbb6c99ccd1390092f7bc801695491c0faa9c01debb0a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12fa816ea4dfc51f3a65e4a7f41068f489db6ea4ec1c8e9979d0728a3f6d8b7f40d7873fc96b15705330151c4aae41eef033e3dc9032fb03428f373fa2719240d081c12d474c2933e2db86509f98636ebc6c57cb5fae6d722504a8e380e7838fd238afac9ba12ed68d0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdcca6bbd79b84e9ebd75fcc0ec84da09ae5a867ccfec4b08072345709516c6e91c424271a0793f5e3a4f22ff8d191f9dbe61715ff3baae8c0422f02b53ead6d1d6c0ed2651e1c6c8c0a9880814f6a38e6a33c916f5f6346630d82a0d8c11fa620e7de8c9f33954ab25;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1830925278bb30ce267f9b95279a491c4f2b39bd6d2f983f552f1b9fa47d7b084630d9de8aadf1e495d79e2916b20fee4c8057a6e121f614f771e996ac937634d70515a65a4c5d0688d2951afc6e512cd0561cf5ccbf3357d910abd39759dfc1a52151281e5a5dafefc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d47390b922269706701b0f33589118adf921a1ef0c0ecb2f649204d18931cd740437e9d8ef30133c30c4f1c7c1f3ab9e9022810ac2a2089e7dfff1afd50e331bcf687d8cebe92b230348dc4013dbc8efe7ddd91277aceed4556eea52c293ebbafafc3a68967ca1e150;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ade6ce778fb41ad5053abab5cff47ef17cd75bb0a72e6b46c2b1262b55a974c82450c5322243f323da5a216bd7890c3b899b005546e9a00e49a7d62d47d403eeebeeb2daa23e88c0cfdfa6810dbc988f19b4a6d00eccd34bcc47eaef1b27a5340646634409eb3b3da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4f1ab957233073bd28f48d80d16c2e1cfdeb367b5a23eb8ed17b27523dceeaf113ee5ab1bd4cfa3f3a70c08502f44188ce1ed1bb1d4dc61efb716991b7735b705abfa968416912e08e0c26f712cc799ec4a880cc24478d59241e198147b6034bd2fe7e09e2c6f8fb7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16321c6897f088a34582ce7a79975cad6a7d6676969406a479ff6e908239bed5018098907898f45766f0be0fa7633c81f116d743207952a708cfccd7facd8c29f2745377447ef04c74cdd15c218137d4b2f83de8d87a1f7ca015c707437ec7b6b9f142a223ed77be4c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1268f55caf4e56b2405ae11fc39a9a61f449d41951c24899b95b109bdf1e174b04bb7638f646b57cd8d0e20f00e993a3d80e832464f8c6152d00eeffc927094ff374d116ab3a3b4fa3c854e1a14722b9b86f89ccaa0ec1cc5bd8d8b8f68afac1d5d56ed65ec14cff145;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4470fca3f817c836e523598e587a600d2814fea1c851de266911c3549f56d558db91e671d03e2a6490f83f294a9bcf9c57762081a881e0b20b4640390b569d5807cefc10ee7f755c3450e7840889659b9235515b7e96190ffea0033c18e8e42dab4f54bb24066d9fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbfe22a8f9bee70fd8a36224a273cf5d5d6885bdae1605d86624d7e1afd39193f687b2f3459094ca7c0e18991c911b947a1e5c968e89f42f1ff47e62496948b71c4eba0c1ad2867f1438c5f536c4a517a8063f198dfcfafa7ceb863e7f1afbe04c918850d4939b0b346;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he89be03a3708e60b1ee58f7b32f86635707d9c68cc11f37e953866cbb6177423c50011f3f84dfd70f9f9a1546635e9db1eae51e2c174eda07fa7e30d1e4e9bd8baa6c5c3680495ea046e86ea76ea09ca60b4bf7efe73b4d4cd10bfd8762f18660815d997475874f0f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e376786763aec003c5c4e98490abd40862aaa2531529f9d36ace26d9a6fd79ef28fad4cd9ea6ab7a336dae1f703e14573e91d99b7f3aa991bb005df06563934e63bd3346ed87e455b5f2d5358ff7e9e9a6eeaf6453317c7b795eae376c0eb27c393cf74fed2f2f267;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175251cf0e4472ee10c8c11f3ddb8dcfc74e2d86d4e2c1faa2410d5c1da9c8b0612baa412572ccb52a5503f81f66b9e4b310200fc8719e3b8cf00c78f2e1c78d9481ddce2ed527575ea5c39b9394f14933fcca7fd26d0775cdba47206e2b26d7f7c0e1d2ebe85a044dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1216319c04cb3f174ac09c999248fc9a8c549df13fd139845b4ea097ed27b959de52c7847e2ec394e8c604f76ce41a8e089feaf412986833f02c7224d81c33a49f84d6bf378dbf15ed118f674414f48ea094ef2323c8f28fa105a5d7ebf52a0d488188b79aa8f1d1a47;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he7132b10bbe2438fb003c864f01952820d086baacce208a15230b14e0cfa31346b2d5c0cdae543e8928d30680634443729eedaed97c38aeb914781df93e8dfae9007fc250b25122c0a060df5753355e1582f6858c410b6f3ab672b6c6c0b7841a5c6599710d3dd53b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2de8b73168382fceb85326bcc2b84e2712fdbc5fa23d78e1a7f3337a942d1d1444174a3e372eae38566d9fadb2b87b1aba6548d6f8c13f51a78e0b425ed9c794bfe61abc375167146ff19c356bc816702179171e14ab9924b849cca82a872e18feb804ed65d0dc7cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hda1129b6a3f4e6a6bf6301b2d6aa43b3037cc681ac5d777c200aff640a50d9594d6d1c7bd781602e12dc913164f91b4432f18d04f9faa9d40e8fa6ec96413d77a799b65e479c0b17fcd04a0b0213526848a0fc8d8a99d3bf337796eb2536092b2456116ed97b68592f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c2c9f12c2f026a9ef15d339fcd307e17ef8a71f37b0271945274fd3b02ecfa64f029e9de4d13ac7ad443f1fb1238324d27e568c760586647419072c44b22dd9ba848d8d4d81a6ca66dbb5b2184c1fdc66a6ea02bc502aa961b3fa25ad3c10c0c466643e5716921f631;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12dab9afed67ecf2ccb07c430b52f972b7f6ec1567af22bc857f75e01e61f9ef68f7c5260593d360d290ca360c642413372814b73ba9e12b4e7a73b70bbc471e477ed58517507db44c977f09bbbf2a0d5c129666aa7a179deab449139f0651ce9593be1c1dc6632e5e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a01e7c94faecd0d03108518d0f2217f22961b473e603fcd03121349e9f9cee20cb526308b33c2e07e05c3f768f30def9fe19bb775b410081129c1eb5320ca993f80dc24ce1063abfc9971983bd686fdd04b6b8584e76347d667f3e04d52c9fea96e002f8a2fd5593a1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h47f38859b4f9827626765ab584c4af59d90d4835d0014b95c73bf274f96ba200b6f654cca7d71bc06c1e29fcb10e7104e2a2bba55b0d42862ff10a9da56ab4774a303aeeb3edc56352eab1b443b44737c1b8de112dcfb025af08041b59f2083e95e3bbb9f65bfdccfb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c42bb487bbf698ae0f87dbccb480873b312dc5bccdabe447edfa078630365ec1eab2b4833694a38e2110c178a645ed5483cb2294e52c54d9650527eb1ca86ac1300112a73d58de0ada6824e90b8b3e6ae238c9dc19764d6acf58cebde5d9ff5b435bc59940a7dfee80;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h403aa936611fb3f9316faef7a1bd683f9e6ed8218e919af830571796c8afe4bb82db4986fb80f1901efd5d805295fedc229b89c1ae0920fa3898727dca147151a188e29c76e10bc6ffbdb25ddf77605e2d324dbd74f213ab2d7be46d73e3d575778fd05557dfcb0eaa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f6204b678854ed7b76888d88d72024043818cebba788ca3204ecf076e5876193207c067efefd604cbd65c010b1c4ea3ddb1e9841c9a2570dff35daa42500b8b2a58c4ee064a731e3cedd7e08ad096063e2b57723e994168e4ecbe4796c22324e6b0b07e1c82e7c35f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5aa61b027df34d700a518700826a0f195b797ceaf8ee8ba55931fa0ce55228fc1033691d4aa524eea06fdb61452acb5910b697311463721d9c8a09bfe60ef124b83d7d75e62e417d04251694c78b3a569b486ba21206206353bc1329ea64e6ac2119f784cab02256f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haf42db11f85ba10fc8f1837b7f76c7fe553d9dd03e35ea924fb341a9f6e9d643a3a377b9d5edb8324b8282a96debade852f8c6546b7cd9dfb4751d1d7d4939d7f10056df26168a8693024c0808fb4de31e4717e6ca01e1a0c33cf9683b4b48188b6df8f3ba4bb2e2ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a695294aec29dcd2b1be9e62291063828509b7564937850577d8337e74567d888f6efef4bfa9ebf4bb934b4a74e4e2016adcba583a6e9071b77478741ea2426caa2bc3fb3c30d219c2f725a35cf1d4e4c665f4b85796ddbb7668ec523baf3af0eb724015a5b6e4b01d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d1b83efe54902b8571f90b6ba76ee3de3504bf07cdce137d6530475de86e31937c4258bb83c3c5ebe4fdbe63883eac72f4f4cb739dcf6c72e267d605225280648ab1c7624bd2112b21c184fee127362c2ebd6cfc4023ecfb7927d24af437f7b924baa8662da89d9e53;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1603e7f88d9d00e1fa7bfeb9c09e9bb2e891bc08fbbbca244736eaa379751c2c2b582ba9d8d868e6cf7ca8117567a19a2b302cffd5058d420753a87f5669059b1ac370743df6bb37c8b818be10ad99b30017533e9e0eb537e135905129b2db6955d5c398c7c8ef65fdd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb35bba7bbf7cb1905399641f7b3f73394987121b2e354f444c3b172c8825b1ec346a62ae316b7fa207a8114190138acb69c62616f16dcce63a58e0d6e16557fec42b2258a2d7b7802e370f7166c2fa1ecb593a9683040e250206d913333e52b81dd5d3b4253d36f84f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb923b5d63e1c3f2b07e18ec72a38a22482a59362bc187c01c8538376c9af547d799c34e26d8f1bb73035435e35969b559af1c84b5c690953f56365b36f43b549e12bd6a8c5436e328ae0d748beec7391c0e7d99f29a8b37465b3ed687d9d9c3164bbaf2f4deb90a46d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h181c880c8b8f6087a082d5c1e1631ade58fb53d6b635a8456634daf60582395870e54f04b32e2113667d33714ed923f1b52c582500091dc4dd27ed3d79b0270cd75afd51fa0d62628559e729f9f8e2de844843aff1f4edb13c815a24caa1989b6eff442476633115a37;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197533534815bf4f260620cb018cbf2d8277a7f7ccd67311497a9c13e706590cf0cc7d1a11a17ea507f1b06feb9f610a76b9c93484d12dfa34c1d53ee1b2d57bd10c72dbd55f42b3f6d4eb24cfee28bc1de3876d36483fc88775f32f3d96955877650b13aad4101e4a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c5b5e66758a96ea603ddea3984859d67f77b71f10b858e1d2af6efa728361482784598fc701c11a8a1ec90d3df9961a0f73954c1a996a683da5c5aa7493d6907264a63d5410c6e9b0b40cdcc6d6c423331eeee05487a5c1226923afc9f37d774f5adff707818fe163;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcec7ab9614940a656a2b1bbf4775ad364e967967fcf98cff9c978ee13437e1fabe1f0cd8682d8ef79827e9a0b5226b702327272926ded72b8a71f07e49ae55286dcae053e5b6c77f246108c7274f8f353a2b12c5e7788dd8769e9f19aec820e41253e33b1c89ecbb7c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h35dee89be55ba0a194d7c9c13debef54bc88ca7244e020dba69420c3ee413acb4be14cf412d27aa63e33ffd786806774e1eed5a448fa610015108abbe26bdd30221f003f700af802528aaaa1587bc7adc0c483b473a28e01169926b11b2d252a594d894a5b238d8582;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11f9cd32037ac421d2d9f3c52a1cb28afb2588b82d4ba9f6f2173e448ddbabdf92a8f61ce1bacdcf17edb8f22dec5e1dd62318ab13e08b5218379d7efa57d02c59bb8286b0a31a5fce026518b1d1a6eab7f85c2fda80910d97919d6d30909b76aee9e7dc13db2abfdda;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18f75edd069ed12cc6970fa0b82cfa85eb3452240c99fd9f9609ab5943ce4d2582dcd2fbe67d374b9019fa4d3e650bda2962cb100b2324ea1bf9ecee714859654a1165106d96227e0a5a5159ef744c7c9a90e7a0749f7ba99059b04505d26843536502afa73b33fcaea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ef38f5ee94e2fc6f31d332dce7ed7e46785e4df56be143a60e7a925df65c351c54a688d4bec151c90884c5b93a82a049e6713201b37f9e72c8b86cd44019bd6face6d8235c5b564043a6808a621ad42b96590b7043d4446d47af98c4184e68c0e2688cbe95ecbcb3e9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197f4973dcc435ec469ed12203cd1759f9b4c504ceebaecb0a70cd684840614bf52c0e853c1d103435f65117f4df47571e2e4d6b940be2114702fc4b725eb9f5c086c00dea51877b9465c07f3a6c2a5fc852fab14c3b3ba23dc03db70c95282d8e7ab3f6a6fb40d0e44;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h157c5225cc7e01982739704cb738d28279dc6d42f2cc27f71716ee9c1bf0067901bfe3682eddbbdff0ee3df979b33049776ad32d6677c01890078175cc613f5b1dc21e9a8a42723cbc278c41a6b8173d261cbbde0adaed00baacc04bd8a3987f535611cbc542f8741e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h160a9bbd26c0df0b66693735cb8bad0697dd0b15749dcf7c8319595320a8cd4200f62db4d15c1e5ecbccdc8085215d07f9277365b3ea2b2c57845cfa65f8d3507bc793eb888006154227a34815669b51eb50503fd7cb364ebaa218098595b364762d205ac9ccbd5feeb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h986d1e08e9cdefa3763519ca7fe2d90745783977dd72cf4c25377575cc3275e5a738cfbb009d2c5ead001d30e15b4d84bf4d7dd8b957a68feb6e433c3cbb271360f90ad34b2a13eb32ec1093e9fc64e2f48df16d503dcbd1de7bd647643a475a20f506fb7822b54fee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ea11ecbff7380a540af4e62c2120e975354cceb6c27b0c6eb911a2d49e5ecd5ea98b560b43f997e555c748af7fedd90c8a58a807276740e5fd0943b7797b2138a8ef41aeee2ada43202043104622308ccd8725de1c1d26af0dffd511d69d4cdddf4a0b39f0f72a9259;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ee93cc3dd3408c6623f7f2dc5b96f9db85b44883e470e9d1df366ccd0c5b58427a85d78e901c8b03a3f5a65fa1a0195dbf9bb2254a5c409852c001dd3b8026faa69025fa1a1924fddd815aa3327e236acc66125e09fc3960199e8487f7f43831c60227f73b626654e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd8069fdc1e471288ef0d83a0af7fbd9f9609fd053e8cd7e85a93108d21c11cb5df1636532f7f279650a74698e44378326dd9cc31409b34a9f2ee4b6cd6cea69bd12a4d50961ea86a1164a8288395aa93a9aa0df4debf8d173c776ba6a7fa3bc52a0cadd5071dba93c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdeb0c0bf8a98b0ce1fe427d69f3bafa3b9a0d9670333961e73c11dd15cd9075f833f5598d9ef60f34202fbf055c3f558d9b46a18a69438fb7caf6ace24527f63db66b11cf07e8c0882d772fdb47d252399beecf92c83a31ff3c7a872407c6f0e2b8601c487eb6353ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1818a649873ebc24f849a3586b96b5454cd6cb11829c24540058d04d96fc3ec3b84b7459c48ef50570d7dcbda9c27669be7afed76d64e8cf54b1e922d2da0983b5dfcfad53a6b89b6666318f3fd45d9edeb923cce4227edaf01877526cda2d569bfc0e1e663de84db5e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h80b2fc3b28654e38b8da5b14082938d20e60fdd4daec0b6d70915a10095cf33a4c2176910d2dd347c17feb8a56a99934f5dfe0f359581656cb4aad76db23787f30c2ed6f66208eb7cf58c0c632f8df2545e8054acb39f3001df19fb5a0e2455bed136f9ebafd3da25a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heb59c2a396acd12f55a4f9becd105b97948a6d3556480baaf5ad3b5b26829ae3da1e306c50eb3517ab49c803080b9125cb0685c9f9576f1d0dc12455944c9ff03dc32d5d1f9bd000198b7e200565298739edbdfd0b70d078d7c7c6fc5b44e3d49da5db6cdf32f09c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15370e74ae40b2ace4ee17b94e62ed845d9d877880ab1a0c52b4c1b7d7b47143e191142aea3f7ad853c8b766bc5f98f7ada8271e7df726aea7dc55ee7bc08335a04f8dac66a989dd65f6ae7bfbb2d06fbda0715c3d67cb2465287870d91a3a9c97a9da10773f7142ccd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h97f4790efe94572e75b91d10ac92f37982a171b628f45bda201d0a422e6257996122565bde1a01d27d6ce92e6405d53d3b2400df06c47e5a6b4cb04fe794f4cbefe6fea33f742785f013ba1f5a772a5adf40c596ea39b771a6de3420e8b2a0ba67e47a7a33f436036e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he6b6cbece100f8bb139132b342f05f1323abc4749e2b48fec92c4f43857cf8fefa65b91f342724bfc41c544e29cfe63a71692fef2abfbd9ef659db9b294031fa9a3a73b89339df657b5e95c2bece0712507692d3f8512a060134dce51e9b6ab64ee7633e3c39dac720;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1486d0095fd6541afc424438bc7f1947d43f0b453bb72853919f45ea72aeb55482c6ee2bcbb73cd6acf1f16a92782019bd2ea819f8e96acc0ee813e501a187ae10814c991ebc9b15cd05131b5d220016456779ad705d29752bde42429a980b6c077357a8ab527ab95df;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h839897d33c9f0d1a5d6ee8688499e766c6991414f7e981b8d79e91bdbbeba7338c3790535299d2f500aaa12b5389bb6a442c1ca38839d992840f06ad1fc832fb37699db36091235816b7df93f789d448bce6546033d34dc36c6532e8bee03420bec226c5d14d2c89e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2bc5e0ddbafa3a8ec30f2db94ec7271303f0a8ab3103af731ad07f0f9bbb1da4cc15b0cc9e404ee2e6ac9767922492111f6201cd4b517752e697dfbbbd8540d55ec105c07bb9538edc1a842398a75d9e0919c06e7849ec8cb84b164f34bcfe7a3638947c38c91beae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h85514af0c8b12a5351d3c09a2ec1f09e1543a824d44821dc95c6b463d2c94ad0eca664688d219dccf041d9d9773d20e4a16399be67b082448007bc6f55310eb3968b1c30e445999b5baf441372a9e96b90afb6411b4a1099e0edb6357a2683554b5db42ac059db10c7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h55362462a3e8019c07acdd29699c9c8fd790f60863d4afdc83a286a569c3b72428c33ac6fad5616dba05a29bce00a42d6a5078268ef85f650afb2c985548e8264918877d052269ed5ae8ea08c3770148b34cf142d7b18431b5ab89b1bea65449b5aa54017d8156dedc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc1014a187045251e453c0a956cc31d9d94e42db5a9b96d267470fa764e3ca4c90fb568acd26f4012dcc1640e6896ab0164f7cedbd6c2c4075b980e36a2fd849cff98331adfab49b6e5bc6c1d004e20084a13588d4a6e4e2148e2d2e2e85468cfb46ef1ffcf8d88fa83;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c6cc474589a9edd3566cb0a8014e3095e9cc45ea2ff3c8de3daf0b15567216f20185e1a8765d4d0ad701ded09b69bb9919d99aa4b0933d84f14282e2ed35d744ec10e037d0dad41d0a2bca0d027182368c7988ec34b050b073fc2fd121e4f6514531a12003fd80653;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h157f1516fdee302f860762b118ec9f21df80c8d6b0b11995e694fd3ae64bbab16edbbca664031f0243ebd814611b03cffdf13c46f7f96883638e50dc81283be2cbc7e78d3f21d1e80ed2bcd8846abfcefc3671694748f98e613ea639d7e914f1b7773c4e3a261ae7179;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1925da4fec192c220bf1b46598e465ece849c1ec73bbadced066916c4ca4a0354475ecadbf6d5b79624e3451068868d7feec57f7af143a8194ab23df15ace003627d4889a374f7e3ad24d01e378a5464eef6efee06408a053b096f1ef9e2c0877e5e4fbbec134a04a7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4815d3d94bbc24b88e99b1b72d8de887f76619b8f085a12cfd53ca7c372e37b4c1ee6418ca4cd7f556b2b3829035928b22018185fd3e34f63ed1e45372bbe06cc243e73409d9a6a508a78b73baf1a5262080ee5452dcfc84ee0c0824a8b58bd58a1af5f4ef1acbbba8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12b9dc5f775236e4f439d26df626e6a2bdd32bb8121913fef3ab75c31f2933971658ce240a199507fe49785a5ba6922295b54f0a3ea6de4a98a1179eb44ceef9126a72fe032ebbadb22ac311b2dd165ee2c1e8e88b5e06969c4940d47cd8501bd753fa9c80971911759;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12e6fe8a37e448477c5fe9dc3a3b292c5e4ee40ea5a2973e65b103cd9d1c7dddbc3e6db6b62436555087b1b7372659bf4ac96ba87aaafe4b0f20d59095693fdf642010df50bfe75e3d5e6807ebe606697695c9be74736b588a3e9ae928f4c9b10a6163d2d0d2d66037d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb2642ba6f40a3874239ef554350bbbc5a5b66d75366097476b470a12bdad9c5c43297cf69fe91687f47656ac090675cb049ad706ccb1d25a377d1fa8c798e564a23f96fabcc70ebdc5756e5d86471a5118edff6011e39f991868470ddaac31054422423cf67cc89c03;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44e8dcf2fb9cd3dbb7eabb1f95361c894fa1d237590af116b2b8262b3ce3ae6fd3f912d080c4778b44710045f7f30dff2aef608540fcb2b7e8fb337c11f957d718793a243f800b2ff3d6ce4fb08738970d3f8e7d52a7c1de76fde0aec26f8df568b4d3536681e870e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4dd1b18dd34bbe035ac6677461e567ff93ba9b10cc83cd3fabe719570b8ff0a8472ded737e0e70fecc260753f7469ecd104afd985a4c1bad00c63f08675de39578a8aefdbf32a8952e5cfdb38ceccd6b8c2067596c0ae7bc82e928c7cbe82067f47d28c5eeacfa5892;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hef04304fa5d6b57b140921b0f4c709d4aee8acd207fb2173c0288cb2622f1fc619b6eb82f74506ad83961e3c1383e46610d17948f7e0ab807cf1e40e060903da9478af71ddd5d61631b749e4b6f749c1b60ee4a31542ef45b9f85f1d33e16a1bab5f8b8f047afc74cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha8a88073d750f24faf33b841864e8945e538b482ca4a4bb9960b5821ad7f098dc3369da2488d35d328f10733da530b8553c35da59ada58f2f98e551a0a0f1c81dc35c9cc094f7b49ed3662c74ead633f7be161a863033a8903ddd70d01fd1298e28398c549d4027440;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd9b8ebdf8ee879edb6a1fc007530e9869aa718b354a4aac3e41b88d56ade2374c7e37cada26b7c1cd463c87b19d2c311939f81e5bbf57fb45b6bc98f35802b3130a29a06a0b8e0641e91cc5b713f645d1bb65f6b266c853a93b3791d660837d7cdbd148855ed3f15da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96fc0e58947ef1d5f5442cc58835100000fe5307b1bec6cf694673a58d5fcc0dab869257e84db575cc72ee9e72c799ce79ec69decdc9c2b7bf4b2af12efb36a5c2ec4c6ce99fe1939634b360412ed0d162bf4c6d8c0d0d98d9cf9755841d896ffc5bc4bc7967110ca3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dd9488d8a765ebf84546a583838dbfd7a52afdecd6d76dc351dede8dade2f39ccf0cf81a5d1c02c7741638aae4f535f3e815bd08fedeefb4fc05036a3824b923b31057f7cc54d85d9ba9260ac1aa1135131263a46f7231ec77a8e230cd0deff69701fcc7eda349c16;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a2a06bcc527844cd1b6bd058740f745bca17b2d0b69d32b323bef0839cf940704b6405810db8081551939b2b426518710ba8ce562385769a6b39b3b3167f0d9c695f744cb28d29da534389e994329f58ab60a1c08b51752dc0e7d78f51625a0f8a90cb1e01c6f64f21;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9adcd65cb368b063be2bad11477fe138178ea6f508613a100a6f7fd7ecdc3e313e591542a2480fac7de521aaaf3736a66aaedae41fbbc0cc3bcbd25dcb1316ec05d2bfe6d5601ca5eae3a554db0008d4bfe6d53976572e162f16c0fde1e5f34409b6dd982b055e0947;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c0ea6e5efc617be2c9fb460057ef60876d55aff552354e71e8acba247ab0dcc4c27df2f6649b485d442d63e5a97abbb39156534317d007d56a513fdd1368633b5c6676a851fbce26d339038f38a1a1a54f8394add08681ee68fbdad6a0714703f37007efe379fd4a74;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hacc66c43f8ea78b31bf3cd7b2efedd7be661d15982bf608f305a3f304b133faf2c93becd9c72f1fd730ad1ad2c0ce1f088187b15e21244c1c954aec69ef34dfb5e3cfe0b1028b3198076f4ab0a8876f735f7e6e6cfb1bfea6d01877abbf5185e8519923621013b12f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfa4ed7ec2a537b7c2aa1fc454be4d352de73d22f95867ff15de28914bc6bd08dc4047a12fbba5091baafdb398983c4de0a48662867aab61c2ad2888943741bf680c3c3c8b0da9d08da836717333fa9b700252794af2e8755ded913f64430f21f62ec3cf4384850247e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197e1b49ac9ca513f2929dee353bf588679c58bbf0a0e4b8b603512b63ee59cfc70c61cf29952b9a33cc079bbb7d06da26bd044abb2e960de21f440f61febaea4ce7c597082e8135090e4cc927352404711a04d6fa0822d869e532ec6a9cb62f2d0b60d4ab6dda6cde1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1002dd18c9c5bd44c9578855cc6e1902da70470e228f28014bc27df8f8965ccc71feb7550b17f5fa25d58df056a6df6b393b9d7102328c842aae074102d67f54529577e21044aae1a794b2b02757cbf4f27d43949aae0468737920287874a43885221543497c1bf3560;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a38870c862af9f29802e6454d7c216c98362402f9bab84d78f531e1d44a4893d0d01aa04fcf6965a1240bc4ef4d10f71c153c049c40de50853e849cfb20b0ec97af352fa719188e66a64f09eeb41c7f0fc4784a915005715fc8563efc04e3df9f676321bd7cd228fce;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf86619df793a944d1c67f3789e46e8d777d519d60236b28f9422896e724e0ffbb6ad4e5ee9d7ed02e3cde0b53b19df1d2394916434916e1cc49daf23f3cf101293d2f86457bc2df40a450317ea9387a84039b0025a0fd3bb292f2eb184ad5f6a84c4dc96dcc543f0c9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14184c2a56234a7494a26e97e12f6d8b20fa39c678725275bd11d983768a1a4f158137d24a6d5b60571b29a38a1b8272bb0cbf59ca0f27b586be6653bf47c8a7d0bc7fdc265520ae5e4b3105ffb240dc54e3e0a1ee40ab7b1760cf3e1d2e587280a078d160f8b7a63f1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfd03353b82043cd843bac38e967e89e0d68b57ba962df99512f962881a09cfb472e011ebc9f0fd771a6f8a8545eae4a602186d802fb910559da65c5daa47c9e61f0225eb5a9afe15b452e230bc14cfff53d0e5865009aef1fd4962d4951ff37703581622802e9ff66b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af58c0b838ab7f24f1030102ffef10fcf94a435eca7d23b0d705cff3f7acac21fe46e01a0d542616a247197ae7a117bbe1a58aa7fcc81520b518889342839dba8f64bd9dd8bace3583cbd5df665eeaf3bd16f1462b0bf3b8364625f74e0c9ae9aecb53c254007e9f2c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14684f74bf80824b2fc4eebfc0b87f58f3f231f6a40fe5b4e81ac456f7e8f371af90c24121f52c906e2e9afd26f516ac927f0b315ef5b5d33ec4c04afaa1999af09f4a778f33b36768d02a3757822ab1066e3e3e2a606fced59a13d3cea6063887d0eafe0b386684dde;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4de20181f0bf0e545cd69b4b91b4da2bdc7d2b68188a9552f456a78b183da7506a4d29ad655b47b7307575b95849c79d6d89145aa340f51b06b0e651136b271867dde4ad0a0f7b01f2b84aa6d7015937a7d1554b66c73f0b3d6ce9cd40cffa82cdeab4bcb1f681b1a8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h31a6514c5a7a1b6d640bcfce1bc5d44999ea049818897211b00997d6132e49154e3059e834285c68f7cad854fb1fe0c6580c578b681fedaac095a492c952778224a8b001bb01b8a644623e8de263d8c9d85124bd19ad47ac662988034ed03508d63c4ed8a6417abeee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h132a96eb148a587878220618143a171d737b609ee60684c2f78607394ce1a6581bf1cfc6581194c152cd868ec2cd32eab593ef094f750186ff48a81bfe9f04faa3122bfa19c7f08a76523a3a9a36d3aacdb3101d55cc90b27b2459903906af84519354b15815d154aa8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h102d7060e37d8d0c70a1bfce0e2b58b07350d1d7db991ad3463f49cbbf4612e7a0108ad5eb6849d506e5a05d8fd40dae3f3bbe574fadb3996f3e0f58b90eea1abaebbb88c78d40893cfbef7a55ebdc7d2bb18463956b663997d3888a9ae11a439efb74c355a15a99cb2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c4e8e49d7a386b8aed5b3cdc22ae0df1267d3b5599889727f9febcd2403d25de0c0399e5b175f02d5422a955b557c7221f6abb01758403bb408a948bb35e50df01d7dbf34694b5793a02e9f4dc0a262a28d52fc37029f9b3da29fbc3cc48c9ee8811fc34366ccf0833;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hceb05ed0cf0ead2cb9c3503d4d8b59d86ab980eaf81118f68b2ffbfb89895bbdfe9d5885992344792bd51b56f92ad01a1734c942ec870c465449a159a5ac2a067552a5c403f7bbb53ebbe5e8e62d827a9e1701273bc84d4586d50cd4000de8f52c8a156fd45be0606f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8d9d8bd1d92ec9b73dd1720cc16329cd8ac35d3a5cf5fc88380acddd6df22591587cf6c53c7a7da587a3b814b83112a2a483bb516f75753d85258f6cac5eed6bc64304c96db7d9dbe76e7d08437d62bd94d1fc2524eed44b1d92c8d4c714973cdac517da210cf8879b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e39cdf16c8b010f307af79728a82a4f913e6f0175e6e7606f0f111daf9c1db47f275e67c76a72674653e7bb4ffea124c18e8709799d26483f4c7afea67d339a87220955da295a418558237e2770fc2a56f5be59e24edf562a93d9b32668a912ea94400e857762a500;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177e850450127e94d8a9306552bf2e562f435ee4d20e0f111d70bb41125ce21eeaff44445603f2bf1289d47a3679200075ed4eb95263c158100b36a7ac1c504f7d39111835af169bd7ec14d94a383121fc61a4e4930108b38ef5e736faa6020574b2aacf1cf7a7f02f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1205bf175a11217d51ace52ae194beffcf5fbc0f8ae8a3f34ea2ace11907ed976332ae1f7b61ddbeac5a345a7efe1420d384276ce8c269ccc8cb48d0ae27ee7d49b03db25dc471d52d8bdfc34346bc2893f5cc5b1cb26fe485cfc05a430a7a7cf0d4de3df7467308dc6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f8245e7a2077c992127db8c89f8059f217e02d5caafa801bb055b9bff215065bd77bf1827d98c0266e24a5d6b00543551cfb0895d57710d2f71851a11600f875d03fd6136575526d80b2acfb8920b5b7d92db071aaa3edcdd74742e094ebae623f18bdb5d72078924;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hacd4d222a24e1faba13df16d649358bf1447f36eaac9591a61a286fe4fe5e538dfdd488b19f16db0e80a90ecce4216e8898aedd8950716a3e9d44808490528131a6a9516a08ecb2e4666426a57d11ff797f94b694875e73dff8bf7176ec7c22d41116e1abea8b483c7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8310766d3b449ead92197c443690acb33e51ba7b580332277bc4a67794121e2cf67c90eda9394428ca7160e8a8beabd008b1cfc351fd2be76b2570534e2be60a3bd4441bb6c4b3a7d94ac159f96462096d67d52266bce0368aa618b3d2dc110823866b6d3a0f45e35;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h81e607cbd29fc39ba8b056471f26fd18cf4d12e6c42a3892e1cb9877c1b218452fe3d85102387f96896b511569f455190b8185dc8e075b6eb1c6f6e12edeeb978219047ff1bde6e4e5234757f9822e6c13ce3633af7b633531c5989c45659918b37845b5614debe091;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197a145a8eeda1eb8054a99cd7c87a74e8823615d3b8be595924e1e79ef0cd483b89a12eeb43b413ee3b7b2d4038875c638a0b3016bfbf72ea59ac69c8895f4cdb0f9c18e7b9959a7ed46cc29c0b97d55ec4d231e9120bb5cf4855d7f003e757753bcc57675302e18eb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11908ae48588e28c670eb2e689e4801b46d8ea0c73f081e865a3a3c96c89390a6030aa07a7d8849cea4c834496a2276a0c1902e3ae1f32656d069acb650507c669eae9087f93bf25901fb737f47c886c893466a5a417e25a610874ebb500e331ac957ad5bf5529651ad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd7435012473c45246720560b32850da78f4868a9327a8786553e1bf1c445bf72d0be2f92a0d4cc0ddbb995289387650fb5411336228d0be194e83f37fdf22ffd637198979dbc4af31c8b872256d153f9cbdb82f1f4fe325dbb92d5b983d24392a72e46be86c7ed1246;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cd720130ed73c0cc2e1f982f1755d9f5d763de748f82387e21f5ba25ada5e6a5fa20c6c347d43ad57fa72fb512162a781f94f06c081029bcb5fd76f67e9a8ccffae9d562a72ce690ca65293e6ff474247f5340bd466346cfc51a997a222265c495b56eac00e312e3dc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18767dcbe2dfa2ad6e7ff2cf634d9bdfd6f8d5ee1ceeac7636e80f1c8c6ca40c9126c436bbdb9dcf251212f2fd31aff4320a75df3324e2cf084542c5f5f222534328ccbbd9b002122cf3c113c992226aef79e18242c4cad2e518137b4067d33a020491df95daa0d21bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb893d213d3eff0bd24a7a1a08e972ff4be39da92d7754fe4f0791331a57156571551af52ef0ef08492a7b937a5ff88fe559530ef669520a8bfb067419d6bfde7e537d9e004e377bb1f370bfec6926c3fbe38eee18d52f2b7a3fdff65235062984e8cac6efcafdc225;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1997e5402989f26fdc5a5bfee9bb1a7dcd5d188e106cd94b683902ebd31654af344ab2db57e2d8e5b607a3586fce7afa336559bc19160b86c510b3da274722753ae6ea4f92946b759988fcb0a00d704fb008dc6d482bd8693a55b6d5135654294a2e53933961a585035;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b47c8dcb650667a54fd5be8a09267fee89a2d6c606f778126c7a20abd513fb2d1f962cdc03211a72c1d4e07af66080070067015835b4f399c6db534738ba96e4378a860ee831a387bdfa7488448d249e3096e5bd5c25167141d030daf0f899b6b426b24d87f7c4a2b9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h984942b3cbe142a206720ffc2cc66d77875c3169d69668ce2c05fcd16a1d3f9feb6d02d95d2d23fe2cbdf86882cfeec1509ce91e224961ffa28781bf23351323600fe67f1389d1acf425a096e11afb0e16cfa70611d93ccaaab204380bbb012f37b33ba68c4abd6e36;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2bb3d643b2293e5c9190bb89eb6c1f658abe0459d12cb8eae6462a684f3a8cbe44992d06d37b4844255ae81ae0b4becf34ce2ca98ce957cac51960fb42ae2049325254ba0d4ea27bc3d47c72a5b74cb32ce1b3a4936df3dba6fb338182a3f5c9841b44af6466b8df9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdd10a12d6a4a3787cfbc0afd64318ec62eddc0fa80ec85bb78a21bef0a8ad8441015c7263c5a40baa13bcf17a947156d70b820af244120be61c8f0e23f572e2f0e9074d3a857181af1377c6754aeda0baed9a53576cfe0d4671fc9b0faee014e60f703a8e0a22a6404;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h386b67704a4fa07c77a1730b977d3858bda0846476828d37534431faea81662ddeb7fa2c4c5d888aca28e4c188212a7aa08a1c8524d74e230e0323d1994333a821396b7100d267e08b1118c74b146ffb93515e442881e2860153da3d46d928a3346ecd243fe7a7f618;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2898a1f51e3b5ef39d2081df5b7a9627274f0ccc31301740a2fedcc02eed7adf78f64d0c8752e276a14c61ef5de2a589fbfdf80614edc938c9fad97c8a18453c3fd16b10ac33b4523f63d5fd593321d14e479af33c56eac661ef39d10b64b00f43942c21290a223cda;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf58aded1e1c77a00e2dc5f33a817c78d321037d32bae73cfdde4acd6a1e4e1e8725f90881855f8bfdd6ca3971e33d82704f00751f09251276bf32b64964f02e1cf6fb47ec701260b4bc425b4d39192b2cbb76c85b6e5effff97244c7c4c337b78fd6c4f30c63fb30d4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17791e34d96d4c19eed2fc7e0005974accde73c5d9e8b21c25154941bbdcd45848d49de119eb474ccbb3fb7b67e8d66de51e7058cba8a2c5b0ca2dd54f11fba2f3dde33873b0d4d24b2fff8034951187dc3f7dae5d3e2341231f8463d462f38f74a53f64b0876a04042;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1515f4f4057e62333a74aac73d071dedbe717c70dc6494147dcd2fb8164932479639eb194fb5eef324bb62c3678dd6f1beb878e2db29246daf0d8756aa51a84e4da8c64998a54ab01872e60ef934ac391f7717a6456dd4cbb519ac58000ef50b9dfb5a6f3c3fcc195d2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f01d488f656a749cfa7221df8d4916d70bb90465320e4cb435ac254c0ae450006feae37a1bdab88835982cb00cd81a49e8d82452854255f15486dbbd979a3854ebd1202f14aea6d9b8d7565a207cad136bddf5657196a0c7a6970e78e1416e5f74119297bae8c9e0dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36af00055da6beb3f5470631b7221195c8894194a5602b8bc7e9d0ad176d841b01e37ff04e638e37453967c06967d19cd21c37cdcc008b4d3a1c406b1005c5c4b69a82e8957757c96876e1ba080e5a4cd62fbb5cd569871f19be533a83c430b8a5a0474bba75926c6c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4d5862357eeb39e80afde6b7f259067e107c61c0bb50b4bf96bf19ccab1e056480ef23dbb0bf006573c89c8f3cb7793ac296aba84f89582906c00bb027fdd43100b1e37bdb96afe85d6edbca0df16014c971538a74636de01b6a93402e60a5e376689fc4ca7c018dfc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h97b026ea6583a813187d4fcb17bbd35574ea3b888be00fd081eb9ed69fed42e312f58096d63fe939c32bfd15c6092e0b00eecc95ee1b375be9c795bd9d50f53ef5b45fcf85a9d660d4c3663f257462fd2af29f77aaca5e52945c8cd53109e545b9473440a2801c6320;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h127680b23038ed88c12111e1fa22260ef1c3223e0fed02f0ef533f97317d0e3b8f772db8592e255cef41cf89bc238c2f07fb5770d924d2e28fc9ee7914cc0b86b1e209ba03fcad9477c582f61e9d19a7a3b68fe770310c5b24e104851209905dffb2a02cb89e9cfd0ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15e9b9bec1c6d58480ab341b74a648c414a9a66d35fbc50d3936b4d3037ae4117c1ee1ecea27ce423fa84cae67e835234c0bd6b16da20365676e79051cedee3c17924e00af17ee0139fa54fdf68cf41dfcbcd4eb6639d5a2650c8648101fb931a3dc931d94a672924f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5724d52387beb12c4a4b7b6c0936d105ca522ba858707db966e80dd3490a7b880e8ced697e1c29a2c35eda817cedecf6dc8ff641990a564ab4d28ea59a7b3a401f5f828e0fd83cd921d65008e3d09f65a1b21cb64eca491a424ad0f8a82c107382a4f582a1ce31ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbfe2e9818288611ff280c462acc60307e78b6975007b408d30d8094a16bd5681d2f2e5df5b9ba5ed4aed5b9b329b80518548d93bc160982dbe390aac1e04f58d348c9ea232be796f0dbdac69c4cea5169ccf02a675436a689ed084a965ef41a98afd4f049259f4dfb0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d4d7ebc69f8e527f190943cd53913b99fb8f79b8019a74c897c42ac34e5192b1a159e6d9c68f96fb45308f5821c1387a48cada85a0189d102314e47755cc2a177e87e9a8069daf61de2301f5e6d5b9935a568246d5c44e865b1ca9a3345c1a697b2c741227bb618f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h309734c6e8f331d22c575bd3495a5f5ae130c4c97e70fac4abe620e7245560c2fac33c8bdf800f6117e73a88544ac417676317d3e47e08b471d8b6cc3e925b7da0bba83f6f8aa5af7e6a3fc00ebd7a5db73cec06bdd282bd0ec2e7490fd5833ffd952646a24850958c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1feb6e64fd22b9ceceda6b0511dcd9bbc0538d09a4bf4e9a452b9e8facafa6337e48e7262b3a56feabbacd75004d60de88a0a6fb62195e0aa4036cea555571a3562cb743c64f34959193a9ab3a850b4801b27e5975ff8a84c9e5a8794cbbc40a9248600bf442c50a557;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12883a6444ebe0f42654d47829b2179415112f8a5f0fde526630092ece52fce52d9e9600e6eda64d5fa266b010a22c6c4fdd9835a78c8920049ee99e54cc13d24a8e8cf36b73aa66048250623a2045205d6be708d277d903223a8d0d74dc71dbacf2297c75150d542d2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150fee107b6a0af4d8ad208b5acb58240b448a18aa1a3d98133d1f170f9c162226cd2fe3b93fcf9dee86059c8b2ebb31674c3270c2f88bc541c6cb9f37b710e8342e57ff3f8483d0acce1058755bc5af10e88e9b153a9476001e95ff9360577b6c8506a05ce555992fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163eaade15e1265c91cd2fbb1937a8731c4c069af1b8c9d917468c585c42fc74a8b41c39e889a06ca664884d6167f3f1a60895e6d8f81f9aad63577beaa3f0e576dc08790f0d437c509f6930e86b60e32a3b1dcad7e9d1edd5bb6b363890c59215feae285546819384;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174ff887bdf070cb2b1f04bcfb8214f6b7399b3a8a5e784710d62fb0457f2516f6209531212fd73ceeb33f94c222d911b37fdc3ee51e5b13f1c6624ee43f5e32ea1896c93bb2ea1552be77cc344a2932253ce3dfc91d22a8ddabd39b63792cdcba955b4908b8b48670c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h84461b07b07322e47d8e1682de7c0c3614bfd2b11273c6bc913ab11cce153055e1b56b3ce78887094d04320180d93239c5c4fd57114d3f21e2b283f61b8e58efac71e1eb7ae627981948a7aa8785d0c34fc0e3fd744c7d9907a0d1bd7383a7ef885c019f5258966a89;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1af484273e5a4cf560a6698c15ebfd46fc83e183178b28786838dda71ab6bfe98d79c6a221b00597e491c91081b8c9b5322a4adfe1573a6739e7255f4e8738543d67deafd769483e565e636fe99785bc704ec3d8c65c360b43085a493877b4be2f85066d2d8478582;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1532af066eb948fe076df433ac36357909c7ae9745875cdd3b2dc98af3e5b64e2e3f5d0d06c21861d3cdbb2a635b2e4a63dc1c836b412c2bf3f0e8fc29013156aa720e10e5a327f6fc326b35a2ff553d7e8ae8f6a9612a475a061f030c91d769196f3d3ef0c1037b603;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ca62c73cb8c12806b3bfa78fb83a93051993a66dba3c841d0508c7995f579b415d516cacc026e762cfd0b5eb53403b9210d9c4e289cfd076b941230a03821279b34e052f08d86db623df314b9bda0a7194b86872e3ebf7693d956733dc97823237e70892f029f9212;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59919c060c774180385e9ee37c134843b9cd803286a52cb01fdfe8590668cddab3316e7ab1e6ba6e8482a7aaf608d398bc6644dd6af91b716619b69113efa5b931cda34a11f44820f3ecdb168fbd02b23c3f8e5705e3b78923d0710700e8597e32fd7d6fd0575154c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha397d76be299b10401266d049da24d0556083e12753c3122c966cf28c8ed995c19f0a5eca5ec8a5c1e820b5118a5b81b8a258fa10f1f388a1b8db96b9269d509fe215300d2cfe0bd75658a3fb7845b0d393b2fd51fe9dda0eace0f63f551862bab697b14b0caa8cfc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bbed6a3eaf9fc024cac68dd867054410d4eb0d36762c790347e4ae25c81cbebf5cbd709f5da8e97e9c59488d35553db6d48f71d8d784a37dd84d05786e9fb38e15008a8297779ac13dc3c3c379a31e8420989948142c77525b7439e55fade53faa90c898885b6952e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha726dce939765b2bc7c3011739e65d7fc4ef4542a1797cc983e2c8bfd57769cba9dd1285b4339a9763f5677c84f62fbb7abc227486f83a57363d25aa3c8ff707ddc007d31702533aba8288251d75420d74dee61cf0b78ea5558fd96ce6cc606526d7bac6fc14cbb440;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d80cf2edfcb3cc5bc9fb2c54bdf56925a79054c08c37ef36ed9cee7c67a5a13671bb362609a0c9f2711f8deddb5d7cc2840715aa2cbd5e789fa426cf686bea5ad30f26e08ded330184ca0c02dbb98ddeb01992df83ba6e1aaab03e9b78ae48e244ae461c014b319222;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1285c3d8867b8ffe83f67866e392ff30e505d0339ee619876d4f027325fe0680344ad9979b24a81aaebe7e8670a0e311f0c3137943666589a156f5e5c84bbeb95914079168bb14355a0305f16d575c19c11763acf5993ab0935c03d23bf237eb0f32f74817abaf22489;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b4db62116e5f8c7211b3fb07f803285f5d942f95ca558f5a5c8097e00a8abfc153c94348933b9bcf324dc6c4e163447b2fad597659f5db3dc2f04a4e7f8d494fb797c45b94170c04676609e05a36cb251ff2a8ed0c13c1a1670fc9cf9d004a3ee123d515018327439;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a0078501be991484b7a2a85d4dfde3a25b41e3e4b39db3240c9d1f1446d895157f1b4b88db54fe5fb68ac9c4383b2788b5bb33562605e74dfdec791843fd4a4469661dc707c11d24bbad55211364febec8d2e531acbb03d767bfd83e622762ef645a27240c966b41;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174a10c4386918d5aca10ccb1fe751b35143f7316e3be2048365928b7dac78dd21445536420247dfc169ad4f3744c5ea0ba98c9e3a544c6858bd7b9de1618da90769b2aa044c4ff20ee9ccd4e90ee4d96470e346ec125f14715e30d675de7d0c5f7d1847f6433a427d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h57ca55602a59289c0a6c06e44b9dd9d1204eab2be2cb2b9169b61de18b5a94fcd34e214b607a35e272f8cf08ab08076a4648ed323cd192e243377627ac5f9c850a50d483ed455d6ae037857c2721b2e3b011b8cae5f815c3f6f22402539683db132797a62bb3ab57ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8d39d2b4e276194d0a05effdb40c775ad272ae111aeeaaa1d321be4aa8d5dd620503336e4a81de73feaf17c2d93e6d819d18fd2c5c9381f4fd87f0ffaa227bcdf8a20c54a8fdc23d10adc5067527710c980719359636e4d1eeedd92442950db10b0528570e2de4faa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd756ac50078f77ff0ff7177390e3dd5bf170637eba63ab31978821f013dbb86e7345a975250feaf3f59f13f839f57d96b8974869835525e0c8bfbe92ebbdee59b496ea9d7941461de7f13d45a20ebc03f9d0402850facdbdbbc532a2ba9ed970eff4ce17dda389770b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha670dc6908685392e9cddcffc48ff07bfa6a292d01a02dd03995aec7fd70a13512d731f36a1cd40724afa13352d75ea9161a38c871b77202fb289536e8093a6ad3299c7c0e204ec30479d3713f623e90aea4dc1e83db74d683b242b73ae692da7ded28973be01ffcdc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e597b645b9855828fddbac443cfc0659019b5cfdbea85cc55fed3aece95d8b7627dc21997b996c7f781908af093c04a4996ac6d83fe7e9511ad6edaf0095a77f7f3ee09089a6de90191b1a95ea1e2e7db71352e0e4b20ecb1f1160346c91e246638a7c5051b0c54a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16d52118f9e19b3dcfc97cb6553206df2679ffba43617132a1a43c0a302d285c55d010d4da4a24c86e8f3c3ae73cc8bc5cbd0865002a0afb113e41d0d59c4e0b00e30ecd248dc8caad170381e4ac57a2eea4cd4f3c25f40004a7fd1ab4e6c75f9adba6bdbe90fa6177f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f3a7d9cd2b163918bef1ebafc9a51d392a1636339ad460cd3c18333b3ce510251d8d3c28fbc15a44df687c3905d5d847d8b6ee5a0a303a1817689aa434790c20ef886e055d4380debe87bd5afd0144a1328de22848f337775de27a2a358f62b2be609795f102f564f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca25cafcfd86c0fec65e8f7f619dea2c1011b57ce901f35e44c8ce96484e2d0f9fdc9214be9613749abba0e523c6d9b8278e77a943e809253907b9fa43acea260f6f88663d258ea6c3f1871f7a1391dbeca8a618f85bd404e5308b13f936d7caa9a1e936585e142601;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14da9a60eb3b79a315fb6435f9ba132510fd63c08441f94822ada730ec439b8b49099b5890b00d3a9244b2eaa710ca1dd230a4c1151d89dd65279c1189d2b7f750a5008d741e2b67dda2607135d1675a4f75c9fa3b728a5cecc7faf8cc3b40c22de6e6f4f21163784ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a627373712244d14d1f00a6ec046172de4e6281ed6c825c0f5f391d7319ffc0f337b841592654f40fd35eb6bc87c5a632ef289e2b59b95bd949ac10ccf7f4df9cefd909331d120620f3ca6f2dd493180181c38f4a1a1002e0f39e3f46810413a8f4a79cfc04c6587f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0836481dcacc6f4f06fc251c6ebd5d5b0c44f7ec18036c207dcef4890836074211b7be99a95a6c81277d2afcac90aa094482e7e995a4b92e744faf7541cd0ef4bb7289c5b1b5c0807f2e2c7ffd3cfaeaecc455780ac5e68003dc96af86afff13f7fe7f745217ea37e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf319d50d6e621ded9a8c0e197e012dec1ee100c1d8c22a05351dacaffb97a92f06ab15192466a91239515f5b301dd6e82b9351585d8a1edfa0fd840b55838b4620be7151b587cf69c0063f12d84f6b73e25ac02c347e792d48004ceea1158ebbc9672cab28f0b18479;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f34ad04a4bf2e03665771224a8d238f700bd396fc3afd98e4b6465c574f4110844051a8333cf489ce185ea253f1dc7d15869d4bd833913c058aa923ad0ef392457853eda6196b643a6603258ae7c0d5ea7446ae48d9074c895631eaeda4fc25d0f54aa7660f203f9a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d6e84d9193ffeabb98601321b98843ab04e12346b554a77b60c2f7ebcb59f91d62a7f3b808496ef91c3e3f683e2f55fecb31a9002ca24f871f625ea829dc8fabcb98d765bf9f10229bbb67b3effbd1ea9e524c2e11bd0d1af666e0e544265af9407c91ceeb83bee95a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd99a5926720b9044c68b6cf6b8752b90b18160be0c109b6b5e9c1d50839c11a71c9e986925eaae4be4ea038c275f10e23179de9856c03deadcb6e41b16fb9ac190dd503834eb5b9edc953de38ba3d352ff2a13cc581a0cbfd277a310a3b66371cb4965d473fe7fc5a7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2938a373875926884a84f935e450f18f8ac556e17b6c73942bf228a99af71858efe640abf9d1031e99a1379deaf121a87330b6c3f58568d0b980b0468e7b73f9db64d3722f4f2d4577467ee3b331491932eaa6c79c68fcfed312e32dd492b2953cf2a5dab4a068cdc7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3f170c9e44d97b82223ca4031f0a7d447bca261b599badf3c82f114b25f987b6496b037d53d26a6f465e024348fcabb805f1a6cde3fda62be6f7675a0c011e9225d2eab2624e7949bd9cbd4a6194c47fd156fc2b084302fedf7654fc098822c17b8d4d75c0fb854e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he6d4d8e63e62bd579ad1409d6019ebee83e510b039e92f35bed6610156ec175ec83c4184fdaebb14c42532b4a597bb600f2917cc6181db45ac41976096422d9e4e7cef24df2c06ebb77f2c3b9670fca4a743db085ca24ac2c1dca7660752c03ca129840629c6d228fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10adbe5a97e310a2d87ee334f0594a9b0446102052a725e5249885638d0e21181fa7a776a2af56959f884d9bb75b81d79e1dba49c508a2c1703bbe73171d9882b18d2112f27ca83725d28224b441c731bc288b746392e20b87f43e40b473392f91d33ca83e6491c0a2b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbb6307cd8cce26b4958952765f6f4e6d91aeecccc2c9945ff5391feac9612af3ec5a68095661f34e1f21b2e2430a8ab74a86bf465dbc2b9d712a07d89c57412b1080f8b60b8560d564356722bf8b2fd31586e92ed04409b28694013c63ff048a42fccc9ce31d4dbb4b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19ed77bea25b78d9708cc86db922e47fbfc8d2df62eac1ae2b5dc01ab7b968cd2aa1c73a1e7f0bc06575392daa8e835bce18774c56f1dea46bb356e746ded60caf23e6abd79fa207debeabc8765c0b9e6bd75449fe8336a396c8aa9dc7adfc3b86d1565d6cc3a3c50ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bcd3486ae7c172fc659990247ccb590f3076a360f7c459105d5ec37977712447a8f1d9d21240ac264a821299db06adec6b483ac7d51d7702cef78e163a3aa07071fe696811a8ef7b9f014b30f32cc95a3a1399dcaf8a1349ee70fa2652209ca22191930d65e234338f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8d5ec24614a5d100d569fd62c7c8604789c161962b028df2fb45b2882af473df79ee965e8fbf78e9f70c271eb81c988fc4c04264dc722f5d4f82e456141f2ed5483ee390385aedb2734f9d91e34a026a5471a624a8f7868259c46fe0bf8f8a575ad267139a6aea6b78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f08d4dbe6bb9abc0e682816b909dc14617731e93fc3bdc7cee7f18a75b01a476f0f29e792eed9abab4df8e79cb4dfa1432c79a69d26cd15d4b811b2aba9c671762ceb65e2060bb31becd519f7c5e25e372b5e20b8b434d42bc4bf101955fa9884190d7ba0fb13f9ed4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1622026696f06dc14e53a766b6c142518355a341a82a6b88928e9c58407547cb726b8a9bcdcb73ebe782f631a448f56e52cd5cebcf4c8cb0f6753dbe48ab8d362b11af4c252b52c23076aea1ea59165c9dede0c0552e321ce755d98934806266a96f9da0f1b522194cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1511e6b2bb765ec32e85cc03e27d984f75b6af6ac51487be4d4154eaa15cea08cc6b366adda16d3c51ba85ff0f295fd242f365af76adbcc7f89b1be545fb498199b555932bf36c77108657746d5cfea5da67c7d83e1abe0e3c16b8586f9702dd8ec7f5ac0a327e768a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142620cecd5f86323a0e4f348d58c9197e3f9841def241f9ccacad39dc2d5b8cacb19962e9887acbfcacd8752bb85c6254fd12b96df6d417b212b665cb007af93f8aff45d60365748acf0894f8ca946c10ec54aada79cb8af2995df3ca6fb34b4e38b2bcabf2c43e6b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h93eaa69ad0ef1c3ca0927163781e0f00ab4ea3363e9af85a4b74eb1f5074a895535499ec24f161ad3b9b7f8baeb3f702231290cee0a2ff930acb725f969405ba3db745aacecdb5d2739a1947dffcb34681d7279ad371337d8e0620635863b6ab95bde94a56c326ea1e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6af886b1d7c2d7c70d505c7b9f87cc083fbb770a7a4dc0e96e3a77773f837aa8b9900de7be7c7091e963587733fdbce21888706a93c8e64dcb4755e22fe4470f3d692909a37f54a46824c739f5fc400420198b0a91c2eff2693f17292de4ba16fdb613583453c66d2c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1b4a2797c2a46a1d8ad9579b228ebdc2b2bd54d4935235bc053803bb79700df111a00a7a3ca5b80b5369c47bcfdc6c082f5410fac98c1d3f446ca26fbd647c5938489cd6b3af14fe4f539c4542ddf46217cf611bfb234c30486d2bdddf5c240baf1fe404ac9918e1b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4b3a023e1bbf599f99cb140d1019260baffc596f222c39654909b4a2ac2cba564ab1d2baa8bb9d56bdfc14164d1813b85781b7f45576c422766ad78a28ace87a3396ce41a057db5bc61a812f387da2d239bd1d979dd76661f7f33cef187ca2085f9960f9eca196ae34;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d185f63dfb01d7b75cb10f6525e46323f5a6cd0c7918ab3378741e1db043166465ae6414678e49d1e9a7fbae42251337ae5ad21b7456158b85cee2b7d50f638fe54b76c7c81ad430eee9df155837b7c4ae902d852f95b81194a34e039e6c56fe5aff7fad669f4235d0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14512452f14cf11aa0662ea5633462e63db149c9a1d98689f00392de5735b5312ab76e6f5e0c6a55014ec990f469681172a9fc39ab975a0f98a715b82a77ea9fdf0fe1bb218abd3ba96017e1ac6f0ad79ecf24686e801c10f436ee45a218f7e6d1201e5c400ea6f9e27;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fa4a0b1720563dd760de852fa1d94d02448e65b02ba6c430fe2d4564d3b0d301b78ba60276d8b52482df4266fdda51dbe06e653c9910b27c9ac8221aa7d74b4a8b9002579b5aaf0ae155b74a92d26e149444701d3789f724ba58f4589c4cfecd4475a6d0603dd33fcb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd4a047427d8e8de84b2f2cea09fbc8dd8530e416e06f4e481e4944b4d76fe23488c2f85bb85276594391f6fdaa7e91a53dc9a1cb48f59e2b6a0b33df2a75a699b0364ca7758eb97a253e7171091d0e9986cac02599e1cdccd39941c3e7fd6bebc86b7c0ca9c57367c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h50b592788f8fa7d6094f2e9218b0fe589d9d393edd0bb6e512f35ac1b1f9c303468a35b531f66d4a02e21ca200e9e2c33f975a4bdb8b2313144024ad76bac4b59130a48569f7626040f938cd6d8c53355851fc857d584ac4060f6b626ea74e9b50a498bec6fae345;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a4d1813435044571842bce24284d93cf53c89788b814e1f01ba28e7c915651bdf0c6065e1c6f67fe0f0cdfb5125791e32dac8a6bb8f340c04613d3e7ca0f0b7f8bc2ea288c43f00795e1fd05f97026ba70ffc9bc75e1087840305228344157bb9f86bd43dafbfcb415;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9009c43a0e730cb677aa5619b8c2fae379cc015d753b0c4b048b8e09602aef11cd9e51e6ce91b9845d5daec34a88f0b18ef2c5257eda812da6584b4b051339163197e79aa7c93dbc73cb496bced455dbbd2d17ef1fccf3bd86fcc6801fda91069b1f181a78650abb34;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha526bc824a1da8e3048aa0b562e281c0b3b6412930352d286a32eb0b2eeaa2da3cd5cdf9a755c7bf40ed6f4095ed45d903c37e51a1100afc061e4622c74f7a18213c6843fbcad7a1ccdcbecb7a1e73fbca26ab05d15fff642d52976c2152328ba745e0e3c7d65c0318;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h278cdb85e415556c3e2f7a08a4643db8abefe81c6e84ee548445aaa618c6473299fec738cbe94359c769f408aff190ccd6b8302ef7b01580274eca306e21cde2fc6bfc77eefa7dbd21ebd0e6a783041e3bedd322d4e6755792e869a83b34e646a29ab0bfb5afc2878f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h129e6589648f0d0ec3fa4cd680966d0e4110f007c46bb8af9fedfbff8de339bd66e17d88b33b4615e6287782c87f684b24141e90914a470ab971e6d0b6cfe2246d9c089ba33dbc29114442209c291b6a81d910742646f5a38420a880c6d107ae166a22b2ebe1cd4f84a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd64e82d6f6b7fd61a901b52e3d681c275cd64d52b9081cf1194c9d157b97d9243daa3f54e90c0c63f4183b0e711490e218271945d5abc83de09986b3a1d7a2f1e6cadd03c4602b419d3a5c898fcdd3dea30d5f29ee23087b234758e429154de17bff316f38474001e9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113faf386ee4d491f362858dea9ddc0d8c9aba06cbb7ef34e939c000b4228565c8bca75f1c5c5e7f0dd6d77c6b7491271534fd88af709c3ec7b15ef4a3ea367d60ecdca28e1a67f335cd4101d41762a5cf0c9cb520118514ba1692bd130e7cf6ade2135b79574ce6380;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175c7c38855843b3a69cc86c2d42a0fcd1da414b7f53ce94eee3aca27d899fcdb9b43c626fa8d9a4bf6e8dae2adabd089ecadbf830e943280908075182096aa70084a105c134401bba2faa9371fae6274f57b2bef6b179b78122ac826515f336c0a2b9be07cbdb91ba2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h165bd2a20d6205d9c4bba86652826512e8eadc3757c326553ca4f3280aea18c6fe6b21a9ada7faf9215004c8cab3d8e830c45859524d32856bb3b8851815226bd83b8ca66442b51cad93448f80a5703b8e41b801ca6e10019a7e9bdae969225300ecdc85ce98e40a9b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f9a6f2a60a25fbf44300e481068e12f0b4e17ad46e8f64b92cf269ddbf2f5fecb9f5663dff631530a36b59fde0d46528325ff651074f8b5a12d639bac57de36d6f760bc7ca2b370006587e18713b8e2a051a81cee51e0e7734edba2002ddc48a9c8829b7de534f3cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f99635140e0cae8a7016388b4a6cb361499ff7bff358171ef5d947c3af56c07bd8e8abfdeaf6d4d32fa4cd3a02543bc12825f1899daa41a4fec9d4f648d9690bb85420637a0d61cdc97f395ceaa18996ab2222b773f053ec45b3d4f3cf7ad4797d55f71a8e09d84c7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1735b0fc5e7ea1af194da7c23e101c39f9ec904bc68143eb27c6048789d38b9ceb75af15a7de8d69b2afa1a7d82985e3e389e610c8b3ec81039916741e13d0e9cea13bda73a843f6ef860def59bf7e5d7c25964d71ab15a064b662c06ac1661690238a46ff21d1b59bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15494417e84cc3aa85155df65555cfa985ce6d25466aced31c747e268ae90467f883b28efc201eb77655748e98753c7012880c19b285672a08f0ea93527a3314e9377a474ad1facd2d6d17ca9d18dd0f332fc75e6a131f681b40e68c02f11c1890bc7a9f023dc226e6d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h66420d261c2e7e58c3678e324fc876c7847a04b567c0c890066808d70fa027b588aa6b400b51cb763f3aa1c67c95a26943ad22b40c9f4f46a10b081fb69cd74def91532f4ecb3aaac73eccff32bdb26e076eefe1308c053910ee47a3bfaece54e23f87fe717ea7b0bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h987eb0927283e01b1ba28506bc71634f7f586b227adc588694d958e1d9132e0aaf124b3f83c0e4100bfa52f274e6593cec4b91c3bcac8f2dc3910f4885209399deaa60965c32d8f2114f1116884a34d47dc497b0a3e107812cecac134cce5bf50f94eafe6b2cf7e8fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13926fa5bbf481e42c86ebc284fca280e94c2d905c26cf88894a208033c685fbb0fb4f14b4c1982c9f7800604ea62db0597a2109f67c10a49072fa1849ca9688db10598291132d666937cd2c518ddbe00a15636ddb47a022232c800fc00d3043d795540eac4ce8393d5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146594653a6c5815677d338f0efc1906cdd32b93af22182c00e481f17ed6be3fcc5bb4c2a8e1009d5dfb4151afcb2387fc77979c2ff5c8d30f3d49df1bfee43065cc971d305393a44e49e0c266e2069ca6090e2a23b920e15a526b3b1e54c6cb116d091e816350214da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a19d6a0bd74eb29f26ba99c5f660d900357e40f2176ae3beb8df43b4cf568fb85948ed65d8bd2dc907eb49622ce3876f98d09022e48d3eaa6efd508779c0bb76c256aef3a715bdf97644eb27d4cdba11882b2eff9a402be9df28e54c1a4c6065724873e03f321c1638;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1252f44ae530f39b4affc13f2a586416aa8bd618acfe8a68b769bd66a68f5519fddd1d6987f50035d01089bcda534a3ecec6d5b5381abd7cc06bcf7e952f76cec42914ed410dea47bce52396ee2b5b6e390e7bccc099b9c257eb281cf63170a20e1290040e42c0f8b3a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42a4cf46e7fdcbb2f2e4ca84191b0f84fad0a9270559d10b2baa3d6442bbe73bc0c540142ca344904e044db8918d39c96b42551f37eeb0481fba4d8f2ba3c35aa0acf7cbf6ab88654659d13289c9b976684aa184a516f73e9c92cab6db9a081d26d5c1b8224df0903;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c2a4b584c134e3b89f1578d21de44ab846a6199f5c366f476e28762e153cd26e67e011b0df8502968eaf6631408d073570b58a73abeb2e04139d31be8276ab1587313f6a547d556e6d1a91e153b78a37f6f0b1de70462b2b8b07c2a572432d52bd7fc426ea4e8ea603;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1294c2207c2eb267849332943ae39298c5a74791bc09ad82578abc50b10da2adcf4f47eb157a854fb554dd0cf99cee24ce4f37df1f45faf6f7e39afc11057cecc04ebce180d052d3a0c86816fe358901de22c9890f066b56730646b7218582b24742aaca927b3a881b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7833371419e6802664d953423b6ed80f9daff6d41617879fe15ef23d666f0324c0570fc50121c1c18e1b964557f222eaab89b7530bc15331151804829fc7262463ff2c528daa8fa444a4360bf0634d430b2b05ce8f93fd03da8df3beb5b5d5c8d39741e761eb96dc67;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h554e4919df89f04cc4cd0f7f1edd9fabf7545f6fa05cc21ada5dfafcc2b8d1390a41ff396dc8fd2b51e4c9ad64d1bbf218099edbeb543a3b65f49f9fa67686a52f3be738f7affb71f3d8f644a326f5f096b160d3926cdde9739f7e4e47a241b1f4ac6998435002cf1b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a9f50200880ba3c81fe403a072bccf4ce29ff137df910610a6f6ca7500f4a61927a56589320b0e5083f8147ee0467b4eaade64926ee269c158755fc2f316b41024cd936735aa7a176dbbede186869b0e63920f014a04911d6a4f9c847e8ff83e636fb6d9fc3bb647fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f7a01362d37edbb88de7069bc6ab3fa1e426d614ceffe78ac6d34d7c083ca178ac59ffcd959f2298f8ef767c32d9b121503792870e1b0078f6bf176b5f56518223f40141166852fcff4587cd332aaa0eb01273fd3f013bcb8acb36fe7b3cf4d3ce4a27677c2a35cd64;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haf10955beab2cf6ca362052e07b8f4db906fd48288c439de534ac1b617f6bfd71bee86e78571f9899a944090251d078b2774c1402c8e70101f31d6aebcf1d327f0fcff5b8dfcdcc9c643b8101110c701d8c829666b9c62b840e701ba51c00272516c80f88fe2d3e60d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb83d4220378646a74ca1572bdb0235ae0bfa94cb45f3bd09475336056e2c950f3c72c3a6826c6ae270b8034b8841682ebbeed278796f52830fe0ded6a4e0a2f4c261e25b5dfd7fdd9645f2799d4647011c8f4ed6b99572fdcbfe753d3e7c7a373c6e3c07f5db0026ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc13ebd634ad4ac565dd562092c5126a8f5480da6ba3d3e77145d5ba738d80c2e91f3a24aba923489852a6970f5b596db23e8663c1d791a9276a772a6d4425e5c934eb0eecd6a04fdb0d2f6d045b09f3cd4489ac9396c558b2d59d352c47c23ee37d8c6a34b2a671f38;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb699714d9b6fa23aec018aa431bc218c6162862df176d2851e2bd4e61a9acc002fa2fcf82a4cf14603b947d93bf579f03b5843b6b71494c00598e9d752970482278616e4487ae0ca73b8795671d7e0f1c77ce493e0817f9ddc244cd4ad2f2e0fae9645c41ee1d8b507;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ebfe1d78ddbb9413d311945ad84ec776ddfcd03eb94503e64a6a26b3c03f7f6df5f45775fbb6d8fcbc4a04dacff33b4f517c588b8aae4bc34d2ed2e289e09febc92e02ea05a0aa02aa96eeeff6b6aec9c28eb2d2756d662bf04a9d261b6957e2abd737442b5c8daa8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11668a42532563e03fb5dc540f010114ede7bb4f2ebf14004fb16e0a0b6ec29f8179a3209725fdb284523db104711ebca4f86a39bfcc336512c5a0aae97512d331dc562fb0eb31240b2ae1c999174ff1ca0af75b3f87a6c041d5e8818c001d70cc170460130411aaa55;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca1f7012c6f262ba5d5c1b393286c3bf44e8f7eb2e249ff7f498ea92d78077a5157cbc7894cca8acee33318f47e58a57825b43a58fb90c03026c1227d52afa4b2cf548d87c89614171d6df3144e141d4c3801215d42423fa7c5ad8d345f4959a15d0ecf1e3ac4948b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h160ac15f383ca7bbac54cff3041bd35eb23669d9333bc641c393a5cad718cbdf960caf5d1b3651de0632b6c180153c841e1890ce624c9ea50733e5a63efba3bd6f854d75d69d6bfedba385a0cf0e34ca1c9b13650b370182fbf229e7cc1780800e2e5180dc4ab143c03;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155369386e1d3e7be4c1c96c615c7608a7ec731cb0a37f8d42fb7d8a975b603a6b6c7c4095ce9df40c80e84c35524695f50376452f6493c45eac1c0c142fb426686f3a78b2b15c8614acebeb8e0327010248e0f1817718b4c9c7842cc859625666a8ec3151e78cdde0c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f624714bd508ce9c0ceacc41b5d2f239f86a4508fc8004139d9b8b6b575caff86d0d137eee5c512e7ab65031aa6130e6d8690500091b79a9ae3ee0b9c44e8b437156c30b2d66adca23fdb0b7a66bc8c6b808889f063e37aa992f8ac3fd45f05c10e76a59317e054af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3764072b678ab5d472c208087634a5bdc736782afe91c4b081f69d65c01d9f22fea3a526e9ce5400fe3ec8cd33ca61bec7fa414a6f25b4b205af350047c16dd3ad68b7ed4b5ae2986e7c14886ad223640447c1d0bf78405f897cfa5b62f7b75c16943ce7731a75697f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he2d194683dec6d23fd8e9a618aa5178e85a919a4393088b60bdafb274290cc6f1734110fd292c50e6351ba6887a138a59457af2124b25592bd9cc383dd6835532c32de0fe6eab80de2bf3ccefb4f91c678d96ee974170cd2ec1f124a8b6dd430c25fd1bd1526fcfa22;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1afcc2191064d2cb28e7638db2bbef20a20dfac9e39e8f9da214de415739a535d832135dc8db775d9dc4b70353e92e842cf279a90b289352674c2e9ee1ff8969a9db44cb19e94d5f2dc60b4665f644fd10b15002dc4e5bdf72eec9fe8febbf88894799c2c6163c4faa7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138c59b3a02599c58a859db8930bb1037cea2ae5db38573a9107e33d26fdc9c7af9f87203ce9afd8ee04a3fc2e68696c5758f654efb7eaee3ffe4a7c7c1ad144fc75d9338f1b604db9c2c7c85cc51dc05c1595a0ba1cf41a9a905cb88b440da1f3305c1d336be32ee09;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cdd4723cc09b57a8b9147fd2df6af8c6b65fbb56db19ba9733abbc5c545b0ec68d6cf041ffe31b8ac081bd1b04d7ff8d9162120371527c6add2e6cac665c3503e9b7e3c4b5ae7e71a0d0ab60022c43c0f8258ebe638de4ec2962474baae665cbf7d14e77e82f06c530;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18829e0049559d532dec9f64f5204e09396cb3caa7ab34daeb68985d0aec8fb5a77531df50eab1c1f95edb480db4e0af6c7a79ffd2b5a84f4ba8b5b00884c1949ccd8e961fa0dcef96fb01d97a6f5630628d7b774946f649ee594ac9e6a4d0116606e44ae1088ebcd4c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h938aa81878025ebb9a6eabacedb69ac7d8497d8c837cd0dfe7133de77f24a8c33c9af4099247f10b79a0634a517fe844fe7c281dd86addad83265ea6f62a7bcfedf0b496ed1e52912d5b0a2e3ef55ea6e725125d93d46887621aeab3c455697f691c3e01910eb46631;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2a4883254849c170d52e722c2deac119db29e963f5c662fc2d2ee5bc266d7ce22119396d8851f846fd53d90badf14244877bbac6086d68447724a72a9f01e0b571f8f2107cd66788e512cb26fc45279da2b916521f6ff80d67ad9322999b0f44bc0b58e00682739686;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h192ab0dd28905064e06628aacbf773b3ff50e417dc3d34c9659da80b30703b52d8ddfe9592a59968d23eab1f84648bbc815201ed7df5762ee730ec2f7b4478d3751258fe1e34381388fbd6ca26803ec1d7ff93adf07f91b8b1a3a41e5c94d09e4d11e65163e1590aff9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113f1fdf5a213eb312c7a57306d2fb91118ef2af6c898982cb4270fe6c99d052c7f05bbb22db64c02066f020de2930bfd11bd0acb329e3aaba4fc77ae43f4f86f901f018baeb7c5624f3edad3256dfa0a55e8714c6ecd559b5cc34a4957616d4e15296c111b9859ffd7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1314ca5160dc01f85416c608d17eed57136e0c841ebf65529a42d63ef907ab287b7708bfac1cfd09458375514f8d558a79f94af16952e77c7fec3695ce967bd60ab31b4a1c66d0dd143fce4627f33951b23454acde79e97082b6cc86e33eb4e0ff1496099f059e697c9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18fe653e270c186ff01ef30b41f6521646adb638d87d7a50cc0e07947f225631c1d9d10656b43f27ff0baf499f18fd4516d8d8a780444f23f3e010722dd348a1f1eb4bb4311bdf7ddcd47a2926f08baf169a465f57df1cb59ec679e1aadcf20aab6b9b2dbee27eec1ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1954bd3688a08bc3443bf760610e5a0e0710f76535d82df5cfbb115e8b58c707a95c6bd1e5664c26b41c4aaf1a4d38d5160ff81a096cfcdb9168b1ee5681152563bc45f2b8fdba9fc70577698a4c889f9d6dc1c99919981392fd1bbdb039f91d3d47b0e1d64efa63fe7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14427965924a63e87c07793b83636d15b56852061bf148747f3a88df6fd23485e3c95d75ae311dc4a4050ce890ded9be58fe878461e4d483d52e680fa52f099ba4fea0b3dca7a04ff0b5b687283b5ea101a3e37c636a655b15dffd71175f35c1f06961775c4303b9638;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdba01ebefc2085efb783780551f9380ff37d8c5c34fd7915425fa02a6d71a41da94c0b716b92f30590bd8083b9e8674763306756de460df5c99b5f9b6d4268dcf61418c49eba50ac3dbdc93d81023df484b13af86d70614f51db6299c4e17470c1d5a198805abbab48;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he2baec5ddd6c99cc4a3257f2fe3bfa6ead487604c38208ee36503e3412599617b4948072042ee1df0bc4e3dd805d4edbcdd22d6a4a29244d3e027abcba0a3c07e31a9531cfb9b9c65d3e8e0a7d4f7289f11ccaebd400fadd8f8b093e17c2f7c31bc8e25437a0015b7a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163c626377c7d2ab84f6a4918a1bc724c2db137720adda8dacb850e5effa712bbb70b02294db65237c8720b2b83a5e7c17978a90bb098b75a794cdb63b105befe153953ffb6af8ed545226bccaec4470049efc90b52eb852f28d638fb781b829fba413af5cbb101c263;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c4f45da45c00f36e4c4f100f5d18e03d7fa4c2be4205f0f442166f2743729660b84342eee92524eb31653ad2823b3a4cdd5a36b59185de329f6b8c79ca7fda8880815865358565d717b9db9d15d0dce3cde07430e218df17db1d594abeeef59ee19ccd395bb1088b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7dccf09356ad24763a317561082dfc1f6768265c736af8f6f2be3d0f0b838d6619b1919000b9bfae7f6f5bafe0e902f1840bc5dab9a201752030e9f238b1bd1f34396b17aec378f10f40382ef8c810e1ac4250e23f740fbf179871f09d459a973a7e7fa2333a01a0d7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12af67c12b49a5746f0b349b2bc47d69a7a5271d0c51a82a8817f5d147c99b8f2d12d6b5d0e3cef2cca16b121b82d1b9e14f94b43862ae63974faa14779ad29c0738aeb8251067072e76256230675728641bee13ee9fcb7e1ad2436b2edf53089a92096a4968e29fb3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8d2405e8ebb805bad17b9ede9484c9ae683253714253ba9816418470414a98f374cc2123340faf6350e5c18719b8968903175c4e16b5c62b7615d2d9471f24735627f2b20a5ae3fbf9b9fd13946faab3a621a23b842881486f68bd276be14846f5e1e15d7ea051276;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb54039a4e078e07b86333f7e48ae4a7470adb050a600d7ac038bc6483e20e3bacc5da145a41cb79904ecf8798aaaadbff91c987bc385a602bc1241cfa79c4d4f85b96c03cff15462365fc09ab45cf43e5dcbe6f2b3edf08928ea28bc2c499af901df065bd5c680e967;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d7a04540279ef267e2448e40fb734efd77ec8862b98f1aa6673d7200574a7d47913102a89e32ea703cddfb7d633dc64516a44e2c5a21f8fdb28de190143f706c4acc3deb46ee24d37c6bfa31ea3bbe6b3f8d774b84f25a6332b9d6f0be1c7744fbcace4e86b9db31e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16fe640bbab161264382c8121eefa2a11504b26be29f75a07a0e7ffc1dab99aed227b96943f7fe04cddfc946c750a868af84c9b2adfe4630fe5be6c53e1d24e1e015bdcea392e6c718bcb308f7b194e509695429d7843603ee0b1457609ccdbf43dca1c7e0c334d24ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h85998316273fd677b215a48e417c670b13231031c173253220fd1455b96896bf71f1b38579bad678eb4eb979b283e354f04255f319b3032e47957107555499b21d27d4898e8c80257347c7fae7417269e93d394689d7d864fa3b4187caf8ad3fc06cc19750e7188bec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1789ea3589d0473567355911b268133ff870e2b3209f8364d14a397435149dc38ab8e8ebcaade53104ec5215e88e29f0eee4f5dd45b1cb3484689dd475f7ff42a02921b2ef59e0e100ad0aa4eafa00c33fd29d6816285fb7923ef1da9c32a2964a9a0bc349bfb55993d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h119fc42e878f882566e1a12c5106ec31ae402986feb6061949c2096c7ffb8ade7fc4d0d15b786ff04da4a7dd9a3c4a6eceff7a6b19cf56518190665534fa7ce21317ae41596407fb2b0dfd0f70180325983f9070b7d395098e38a4ef3cac8d133ad45ad009451e416a4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ef6384a1bbd84d51229014ef48e6c7b79f7f6dbfea012ed52ab83948f6d56c5d043b1661677f69aed15722e9c77444ef4803faffa54e151df847741609d2eaa655be085dd33387f0c42de429b34d445f7714fd1e5b4832ffa2dd184be236160da2b371799f05babdd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ee2f59790332e442eab766db6ff247d8b5ef305c86148a9a06475dda78299aef023b9abff3152e68052206e11846693e7eddc15ac1a908ca3c9909dc440165f7450fd3029f1c1bd7545a488d83583bff8c12d014c4833d521f498e1ca882c0a35ca4365d30c9d93b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5fa6ec75de419f4d6c20c066e25a02d73eccf7194654e4333b2193ead25b1fd4c15564497a805ce61e2de7625175d6eb111ea3ba26f2ee9dbd1d7e99d4196d7ead904e743c701e9587a7451963484d665a83be7ffcdbb8a812ebc2a9a86ce60abb7fc68e1db1539554;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8801fbe21f1f8bcb31244fb48388e91ecbc525492de288b6170566c92ca9e2d845f294b8c1be2161355efdf21014f64a2b92465223eb7722e019ba0bb423e5bf9d701045e4e6e36f066ffb7a764aebccccab720c49e15c85695e761ec5a6f2d42cda3f8931ceff43a8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19ac7a9c012e6f9cb45be154bd49e704e32bedd03755115e4e2da8fb4f872ad6a4d24a0ee3aaa3bbfe16d86233e49f7b51c58f0a1bd74614969c189c039985a13436ce1033db8cdd505b3513957d8493bd91843b9c447a9c4c7fc9778ec28077d0cfc32a3150dd3a880;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fce15b354c5a5a9bde3bf91e077aea1672468fb73115ee83e90bd691c17c9bc988c07ef975b3d860353219d33c8dce120bf8b9aa5823fa1c895f4e68d0c4253fa0affcfba032b3c571b3d6f866788462c1445a9ea9bf9ff63e8cf150bed5920a483c638b33687c66b8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h151e722d26e966f28562053019618f3bdda0d3eaac60d0c741c6c5625f84937a735908560b94b7541420363f0795cafdc4bf1b1097c43e9492c7a452fd9082348116a81da6aa4fa0dc0cd8e551b728984955942c68771479ca6eb1d135e2a216bb5310155779a0dbad0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19de74814500f4e05f29f024ad68016c51e26e73c157fe22b7ebebbfdcda2f7b29f4aed8b58a31c8a19784a241e7a423840060e0378d14cdef28a64e6322cfe3f5f7667d43c72c2c963007c7c4730b0df1fce0ef2810e9a9351f8aef7bf9bae2ee2fd51f55d76bd07b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b92cdcf421ba513361c767150f7d830976026af76166c6cd980fe076c70023d5a09bda1b1a18f7e9a89208a83157d5f70fc9ae00b01795b60c8c5d888caf5eed4c6a4ab9e6e16a9e5b2c3167667bcc34d9d43b4075561b01ffd702e26d1bf7e55f5643556ef8d917e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h289a905918ca94dae80afa2b0d55aebf4d23ff35d4bf0f306ceda379941c70f9795d957fe968b5cab41a82434b35f7ca377ba7d8a0839dd6ea8645f69814abf99d88e77053408dad6a6f378637788b9e1c2ae3f2d1e6b66f2dac243d4c5506b6e9d31fc02c1875257d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0b74d0e9ac80f0d5846c4f4b02c1ae37f38ecd631f26264ba88dc5b99a4157e6d2a6a4832d3ecf022deb17d539792da8ec535f133865e24f6b851b56d0f189ca6d75b64e05b7a22b54e25615fa6e74355ae8ed1ee62ec7f779df5588c9695b1d196886cff5ab4ff68;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha85a4e837c8faa568cf33aa9a84c402844755efa1877e284bd7c29257da98fe62de79f5a7d22dd74eff2898020b2de28c6cb9d4c895c0b3cbab3bfd9e0096975444c80c1b758f35f7b80a40cf941b431ff6c321ec913702544e7ef730362e3093dd7236c74d7ca45f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h186bb66ae6d3f5efb2eb393c0fb99e30db81cf1c017d01483606c4c640beac06c08f67d418b09185a89e751844057dd7fffa616ade4fea2a9157782b890087c52cf6bcc49e6b499a97ec1111faa41b4924bef7dac8b2c7f63a6c38320a34df9a4229066496a98c00209;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13286890f4bf24efc0e35194ec137e5a48b709d902ad9c50325dc5e684f7ccb8616a4eeeb492216edab118018d6e8d8522e8cc22baf7502b5b5ae027b5bdc50da3f17fad2315ee157bb98f4d810b5dc14830c7c22d842dc1edd73108b0700303f0e2470454e0a076ae3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17f626f1c65fc6851c878d473b31eed728ff4c17acf36c937e5bf491773d71bc287d0b94bf4888d0690af6c47807b40cdbf663d51b892714546d61a21b12f473b65ea2cec9d3490f3d77633a69f57309d113cc9b5142a88e6010b5775980b6f1bdfcb4a3c6a7eea3d9e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h120870962bc993036ecdbe92966d972827fa6cce7be2bee3ccacb0243842500fa6440d56bf4705243829d1314cd682eb48d9a38b4edeab429c70305ddce0aa22c26d25bff9c399b3c207c38bdbe3e031e3e88d8a6f914a718756e209f8af52d7aa6e24a480d25c2ef3b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a2046cd6b6dcdf815751150467d5d2ab07816be92dc42b09b5de622c04b84a5897661a44194ecf6cbd54c6b07f6bcd971ec9421d7b7f1ef0bf0bd801b09e159356db19bc6149ecb138a41bc3c3622a754123a51c0267ff8f35068e51983066bde477d854a7a2809d88;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d33d9a241b2f466e9dbaae9a9678a9dc9344a5902a6cd75fbe3954b638c38f29ac78f61f46e3813e411c46b8138eab041274032054dbc101dec55b4880dc7d342a46b0f485302c5647fcb7432a7f507e7e745ab011c6be3ecb3be27b6bf10a4a4aec58a723fec816c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ca2e7207d1a4057f7d57ed5e33205ea4db5880754d3ca3a69f6a79bdec77422cb1ea50a113745ae764d4c13b21a9cffb558d8ee075d2ab0aca86261c182134a992c837551ddc0005449c944526ccaa046413f31d0aa98a82a566a2f90ba656c0f8114995adabb896f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c477947e280bccbbb4a20ac459524e502e7f2095205f5bca1ac40bc5f173e5a8ca256040217ec2854e6eba2e96bf0950d95902d7b66b4a130cc7d941bac25092059de0ab3998cecafb9e6ab0a7df074e1b2b4c46c5f676fe92b7829312ed9bd69cf1560c77d213c81a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c077e62970eaa9f2fba11ed5366b8c5a36868d286ef0c7cce0f44cd6191341420f53e0da25b64dc01bf5a7c8bc2414a1525d6fe8b94f0b8edcc7892c2df89ba3626f26572b4a08a891e137a0ed2702cf8e6684d851646b187f885a3a29492123c2b6ae6ef348f7104a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h924556c4a155e1b3896ba4d68d9d2b37521bf6fb196a950339ee0d0d86905522dcc49326daaf39594938139ee361fe474b11643e604acd7d30d0bce5fb4f792658bcbdf6a2756f2c92fb597428a5079d141a7e12993d50650001cff0b364b95650e4f10c6c3be6c08f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16ec0e90542f0a84902c6c56a1af9b86329dde7b452aca23db530b95f3633c2d392e2e834e635fe52043851fccfc1553f36698b08df7e694156cb2f2bef96dd9751dc84b92ee298d7f9d7f969ba568dc9363da725a6044cee96a92960384f94958b6113a8e1e9a017b8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h115a2e2d55632d816e88f438678cf8caaa8e6c6afbe829f3721baa6f87632aa6fb11f23e9e80087820c9641dd04b9aeff5c784d3e1ac1fcb027e80a3faa307b622d65cbc0cff3b6c2d8beae44af04ac3a46d4c1afb9bdad2c4dc102b4ef1c58482273f76ec80a3fe5ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h77651f6c27c4bb208abcea7c0a81283985ab3224425e5074cf2b35adfdaf63f357f4113cceb8cce86fd88ee5eaf56cb938cda5187f5d36c66fb0d7b0eb679cc6739c76abba6ed654f03321672cee5e33a3487aad09f5c9dde0de9e828524f2d978e3dcec4415435a07;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17ea8754635ce2dbad7b7042678f90ca6a4791b1c2cec4395bf7d7af392c8120f15bf19a8dde9bf4801ba749e6c27394ee07632be786028036e300e9c16f00124f3708b368efb79ceb91fceb4edd081a620674e7fd0be8d3df33f99684fde97c8f861965d2054e1ddca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2662d8944d06b00b3ce7dddd2163183ea9d6497b98daf1e86d8046aad28931805cc52feb9dfe829ea25f7cd2b2291bbc98fbd47f33bfe306c0290d88ffe76806986115c2bb0d128386971a9354a20dd04a130b60a75b81bdd6622e6cb1c23d480c46894d5fdae8394f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ad39a8e10a8617bb010514b8cf2c5f08d0d364fd93d5423ecd858466cef80b59510d32fc0241d50ab640cafe387cb8c92f1569bf991bce7d4a6113dafa8b9f420efa90684f55a7072b70644417a50f26ee5c36f1c83b589d02776319743d1b707725f1f83d371f121a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1938220194741ab23be32187cd95c2c05345a53551ae40889e6b257115e0b6af5fbd7fad184bc57557f6edf71f571212c03eb6c225661c03a40035a989d01eaa5bafb88e393d6d014060958d78898633130d84a7a1d48f78bd03f7a4028b862b5729d274e34680b9679;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h41bf580686c82476b2c7a368be64c303394dea73554ca1322bf50c7fbed920d65ebeaca574ec1dc543f5411b6a9502c3cf83c2b5bf3514549c8a4b28c082a946de4a0ae2a9450aa2c6f218968ea76e33da4df86763bc5819711aefdb0e7b9a85ea9a76d5f07bc94a04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h432ea81708398f56a93a96a1e637589db577b08b6460ef1020dbba17d774ae8d4113a7b770af16f6110b7f3ac1b93595cb0fca7e4dcc8b53df01e345220c30746647744c9ea75d13e7fab6a7a1462b72889407f6ff6862644051077d2cb47a029bcaeef5d8787ef0c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f3abf6ca125afb39d10f1b6412506950c5648eecb6a93b39c4c920bc65c71070f93846db7cafb5c90b6063cf56bd8a1a9522184b887c0a6fc529fe702471d198db9ab5651a6b3320a1e5f08c543fedfe4ff9f74aa52c93364aec086f9b8c9a48a43ead3b482d8e94a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h212956bf5c2b1d41e0ce724f32c52aed18e3e6a454840a5959df7cf152604a6b85d84ff159d7306d3f11c01012975be7689ea7c65422d49b9fd35cb132819876901d6d31803f9670e85ed79adb8b16ef23cbde147c0f2ae8f13522851d6ad0a0ef6e7da9f3b43698e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12e011b6d53c8f83d9c0adced55ee51a05285dbbf0453e850c9a8bce141c72ca94f497ac80f91ed8534972239341fa9b72656e5ff7f06a1f89b2dcc047026633659268f3d80c5117c4f5a2eb7ccdc67fdac3910addf4d4915dfe00124a8f6431d031e0b50ce34271c31;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf9fa4e6ff842c77fa99496018867fa5903e078b8d3688c1cd1c52b0f7bfd3930f039b742f06c3ab45e028bfef77d2266dbe7f8de9dcfc540dd129cf378859935fbb8a031390fc6f848a7e97a2ec7f62385d64c15e4f0030699edabc3792ea42747b3d505eadf082d83;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7cec432aed86d3d0070f64b19f459ebdf348b00a4d39e91554c476281be55318db02ebb20b006fb17f8159ba1b0e1b9dea8dbec449452b2d6a39a498799f68616d648e3bd3ceb10a550e88079376cc2be1a0a8198a77e47020f8bf834f50fb4ab53fb91bb9d44f9aea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1945d6608b3dfc6522e0f72aab87e6aa39e01148456fde49de079a6f87650e692ad4981d1490c207b06e2b502142c22547688384dd9f1124c25f8c9f4cd3e13fd03ac8d02fb84105c15ed0e1cb0c1feb7d0c42a4098aa033cf7933f20b0f9d0578d58fd6a4d962f9fc8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h54a8b073ab87fc39676c5d80b20dca6e4a138117f62a3afd76a6e1c8aa19211278b15b01f2d96f3c5d776721639bc0430c28f76da1394f55252b8275e6ec7d157b7285b0da49a6ce0973c31933233a06382a427c74779baaf26d6e1b7c332ee6052991b232ea59b806;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h640b0c759aace096fa0e80610b5664e6b9b17604cf7e19ae2664bc84c8e1b15b6061f2c918960641f0c6b2aea1c7e3b04f7c93f430d837d5b44200e91bba07954f532a28b0db68dcb6e0e6e85d762f8df534b0be1b5aeade4cf0aeadcd7fe43191015f92e67b4df50a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h39dcfcb0e7dceca97a2ddabb50e64b475684d21d9647902becd28ef24672f79efbb0430e1e057d0d619a9e3dd64144dc7f1e18c7d37a904036d2c59c0a7caf438bacc446315be969b477cf7a9052c8418c23eb4ea63cd4c15cb965bd868ee0f74c7f32e64a25a5bde7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h325e778a55fdd5f473f171418b7c090685dd9e27d401730ff40ab49f0264284ab5aca73bda4323277661fd04b819965740aef889248d73d27800759a71798535cb4d7e2ed6a66fbf03e4d992999ed925d28c38684a40a92371473e83036c078acd72f9e69a89bb8e2d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee221738899cc502d61ff7951221e437c948c6be11db08026d36f6ae9c3d85064588e023e92385a1d0bf2798820300286816750fafcf7b906f6e33ecc779436e685f8cff8d87a8835b1b18a2a12f1fe1bae05061ec65981462bb3ca657b5acb8d85a1cc8e71588d194;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h31074f3cb07d283355eb780bb3c52789327619524c819c482c8605627e5a59e647ebaa119076a407666089c7a5e85e1af8796880dae32a94f137f74fddc372d0f10793332a4641568a07f56b4afe9910331e1e7afc2a90eb7aa5dd4c84780d7823863ad38e2d72e593;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae22d4a978a197c42c78ad64f2605fb8165f81f5909eb8e01d006d8bd3b9b027530350397fdd6cef9b6044e9182ad68aaee593b7fb539fb52b64caad0ada1af6d52b63b44f03f8d5813331902788863bf0673c8ce0a6937fcdb627d4a0f3d8d6975deffa36a0381f47;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2646563a8b6076872254805eef8710bb6865e639582d1f546d3ca392716fd15867e1ad996aa057b4cf107b0b6df8bdc36430b30c294f169efd4699af2e6cbf11663b3b387844d38004a36fb3631a42c4b7fa9efdc8ca90c1cf443328289d0913b95fced753d3b36fb1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he768997d553acd75578dd67a1a04ad6c2fbd7b410f143edf4c7a13e174cc4886b68f8f3877c95612ca7f78d917265a118bd267fd74ca6279e6805b4c422e9c34566a44da56209bcee7a572ba4d687b1b1b9d9665193d228890b7144535183b1deb61922257b1a4165b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1afe2ee8135dd0e5d057f4d5b9f1b49d7736890180da2a266b9e52f08cf53295310cd64044e5a97dbd81df234d676a0591dc0193723b73f6ce5f3f4dc40cf582277308f6497e35a3cb9ee8b1fe4a6e7fb70d464b78a805116e72ab58c35a16876a2daf5a13436b5fddc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f10f1276bd966a843c10062bfb7060f27d34267c05b5afcb3017ae65505348e56ad878b1fdfe5cc7defb02956d49c7233b55972af27f0eac415bdc3526eef39d765fb620035658328bf73a8c60a30018fb53c835f88815c2db778306e97e4809badd22a41c5079567b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de0db192f3762093724e74cdf01c095e51314ac2b9efc463e7f2a955960c3edfa89978fa565f9c02d6b4fa10a897c3bd9299f5f1620da24b5e27da3716c0f2b3ffa4e1d7f0e6a9ffdab08ab5547a50e19315dd0de8e8179ff6b4b61c92de640899660ce2078e25ce68;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d9ee9c85ab41a34a6f16b62b3206bb321ad92bd333cb220a81b4e30bca319f14c65859bebc436ea72546c2851522aa3c1c5b6dc32860d79921ce07056e84fd2f4b6bed6cbd33f0250ca46ca15b9327b6cbceaec44e63b8f62085c09f58b6f719ec5700f864265c16c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbc5ee758b9a1ce6b29ea5a4b63a5d5f7612ea938fbe7349a46f90f2ff48a405d6ce5dfac6e03163c43cef6b79d5c43a1ffbe0db237537303cf968bd33020ff6da7bc4eb181efe0f4749c47e0f283c371cdaf5d3c253c75468d2a6292554621c1178772db249416ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17f569f6287f5b861db49e4652f80c4f6ea6be1e89c1517359b6986f627e5f3899cf680bad4f189a01c616748ba78566de765c3fedc1f78896c7d5f81a91754717cdddb1119a8ae6da59c77258262933fb1122d9842d6313877c3c0f971b8688c884d530662d68b124;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb2706228ac51c48d7705c7ece3ed390b088e38bc9419e0294d829386584ece1ac5e0fc7628c87a2f4013616d9f802573d1042e490fd480c721d05bce8df2296bb3d18433555d2eb5738bdce30ef4117e6ee4185b6349385a462c8c98deab3fefa70cde765b5274bb44;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fb0cf8837e1091ae2e12049d331cac395a1420142607f4f3b2824d10944e1b869e9a815da6bd693f16faa9dc425601bd18d62e24e8665d2fa8d88986448c4b8861d4691dcfc64b0329baeedf97f98f18e5bbe487539622ae9dd05bf9f3ce0ad052e7d7a1e2b1ca94c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a0fd294b29101231b2a06b1cf4ede9e0f84365122ad57152d092dd7f20b5a7e375ee70a8b40fd8e5d568636f4d5a7358df488b1fe4b2cdae13e0dd7116fce973a196fb41fdb47dbc4c044dc70c7254e9ecbf714fc9b1fe0275eca88d67f3e4470e9862387ccb0116c9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha1ca31fbb5021d615c8a7a1c6e69eae88e19babae5f3319cd28259e93bcbffcc1ac81cc35ce3839143ba56526ece30e4f801097c198f1d0a67ce2da7cfff6c8b425a4e575f668a9db9a138e73543de8098b2b20497aeba90728856ee1ec8a5c050e157a04c7089d1a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f45eb019e47d67fc8e016d988dad554c73930fb9ac42a0b51142e913060d9f0b3cb02da7a583818265c0dec5970b9320dc6e89b7f7932ec9314d0340c8566ad9e21485ad908709266457f92246e5040a683ea855ebd5e63102e283572696033b0c50300ca2a5fff02c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8fc81cd9613b528bf79ebd42b4f91db23c0c6dde4aa8f1dd7b857e9a46cb6f570796573036d24f749eb6f06d85036582594611f34b113ec4ce98bf6296b9dae253fdfb010f093ed3ccba794a2d2b391fd57bb22131eb1c21c8cff29abaf01d4200836acb8ee0a0343;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h21c50e803f14dcb61d9da2952a1ed8ef63db5f53d2b3a0c93f349e3beb51d460fdf66505845152b6cdb4feefb2261c15bd55f9adb0ce5da91002f4e66182b2e46720563ddfdbdad4384714efd59c8bc8e4c7ebca2c0e5a9ac8d249d891f6f3cb4d9ef11a8a109e4976;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16838e88f4ed8695f6512ffbca2d58f2215005f5dce0f67117338020fc30f4fe62ff001acf8e508d813ab93557b2b4664de9e1af8f8bbfbbc96fb672ed4532ae8cd9bea6cd2aa570c9ab3127b2c5e0902dba3db77043852c87d3d6ba6aaa6596280e3dcbbb825deeae1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b241e14b996611587ddd5f75a8c8ba77244329932c7a578ccff595ee1a3a7cbc119d9b14a5954951ad882675a9e0869e885f555943221ca3ea80b7c2b5123c76e56ca9c7ee7a5fa8bb37e617aee5016d63ee62ed3a95e7c88d733df15a8e247b9f5a259eb26e56925;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11aa2076f96cb724c2186509521518f7750d6225753acad335e61ae94a2b9cccaddb526d76a4e0661317eff49c0429297d1a84af8b60177c9348812e700fc5ef69785904d9090e4247d400babbf0222885e4df9acfd2a03b019398631f46d8e3b447c433ad1670cf23e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h158a9f4e75a6bf92da1b02df271010796b8fcc1a738538c055ca45e1edddee74d7474b41c9fdb4c23a9fbe02d0205042faaff885bd7c747ce6652ddee387088d605b0e5131d45a78e02df6c0d496d093fb886b19f0590158936c9c79368862390013453bde5f9e11b55;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18c366e44deaf051caff7aca997fda77e451749f53784259d64bdeae6a4576abb4fd899ccd0561452a8b955256c1e43841ee456b778a691d2ef404a7e7f909e72c96670e51174623e91e49c2f84da46b118fcc0413cc980ea3c6e1193b418824dbcf2f8a3b2e803d894;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bf56b0058765be7ecc3685c23b3e9d1ca20679f4f433d2cb0ed9164f2de28b0f3937f29fa08e628124957c045aad69212c14b78aa1464ce2defd0083bef3454d81224982f39b7c19f602abd81292b820977a61aaa923c9c926f04f0c0b2aa0f4e63479943c891b1376;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha3a41af0384d3c847f6d53c3a6883b6c7d6dc87dc29ad9920d340050fa895c3dce8689ac7cd51e2ab0567686efbb5e8a4a49de00411ac09674fdc7bbd7cbdf171b14979e8e7ae16babfaefb189ec26e3e6594dea4211f5358e8a530e193f029ad3316f0b903933af67;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ef375970c882ff0cbc815a8ff33bcf9c911f82601b2da66bcd5f18580851d0b0c54aaa6becc1665074a9c9e2d710c08a3d19368eccbe259b26c2e3076604f94a198da1f41009cad0290fabdb0ec51cc66dd10ba960859c4a91b113ca404a60b51ea0aac0f1529578fb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h117d17d1eecc7b2239fe8b334abcb63a0ef54da54193a6772c29a5f8bbf98d2f778f5c8aee3df72868e93c070e487992a54d190013f66fd7cf51e6a4498ee39df10eead9556ed3a3b5234403b4e9a1b5bf1838cc39d8fb205d194b15ef86e72745ce9f3e88dcee71bb0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f9cf1e3b21283036e39742b52cf32f2323ed5626cbbd88b40facccab83a6643150c2a94a96e696d33279321f3a0ee2c02ae79998f44779c84a1cc847d1d5dc06ee2ae8246c4630a310dacd4d772242bc8a00ce77f76e44935b7e6710cc0cb0097d83f2c15218c9cc3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h120be91a9c39e2eaaaeaf9929d4a47cea0f9796631be243cb6466a4a2146918fc462fb82dc1a0933c3aa4f500ff62d92553723d2c4874af717cf929ca5af5f581f3ffeb1b93e31c24a8239d98509b19d255f31f27db3d26b9fbc603ffa4344ff237d1bea9be0984851;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h191d2efed53ab0ce54f811c54611ec83d3639c230ac12a199eb89a642c7be73b5f71662a29d342b93d06eebc8cefc590ad697e20a11eb9fd8da8905be6bad77ffb47f50ae9d5051ffcc1e7530cb8fa12afd31aa44b019b1dcbfec227f117b643da8e224719de84723ad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15d253cb926cab8c1ab842cbdbbe27fdb0706866aa80486e6bf50b62e5d4bf6036340b60dab2231f49d6f8686603139cd9063823e1fda611cdf98ccbeb60ca52a41d7bde88067bfaf012ee5185ebd44839b4c70847023d5dae8223c80709e5cbbfbb91725c4ba5ac204;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1933e1ce9f86950a472816c255c341f856d9b3eaa28cd3c974de28b9963db834faeffc815f4f3e60e9ca3ea573fdb0deaa2d0339d90b19aab1e924b3e80ddf071a11dda6db9fb05bf6c17d97ddb72f8c46fa20c46d2eca2acef4afb35ae0ea71ccdb285c06a60f36f07;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he250dae821dd0bce8333f67216dcd466cdb89e279514330dd19b0f8ecc8ea624981c347a259863843e71e4b1d7cbe86d71827e55f3ba4cc7949726dcda08ff4465cbb685efee825184228b5513a03b7095c0f0d97c928dbc29872a1d8032f013424b1834ffaa8cc20c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb41adf8bb08d0f954c624d776841614f9d3c553473792c6e63322758b37c01a786fc5d87ebd46fb157ac90f3bfe6e52e3d21e8a88cb2d47d5bbbccd7ba0bb099e970f2800375c2a3170eaae88da9d81cb72731b8d3d32045116db06c2b507573810e85f419d7dbc873;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h191c8fdebee8be8109f19529e742cfc12f92d9e1fc7fa521fd7401622c77b2ee19498b03e8d49b9fe7867175fd00d8a5d10b795d952b3d32bc921ed2f1cc3a4915760bb932fbf2a1dcf8e948297440f6ac783ff0a1102b0032f974ffabb50650df095415e62718dddde;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5362c659a87ae66f2d5071922630cb393acd10237995cd1920849bf3680cb147cb61ccadfa263453c2b40b24c10471eec1327cfd0e56b82a8d17605acb70cb9c58cc00678931c6b506532be26ee86cedd178da72ff69454387034849dd64097a123007b4eb2585f4f2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h55456b1b4d202e2bd59abb1322d13e8aec5a0655d701142dd0190f75bfe86b1d780264a59b110dfafaf5c8feedfcce1fa894b4e986aa126cea49f8c1811a3cbd2aef256d28f5cd480711fe47bbb1ba98bcd722c6444520f3c966dd6dfcf877e796420f6da11baaff8f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd4e5ad6175a6fdb9facc40522e740e721787d694cf6462d96b7a39c70230a0c3724e48e6b102d81ef595be99d2692e33b50a30d76ee9fb4f5f9a323ac1bafdbc3ef5cf20d6b7b7ad42af0eff12800ccf205a442fa5bb026218f8725496943107b393c3bec565caf10;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc6ac1f761e2c58c07711af1c802e079b5a88905fc9f0124e4854f8c89f74ab486bff89049790f3a41fee871c1ed84b2718618cfa856365634b260e3b9a2a16c2507bb41448812250c57acfbe1729cc2ef5c248ed2d1efc56ea53accd5017ef5931b55a67ddf9b1ca80;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a89b35317afea39aee8f6c8c183ac22270b18206f333921d44a2c879c5fc5bb5908694b937063a27b97ff86e6e3d8941b1b55ca13ab3a6ee19730c529905393f1f1fff68630d0496ea2472c73a765629627664140c842ab44b513b2ad1b02486b88827ec1c295e39e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9080e194025e6f103d7e2bfef731c7a16f6a53ef91eed4ab563a5c0d4ec31444da164b15ca470304ef5ea788de62a22220ba5f7c503e0f45e55581cc84e06c52dfc643293eafaf52e8d2d9e3b4921405b30b4e168d160311dbd783ffaa9c0ebd6ea479714576c42d83;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a054253de8b26fd7d846187ce5e7631a4fec3631ee185c1fff2ed1fc8c2ae4bf76af13d9d08747f158e1407684e9a247e97149c637c35e785236a6ee551e3ffab196c467fc51b995fa812eb2717fb4b0e08952a8bcdca283218a9e60da6247e6e7c27e8229a366c01c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h121e488321c4dda5a7cc335cbafb3c7d733653b8a56db5ca9fb3028c4ab5f5bc55f23dd7e6bdc8d012ff6fac05a6e1ac5ae4374c7fcae86695c2b5ba34742c3bc51b0c857abdf02ce438cb4dca99f0ad6caa3d240be203d979636bca486095bd2a831ef8d27a30f3356;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ff8ebaff6f80cc081e55395f94932b8fc029dd998944d5d31e6b049de652e9c5c3edbd08ea31a8066afc5d1b530564a1ee158ebd7115f2c2ed7558a8a86ae6cee15ac9deee52f94c6c699c0a04fa4afce029c3819066ac4f50b808fcc5c21ce832a3e72d0b7946581;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14b0c183642794dd8bea3dba0184e93151ef9b3bd8bf2c2345a7f32fcef26da8abbe51998ced9d65b85191f10de2669bc34ecc9b01c3afac8846f8242a6d9803a30ca8a6911efef764f190ad207be339dddb5d90cad602c11a0456a9e39f5dcd79b392ec51ef560f131;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19da021e9282364fcf8c34af766ad3bd4629645659f06c03ad77fc3cfdc4efffd3158fdaa2d850debe30e4b2ae3ed0e9b229650993d5d7c4403e3ea9d79d104860925288cf9ed0b90691a86dc11562a2c393cb0b44ca0c7faee539c8a5c7ead3273f70037e9a71f5902;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17eb9c6ac66099e7f0e81e87e8fe8568a3ff81a153452f52810f5291b5e6b4e11eaf2c1d95f4c886c08a9f2d487f3abf64189cd4ee1dda791e339484389e53082f69db70f386a308f23801c58da3cc69f0e6f5d3ca4964af05801341af43e2d3bc6268cae7f8c0a9d94;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hac339d50383a2ad2c60e55dbfbb17aeca1d91a83a4198d2555875e43978ac8cf5310d4b97a76b387bc1ed72b1b0b8ef89e8840659b752468ea52a476c9d8c95317790b126785a47306ade2f63e859dd687b84b2d0491444ef5fdf113285b50ab1d0be53820216b14c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8ba28b615ad0e69d13fbea68105d3d5ff8cce082178cf813c86227f38889538b486b238a897071590fb055b8161a3c5f958a044cc5e0eff93866503c0de76ab06eaa16670a456d74e496363a4152fa033bf4f520d8e034d9c817b6af76807ffa8f626101a3a084284d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a42978b45d6d30b9e8ed8057d799e9435ea435b62aa36c0fe3b3a29a037ebef051b6de6f9b4dac5f4bbe3247824732e30616d1d14f59d27b56c20ad526e318012f9ec2fba3e682537711c29d8e7b195a2751670dc82a41554178ff716757ab52b983aab6487f4e7fd9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h50425fcd2f62094ea74bccd26dc72655230b727021931a9f95a784eeab523319469cafd851a86af6c2e2268abd0f07f2ea822774b8aac14a30adb0b79e000e7bcc801e02905a6597ceeba82862c930991750b681231839514e21b327889479092f16cb99de3f3984ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13caef55d1cc4b15f4c46e614f8dc51d9e48dc6e38092a9f631f30fc85db3642f9f17de53342adc31970aef2c0997e14c2fb6adee5893ba0d037d43e380731a783be73a40d6bd1667d76d1753c76dda2ea887b366ad2a84cd9671dc717fca1c201c610e9803f6ab6bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc64c03fbee83a1d00e905e4fe7ee5c9a2ac3efb4eb05889bb83dad9d4870a3ad70ab15687f8bd9bd89383123a686a1f17ec6b1f5ac18def60c5635da039d9a7560f7f59129dfcac3a4a0c5f41ad4a3161dec302229c55d6bec1af305c63181472385c36b9d5ea7e897;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h91d03086032575d8cc77feff868a0902b9bd7251129f3f0b232afc643760f5b135339c63cba939d9bb708e4df60fc7661f685055e8815087e3bbdd579c07c4982fb5495c0cdaac1f520cea31778ee290fd5d2e9b4d1650f02b165c74bf7d5720d5aba3558a58afa2e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1754334321bb2308031d640fafcdd1c3804fb31d32abc7b6d8eaed85ab471a8d6a493ec1aabdd854fe4aedb3ec848a4b7f854740d848af629c6d64855311e04c7acf5d462afaa736a96a3e0aed5f5e61dfa0e968f840a7ee769151173ddb018cecca8705900877a20;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h65bb7f2e70fed5eb490bc66a988caec9446bd55eb27884bb12fe65e73657a81dddd3874274859cbf9908c657b11385ffce4bcdf40a861e914cf605d84a5578710efdb6cf963f47d128e3d35fc173e94f3ad59c5e973a254733a0ffcad176155ce23bffb3f51eeddffe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h145aca5c9a4c19e90a4981c1f990610b33dd9264e5656d31ce827bfcdf452b3bdf6b5224f775d244c17a81f2a9ca187d7e8f2d40070ab77a030004356fd356ccfc9efa4db75b74aaecf88829aac14b3c772635a8c75238f2603c3e8e98a9b85be9c26ca44071a01c311;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he06caec2be8a050c24e8d9c28520bc7d61bfe8982d60c21a61ad66cf8309728f65971b0191acdb0d6fda3eedd801a59559e2f4bce60b9259e9811d1f3396ffdee147c321d8880ab8876c9f66f42602f5f841ed6564f21e8280979283e534bb69ed0d0dd7ad4bdfdc76;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd965c215b324265ae405d6838e24a95b7945ca59fe1fc755039c94c856c6464c3e6a5f5d87bf873363268afb4c60e4808fc0ef3f29bbb6e76e44b0e3104c9f4251d90564b793fa4d2fec1e55891d1c66d80486e9b560cc22c7df6fc59c79279c7c8d1882e1ee9fb48;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1929589fb6e940882dda932aeb99e995912995d400e31dea32d2dd225abe64128eb1e871925e1989c7a827f2c3020cfa2ae142b8901ef693813ba77dfbada8409328522077a6427babf418b90cf3fec18f2cecbd96907427e15e2a2eeb54900cf56f7dbda74f5af841e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f120453557a0cd4a3e80c11e41b84e89c355d028309efcfb0aa027d076e6b8b8bc8cde2cb9ebe9375744faf2cdec0601499856bcce76577e654eb009ab5f7806731a518e0cf3fa6f6d4a4b1a05cb9acf62ac45af42410edf16061799ca971e1cfc593a943a9f11d93;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83fceedcae12d990cbaaec0906fba62186976dc30b27ba599b2c873a9de2d1cab0550b7afc29cead3065edb87b66dac6a17850fe07673b850457f5b5880ec474d4052eb4d36b0ff03f72b2939009a9c59c6c2ab5e5dacc13b5500cc403c8d56e0712c793a9a227bfb7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d5e1383ebb108a006b7d26f5c509d7858a1f273fbb1761f31281237ba1682b314a9f6046d227141519ffe4e942ad37419112e775a0977bec1383b2aa56e4295b5d9cb40d48e10baa68aaf8d2ce07668e81075729ac3debce1dce17b78763ad54727f4e6fc5d6414d0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c58cc60ce662f0fb0a1700eb81c91e31c4bea32978a6c8136f34e0edc86990c3eaac9f22835a921bd72c25c4948104495ae8c0a1b400c21ad72e9b5b40d9d2700cb6852ccffde0b5c34fd24f0749578d85cba0fab11b7887735c435b4347798a4628c6990fe5555573;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8fb63553a0162543054dfbd3f532def1759c7f5112d4d92908618a85e8abfa8c6aad9621bfb3c2039bcbbd6e7d4d491f9eaff61fa9c2e37d34a732474c2ac774fa20470fb2276d279666f1f289d3b8d029ce8436dd0a3c50da451596616d310c84eff9ab03abbcd475;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161db02c5825f3f0214242b51d8ae14fc7d7342374586c9b70c3e54e22cbec0ec1dd533cf98fec09e5e320908f38c6b9c8155ce8f7456e9eac723b7517251aa33e54ee93ec5a47c9db8521f7b75b66e8e0cc760a6b736c8656cf60fd311a6d9fb4a9a57c974621f1f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4bde6b9b712a7f10fdecd41a11a1c04f8d3f0b73debcd7b4f599d3af3b02ad39d6764f3d0ecf884fe7186cda83336710bb566787f1b82de4f21db8a77b81ab22ebfc953cefc6a3f2d4ad309b0009098c5c37d6897098b5996aefe1873504ab93d273dd1a37cd7a41b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f3aeec8f9cfdd8be6546525d22d3713c41ba9a7b71241161fc4ffa6347f042213daf7e8a8ab6d5f1d22cc9ae4d911f383d55caca3a4d31314e255f621e15a89bbb2f31d3328c0ed508af3df561109171334005e696f8836b83cfceb26519586d7aca010ae990171c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2be305a0f37fa6cb6b3b778ae36dcb29913636917d16f669c9ea6c0724fa355bb5753759e4f427c61b17d71289f2d7cd94e36633aa003fd3428f474a09b5a995f96147714335c1bce5efa6e270c63afeb32613af0e43df2ac543a9e64028c7fa58bb99ab83d5b5efb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a0d3e57a72b1bdfbfdbefdbb8d09c5945f01f28d3f73776bf47de55fc45345bfea5018245e027d2b66644e8914ae93fafc09da8a75ea5e45710d36eec16a5d4cbf1f0b3c2e5e6fa7eacade0f96dc792d3e937ca5829873d466554d1fb4afcf7006a8ed595b15689e5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc786d96f90f690baf3eb973f203af2081824f72500fdf84cf014a30ebd1930763827914b9136308e719c1b27ce564390f5486b52ab08e5528a571c7def8c7b8994c8a26df03d419132a976bde22a06665c0d931ba244a5aed7d8b889fbea4a64ffa18206d86de797df;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1385302ece22b75a82d1862847023ac8e11d85f53815fe9720603365a180472f91d7d32a7cc610e2a68a3b5ba3be19a9fa84805a62a029e7289ce2578d1a28f6132da543c09f4420564ab12e9b093b21370850dcc35dc75b8615fea0bda33cd809b7f45344a3de2dd78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e09bb1d1521a802f9a42e9a14672fbd2ce65a7c2519cf1981763f3c69f89abfb3f4edfe60007566daa10fad8e3fc5609289b1c38615f94c53d78a08b8fd7bb42cd986f84e35bb1c40c4efad74b3ca9cedcd413863981827237cdbf7fb8cc9f5d88b38504953c48c313;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h467cbedf5550a88cec61d097fe139a39b4d07270cc43140b399e37d33545b144d8581f9a9d97f43c60745ba3c19b47f0e29782a3186c93f369a2b1c710f9f7e9e251a9822f58112e11f27e181d617a33972e9f2ff6e96e7cb3d95e2af26903c67d1d9f07cd51087ff9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h438d197edabc3511c471b107390ed6b79f05c234dcbd6f744626c17fd4478d8fe5252eac2bf8b8e3a44e9e1ae31dba01c405c94a595c5f1c030c993a417088cf1feb1df05c99dfea26a794fbe1f5866744072723ff20d4114cdb2fbd48788359b2973bc2dbf464995a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eae1d0f988b91861ceff8d2eaa236311178f8e686d62fe8258433e6939e002bad434442c2ba7b213f9558931294762136db41e3f1505388863df4cbd8ec8af242dbc1d2e846ed997963126aebf3316cb617298074e440a236b6ccc267bb37ca9991d89b8d07a99d0e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15fa82a5ed68e6ec61199a4533a1f42078a07845c825086b55373914e643567895a1459166ea3fa6ada64e80d0471662acb41073be20564a25b0455419f7d481e8070e11086c3e963d225879ca83af242184275e3debd154dd3ef41064408541506cbf5040aa54dec1c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc4d8a98bdec2ce4bebeedb751126fb6e9ef7047061e55fbb9cf5214c216a1ea496b694df82e4e9ce19548870916bd8c1a72b9df80f42ce95e190761b4c81a49bb873c8004d4b7f8a180022a9a2a4f29532105bf9a9ce0e640be9b6f5e90c551809f3b72fabba1cd90;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf9d4a1b600328b67f2f643beb323a2fddc67e3dcdd39b752f097a5c730f2d8947c0b9ef12e070fc9478af13f12061a0fead4c8722da31524db0869be9561ca4b1d055b2b2d218f386f9689fb7ee00179c596ba827deef0c8bc5a2e1d533492d141dd4cd91dbbec918e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d904e46483278c99385c41de31b987429bdc67340eec92cb4a7852f9fea2d490aa5c7fb6726089cde28941ac8618c96a906c04583739df88b1037d3a86914d3824d0117e35d11a0be51fcb123c948a91e70136a60a4267643bebd43c59312a09513528a675a3e6b06a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha7f3d2c29f527bf60d44ed4e0659165adc5a87fbe23bdd603d3a6b95ac6ab4f10573245dfa7e80d46a54ff5dddf7ebe50315a47ffcb3657d7a436b482aae6e9f583a9fee36c8b87d59c0aae048eda5976ef007320031cf8d0d3042cf5a5a4235bbd409c7b6115a814f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f644b4f73c19d6357af670b3a1c5f8c6810ea30f0c7922aebf9bd2f1b6ebd389c890bea0eb2f315b7da26264def73e9baa1aedd93c897d2b27c38780639cc207e80a37f171eee6740d2d6399215945da77dcffa93bd0ebd5e7a09bb7f5593c90ae002267639bdb1e9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hccb16dd0b3bbf70953b1683d14f47f0e56713bfc109228e7e6e4a3aaf4d121105d19a3c0b72aea4e80e99f40246fdff89b79798309df30bef1647d802bc6d315d6aea5c9a513db3404ed4fa4a351ebb11920f259369521d18f15d69e22340e70d8f45856379bdc239e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h262dbf2c7ef6002d64e055787db8aaf6bd329004460494cf6bf6b7ff6da472dd7318db5dffb0632bbd87707a091c61a65ae9b345963c4313ce1c980eba0eb3188ad5990e96a9a3cbe415b7fcb033a557e3be097f7e8b9077a0608279389ca7e391cfec91e62c3b6e25;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8101062b14db4fb6ff1a4f7c0bec184b00c9f23285aed6b6f749d18018eaf5acb21d5805c04a4a9a88e3226e3694836593825346fe01784accecfde49c9e0633b81dd724dfde31a749f4c9cc0efa2a94346b57fcb6cb0989512b60e093d122128236855e5f70dbfceb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2df78a40e5e767b874cc9f16514bf62811e8ea8c4105ed78002c9d26023c5101c07f4fc8fa50b12c73aa328d212d13402b125324acfb83ca4c9ff94f9b6d1948f4c39bff2f6d02c3a9a762816e1f14a29d8cd846c3fdb9a4dedb088d5b854d0a45f981de78bd560dbc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6fa5ca15c7c892b48ef27abc4b61ccff8fd4e1dce1373c64e1949995c98ab36ed9491411f58e878deb466aa79a5cae1b9c979aaa42a1a035f15118f2c56a6709016077d006adbc5084bf6c0fedaf813b50bb4ccc2c1d0031d9a9842834183ce4b5e6a3a486668a917e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17201f2111c2ded094ca9a5b53c3ac0e77ab9d3090310c7f4ae2a0ad8bdc39ae698ec0154c8eebdad7cb9eb7088773c43fec959d553c6e121df05ae2b29e2d7db4c92844001578203748723720a34489d19bae61d6161bcc03ed91d5aafd2d8bbd16cd7959252a24918;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had2d018972fa4666fb3dd8475ac89773bc83a3728832e80232df6d6803163750f9ddea85b0402c311f9dc000fcbcee0c7bcb09c60f552ec777a950df2f6ff640b7de66a93a7295d3da63232d54e3a01442f1f47a3b18dc0e13012571d07893c822e583a04d90c0e85b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h171f268154bb49f6e1ac6a3c6fb2732367e65b74a440bdfba6e38ca2bd4dac8a0d2d48b6a0eadc83f1ae9cabee2e8dd637945cd3b7acc6bd136da8c6875405d54aa61ca464e021d940a975e6e3caf626c3c2865dc8388f6f2e82fb7ca5e9e9acdc45d05f392400aa9b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha64c541d7272877637039d1b46d361d5040bd5b5a358b7ddad852175f4f7d6e977e0af85fb4480e6f450c16bb15c29b6e9538bcf212343cd451d4297e3b46e4a51c1ee90e1c96d1c879ee1555576a4c96c605624b776b8d2b7564243318abec69ba9d8393e8e4e00b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h850ad391b5b7b8a8b83b7e8e33a00074e547b09464e78885b1bfa7c6e4cf4038165e2ea031755b97eaca970631d3eba1a43a2b4ae265f8ef8e8c13b7aa61bdcf1776f155f6a61522d643917c5128b04bef7705cbcedb51aabf19b69d7ff4737c58e062fcd4b63ad70a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1451d8778ec6f1dec321fa0c82b83b7fdb9052c61f044510f4dfef91f72977fb46d2b98ff007d20704329997a2042b1f6673fee6e269af20dcce374654894187c9b773d00b7fe0d58c952b41b55fc1f310e7e97bf497afd5440eb996d93625ff95efa4fc8943c487532;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc812c4eee5427b417c3b06547e13eb835b9a75dcd2bc6f2566633f5a22e2a7bb4084c6cd1c132bca457236ea8f1012869fd819404d070e1457fa79f240f4a703347a48050ca0d501ffb227042f366c4579e7b9f4cf3c4b5642aff7785d2358ade172860f38e2cb8f21;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a55335b959467f85555ca713f6e9717dfec87ff87bb9a6d0e305c018a04545f9ba76827860b0e2465b48c10b57de2eb931816a956356d766050d1598fde903069d242fd2d6d1e40384e807edc8136242179ff287e172eb804de930dca65d1f0c15dc93a4c31cf9791;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14f2e5c0a298cc90c66acef5c39850dae065b5ab9da373a05629cc04c043d54b143a99364821811138b87c32b37ddcbc5d4fba845e10b2f46b38d8ef4efb417f945347871af43762d1cdcc4ed0c19fb6d2afbef77803729abb799bfc72be4d07b044fc0207aa54ac41;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c571b74262fc9c110d3ebf9f259aec77761f2506090295950cc2345c1905016eb4766e1ed4851965d2610559030ce45c1d6c99f8fe40f47b9ad197f8c54e2d25a537e4896b5e838e2f63981ac68e254a9f75ec0a42f1ad270e9c41f30af5a0eae7822ccb40fcf472b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0d414ff459717766115e95696844bbbb8a57d0147a1c70071a390c2ffc12697faf1140d0ab876a8989ae69abf433c9ed7092290846a259e2d12ad5c885d7e293eef58efeeb720ba1ad72fba557be34edee7c2f222a6a2cc04c8b5721b571da6fa86a4e120c7375a1f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd572f33ff54d598a1848dc42dca4826006224c88600b990a571b1ee18af5f25233849529d9ad9129213924bafc27fa742f58914d861573fba8e316ab95a98f3e4feb5fbcdcaf0c879ea0a6f592f93b2d38c9cf17f64357dba99979799deb8e1503931625c24d086aa7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147d21346b6ea663dcd5db5cdfa304e32bea0221083476262f0b5a6dd03ee8b6c08edf420ad228c8b731530f50fa263989c026cd169de05a16f17050fda301a020430afad1af559de9c97fcd5949abfd5c634f2ac040a5db69b5ca028106e2e80143c43956f1b21b798;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13a59373ae5cf0407a1ffae59a7c8de4ef84f0cbc851e1532f956268666964602872cc730a0e42bc27a30a5ce43c876d0a693c621101b15a63cf20ff02a4641d33b71088319c6a9f9222d0af69d71a4d00d3f7ad8d1940a103b91a9f1e0ec70874f246f99a69837d56a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11fcfacbc557b510ea9c7bbe9cf8079e586fcbdff530f6057b29a822eaad5d3e0ad323501b2e819e527dc2ee45ce59bb0fe4caf619895202fc516c40806382c4f1e6297401074cc23391f996b32868bd03b111a8706f2b141f02fd0367aa4cc736c2bf9f5c89a488d17;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a83b0d77a0b4a372581a320716452eec557f1ef99f757f364e950f9440aa73a1bc9e7ccc295a22b2b4780f9a498b591f981e6556eb9071e53d56924ae3bcca9863d652b9c5921b027cfeb2b027ecef93c9d58c6917a012a282add2d782659404bbcc3b1658f7214f2b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bfcbd6a42896732d56c63de537aa8c9fdf1d17615d2023de1da4f4b7de763f211710a69b2d09e4e089c805d55cb92ff624c591e5ae75c34e2b96030de36e1aacb59f54763b316ae721cef641ec241f34e4ebe019884abb66b1ba8958bac8f80666a94cda6d0728856f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee8c22e6a00411980ecffb51c069c5685015d8de97d79f015bb21dfc9d7529afb0e854c3209488d75fd3e7c207d256c86ef8c686dd00ba38c832313887de73734715fbca9fd7adfb071f43539781f5e678c671c8c7e8b3765fbc4192f68fbd3e0537732a46daa72e5b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h175d0f059de92f3c22d168fb2e18fb5b45547cd92372fe8ae56b136c1ed9fd84c20f8ea3585b3141d4df9ac4147f7c9df0348411478e3639afe0636b5ebdcff27e21964293f880b365fca4bc146a9a273fcc3a8ada90876f066473409a685def9cbc0683b0a2ee97a2c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hacb1403b0171b3f86b75b6817313c9a7c26b09fa69f18d114e7bf81365fcb4483beba33a79b398e78fa341e1067b5425b58b8b4151691064761287a157ee33d756fefb9afd6680421aacbc4e9db2ba027d4d2c79897775d9589c1f3ae5273de5e3355956cbfc914516;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd63a410e52d5b5c8f0dc4cd39b27d0d42717ffa1e4f5f57bd617f55360428ccd2ba53d719cf7ed071d09c5d85233d38c114fd5c07b6564ae98af873fcb60da00e43e688934fc830b1f0d51bca952b425c7cd7ec8e716e17bd58251d8f2a0546ec07c003008db4cc1a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f85c430e6bf8533a3aadf3bfec6a0704dd725d9c23c5e903497cd79cf4d5bda9dedc0c84b194acbb936d1737e8c55ce2a454df4786ff7f3ea463bbc2ff7a17b10205b3c258885aa7bb4db4d53c7d634f4e99fbd248897c5379b9d46319c9d59034ac93846fc54b73cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f7e2101e0deea8f71f0bf1d67c3b26a8241ef4156886d7d565429bc71765091bc893746baab9a1c4f65fd789c5c7d5fc64cad8ef8811ad78fcd6c63fae74ffa7ee87eb3d98dcf5280088298e6cb807fa0ad63059426260572d847ce0c00e54a8e413e3ddc3f6c19ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db0d530b0f394525bee2f5961d4c9f00c73a3e2f8ecdfbfa91222a2f2ae87df439e3f3eaec81034a3205649f2c48bb881bf83a7bf5e8d53bcd82d6f6f448d8979fb5ada4929f2ed7a4d9af1db4d23c27b75bfef6fd7efa897bb2db5f0051a11633168f634bed6e0ee0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9cf50f919ff6bac052efbc06494db6f1378c862d5b2ed336f6b89c52a45f3e97be6e3289667fa9e493c21890b548bc8f2b3c2e32fac7f3596b55e2071ccfcb73e619e29cce86a313026756a85c47a13eeeb2035065ae95e1f9e7fb6054a4f8f213feed21a936858088;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1737797f7f1d998727e6f53c7c9c5563ed2fddd6a31092fe2d9002da629a0acc49b1ce2229a9fe5e115df038a17af09c0950ac90989a041807ef157a807f5897071b53401171777bcb1da0a38a30f1f48730d398a5518e7ddbb861cd4c636fcc502aa3f465877dc0914;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5993e1d00d867d6dbf61eba900e3f6c375e3894bad8dc98b4be63a0065668c3cf8f939f84e93ab3fdfc3e1181ea7f12133d5b0352e8040a62d623a24f1cc21a495528bccb39fe4e377dcf6744d93336cff8e8dedcd9a1dfac028da35ffe4d29433442dfbaa8038af71;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h111b2e9fe036d3ff483c9a90d4635d6ff9dce6920a715856e5e55271d831604be394b1cd20a7052494bdc9e79c9753db9f9584951a4d9418f7d2cdce7b36706a836998f18c9d612de91f3bf2fcdcfe2a71800034e1a6860caabcb1832011f58e347af868fe80e4336ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18f25f5b16e0dae693797a7f77b2fd91a09db02a35e3fdc054c65eb309de093670ad016de885d8e5fb5222611b52f55b45f57ab2cec1c685d2e7f9c1131baa064eb30e4ec37069c1317cee318b75eb4ee5616ec0b9a91bcc482bc0c962ff53de45d7b39422d90df96a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12f73518f2d36ee300b7acd9ccde183abe8611a0393a78523dc994358fab66f9279f8876fbcd66909021efa75ac0c569266768f4382ee638439d4bdb7aa7c7bc8edd529095e4017125a2e286be1e86beae8020758d88a9338e9a913309e8ab5f31b1dd3ee36510cb4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f5210d849dde3d7decd4f799fec13beecfcf364b9987fcbf7e0b4535c390216f398e1d8e056b4a6249cd5d8f25294e1e559db4139eb9558c8b43eff1e5c293fe95568f22607e25698503850e205514455fb85d4ab00c83bc562691e6e7331bb6e3c0f666474291f97;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h164f54e5c4aa852bb06f1b68fe0efd7659d43536bc4c7dcd952bf7e2fc2b900fc07ec0db5cf7470b1cf597a7a267b7404e70805c08a4a7f9bdab35f1c181b39817866a93f6e998221ba2cc9281b36a627a72f15019828f66cfae89555f62831e5a9583be2986b886676;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h153216bcfb46a6e6106737aeef37f8a3c810ba003d4d22af550495d231a0a1305abd052c63b662eae739c11d9f39752861a43b5a3f3afae1bebc24fcc3b9aa624c7f9689962b7930c6a82c178b5b5a4784dc2a3fb6631bd261cb9f9a1d069485fafe61f4294be0f8c35;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1302d19ff348a16af693444690e89ffa7697245dfce62ee292e744ffad9b3896c97651979178e78c9b32db21dfaa9feb9d14a4a347fa7649e055de4c77748f4c75a11794ab219189e22b3d844e8f9631feacb0216f3edad37e3d20ff897748475d78a6341eaf4678e9c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b6c075191687f5e8ba38f10df8fd2d5e7f62700ffa550ca5839793bba3aac7570c151315620543c6c2ef93baf15843a3aeb1d611e6185e8716a04d1aa5b0be8b01c1e8083cca0ac550e2787c496ced9f3ea4c6c5a77433821266d0dec279cf37d88c368f4e38ef883d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc698737e3a44747283d7dbefc30c2ed398e2dcec05536cfb83c9c9ae0a328f920dc3f0e8ed41b6ea9562856e9cce9b9be3a85811f0e31a3d235ac1f26cb2bc4550acb1ceceb91c58e4e2d2c86ce2a766587057ef8d12396610956347803c9aaddbbdbba48fcd3667db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h50f60fd4761250d1eb96b94d9d40c91f1ceb51e1fb223f5353288f8ee18e791bdcc98c1687f8b776f66ebf5ca1fb41bd3e46d1c966f308ecefe8f5d3a00c6e4ee2df26f1f69d6a3f3dd6ce1079d13d05883362b689d82077ea4bde3ad10a737e142faea9965dc9d3f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16abdcd5830cb6b6f4407e7c46545f19a6259c3617f0fe83199b09d2693b7d12204faa8a749f9bd0290d9329243a177dc12fb9c90d37444084553652a4c24f7decf21528f705097300b354f935ffaac2c56ffeb5a4ed894c8976cac5e10b35759f0e7b8f34ff5f96e47;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h109acc3860e31c03195fa9d45a038c5351aa3a842f7ffed34e3510542dcc050652860e608eb22a98e3048ba857aa9fbcd12da7e2ddf4c2caaa91673275488216aa464aebd1a0395d94cd401a78dbcfe173d571b3ad2c7d580da0f48b145aef310f72d3d524985116b8d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b4485a5203cf6a7554398a3073c6d196c592319b611571b670236ffadc56b1d6407bb7f63fc206f968cbbce9cc84384146dca2c1c0e0c730e90a60c8a9ed604c667d666a342ac3efd3dc34aa04d8fd5fd08d1c3e2ac026c7908f8c9db61309b3b8c5e945941f105cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a3cdacdf7b1df9b18fec2031f6bdfa8d7083a060feede2858ff8339a243942cabad0cb4a76d188bb75d0c8cc69e8a429b3d5febdeea47c114eed704c58e72ae94076df9abdbf85cfc876e0e5c027bc6e71746dcb17b92444c1a14bf6394eaae41894bf295ca848a22;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha2a2bc6d9a18a11af149af4d26664dc757476ba5574c4a7e45fdb61785bb108df51c0110afbf16033fcb4bb9e4b2ebb585c106375b91f27bf06f6bcbd5b4a74a172a7587260d609ac55f97c30b596e3023332c53df46f34c23c15f90e37a417d6e5d91a0dc8fdd3f1a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c398d061e49be70d751bbee4b7999ba43c60582e80cb61a0ff35f3abdb57eb55d4d64f7b44cb674969dbb06c6cc3b9f7855d73882f669f7ed86cf285358dcd5b86921c415411769888fb245e884fa91d7283fb9f0d9b23f7b0157935135394f5eed2c229cdd09f03f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfb1ff0586e92a3c7d730bb77d678fb37cf30466548c3eb77baa74fa45abadbcc50d50d7a059ca6d09c8f96a96513e957161324c802a866f2836a48c700ae537bc0bbc875d444ae91ea7f16f2287de55732e94130a8c88b53fb266cf310ed8dfd0b35537b3cd2a74f18;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15dbc4ac7ffaf0cdfd838e2d2da4471630d1f17fd88a04d5f5e58fc01025c93846da714b79d646f4fb775f2484405b53304560a83e7d1ec98895a91262d75b0ada009f92c68c303cc9860bf258e7477e99b5ee260796462979c5bbafdbf2499e2285c9a9aa24e3cd6f8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ce63eb5a304c56aa2b1d0352123ebfb59486da71964e1725417210154b8c2bba24cbe764093d29e820f3bef6bcc73c81a842c859b9d272c87c552728155c4c93a7b02e5967e86dea8ec5e52e752dbb6dcc1831446b121fb593f95ce62f4f487873ee24bc57c122a30;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8d3532ea53dedff695d53dfd9211f13c77b1697438da76087bf8bae602a4201c1cb7ce83c2e020a2e4c0cca329c31f18d9ccb2190da1664442ab89c4325dd3b7bba8d571427573d29c8f8d0f1a99c6c0cc3e6c72e7b2827e9ea90aaf8e2f16b136c212fbcd01bb02f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc1bd4d04ebc1409da835491d6217632dc996a54e7ca560d9b4399eb6d2189436d79b0530a6fe654781d0ccb277f8ef27dc90acfc31849baf88c19e28c12f1a3658cae1ecc3b92aae1578577503b258f5b072099f9d1ea70d49f9099c8039957e38a79b485707c08bcc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15719307ce8065a9f4a149f2221b419a3aaa958afe073cc6a50286ac1a710179368964ee33f01cf06b96d10f71530b9682a4d2464bf522a0e1e6cefccb81e83954e98217939e1af4fe97935e2e19048251e6763f00374a071610edb20f162c26d87d4986258ea2c56a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c79034b664df53964e0212dffb38557c1061a17853b99e12641ef3f7dbe3a4355d2683ef075c222462b8b1e716a012aa7c9e7acec9eb64bc5600aff0a9c6d7603543ee344753aa6c13e2106cfdd8ae3e7e726e3b21e261317a2850c27ad05b82e0de4bfcf76287120;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h379bd9a574e52f2f7c31909327773b10c2a808eefd89783a49fdee0a5740ed1d9f6c45e3624e75b4ff74091ca596d20e609a65d8d37516df83e5c8da30489a1abdc27b6a5a18587e030bf58ec3f2f145aab50aa4f2029382fa5f70cc2e80c9a6f045fc865d26caba82;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1495ea1b3c02b4307bb7e95fda81278ea08758cf56b291eb004216e0e01e9af9da5f2746bd0fb2a3d170e4715d13375595a963c44d7ef2f187759c4dc0acdc09f200fab7fced30dd8ed5274c465f385ca5187fe8de798c3c7ea56973eaf759d354ca469a55374725669;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h31fffed372af8411523dcff4682347a96fd0dfa39a45342961bfefc514b99d62a3e1127c386c5194a3a876f51ae7c3a749bfc59e18f6210fe834dd5f66aad6963a240e9b6bf556c28c7abe6eb21dc6558464d6a86a529b15fe19207dc2270fb7444321ead32ae003ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h105f755d314d85da3a90a1d60a05d7f6675750c602f5b1d081d4e5b6a0eb05c0fad0fc85f6cf433936158694589e24087991f595d7eab6a6873025ce62014eac1868f79aacf082734abb4ab5a3db736dadce9d639750e272607d26aea27094c4a0c72ce493f8f121497;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ffc55a597742fff53c240c6b36455e25d0d186355e011327cd46b015e177d522fead47c99f905886c8ab9aef7517222ceb10aa5b18a0d30c77b2ae7e20e4499a9267be7e51bb0f21969c128aa6f804b5ee74df866444c510a4dd33c95e591e175527b1e0b6906bfe4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ea175bece5aa70e97f0dc8e6f4e50f49258b6beb6e84040e03e7a5aec68feb039fda9be9f1407d0af8760e47989c7d7f49552bd63d4c1bc2924d6a6b25ab9f2ca5bc2e719ca264645ebc9ca11f97812fdafbe8ab77c3e8718d80c8501550d5972a5fc25b93cb394fc1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7c1cef1a3a91f908df2e09f58444f2898bf6b5e7fc5f60e91d156574e59e28d5c1ba34cfad9c83e2428db0850f0d17c77fd56713da147743297753860a9c24e7a6803830b59627648ea5b2b9ac995494c3fbf5f677ac2a812b25355bf02cd0f3572a13231d0b0b2be8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h191b9203de2caeb0c4ac8a33fc996372f8c36d0bb0fb3cc8bab202ea0972ea53c0547afcca1e41486066fb29d63e102129aafc7c24d29d1d454b9f3e44df9070d40c5e040446d963d2ad7cf557b716ce764aa4c1c3d8e87bf19ad1bded729191118db17dba562e7fa38;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c0bec2e8219b19351d8ef30839423ff9ea6885c97b0099145f831b42d53127b1fb7b8eee586232da475733c232f268effd90279520a29128c7c804e087ba3d2efe02674d9caf94bdc8f01e8fae52e174d328acc27a8c0cba32f5f3d19cc8ff9245f6858b838103a36;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8361965c6546954a2cd5b6f6d956819a320eaf86db2138487ea401cdf0e3669ba9f5e5d655730950c52647094a1d1e50deddef54bb3054292425131dec6de24809f2abd95a675b9a30f0e8a33fed821002c41304ba108a490895a5ef5c0417facb1d868808d9163290;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c1cd731186b635ae64a19716d662638cc4abf81f622293c7ef4f0a69b857ff14ea6f22bd3f1ebf0a22c913ed0fd1ec11f2798b6ed52648a7ab356637c0191bd2dbdcea91064472922ff3646a38b607310fe8df674504478749b6f3db773123abf5380ac65fce46fbb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13c44a49815bba733582a1fb0be39c15eb7a1ba2d7140c8d95190d6dbc22b8f0ad1fe8017e6cab2f4cc4a77216cf10f7c7bcebc70e0f7715276e84e0904c5a47c60d053b2b2c393299e42d1d220c7c63bd51123a4bd5f2737d2600a0dac13b28b356063beaa81f6e397;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b476a02dbce2835d02d35b3f149950e5b42100628e14cdf0c235154666494dbfe5a7d2a807c3bb31e485e723c4363b918276dc23cb8a63e75cf6b845c86621ed2611804160424a9e821bdbc1440769afdfdc7904f84686b26119f35dab8951095a5c35c3ece482762;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb00f1f4cab1dae920ea4f3d2b74b87e040d90b2bdc2483d4e95157234eba41501c42169ce7b2042ef831498a9f6d7752c574d0e30c3678f0e0f8df5cf3e4071675a9a02a22049384e157a727c39cea21d8edecd92396addd8b47ae7a162f55389993348f3210db2247;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f29c9c9d707e8b427f55707ae511f4a9d7054a4b8a1efc71f4402a7cd821c49d332b4bedc720c37d16e2803696a68a9ac6628426ce55548ff37e19629f5dc979eb29bdd25adaccf14861b83d575c9bc9881cb175a77df04bc54b276c0dbbf3d98178eb365e24bae4dc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h30ccc012fd6a08e170579a774cc0ef212c4a65a974980d9a9d50671f2d25ecffd202834c47339a1234b4e7aa9d63805baf8b81090c622f04274cebaed6af51c07ac25565168bada9fb06f1fd815c8840594758f052bd2275d77f5bf03bc3b220bb2e7bf03a699fb70a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he5fa91329877cae3e2c30008b5b948dd1a0f88a25c86be306b2a872ce515b64de2cb81e3cea4444af81a5a73709b1ab25806d013057acbe7871d51958a5419e8414592ef4e84a28065488f5ca726effc52284dc40fd7f20ac24d0e5129158f71d18a762f9789956ac5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100a5b3cd361d95e9de0fa4a14abd9b230d25763b92574a74df2b387ca9d9176c48e0a18a884c4256a3a77933ffef0df623d871a37e7c3b251e865540e4a87f207e5ea39596e707eef115eb2b8abcb459e49c18400733be012a99109275724da6812334f2cdaade9bd1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1673632ecc564fc6d7ed21f792d241e351be54a2e603338fa79f5e7fbca63b478e5424fc358190fcc665402f0dbfd149e4382256eac261b9a73a950eab0737f0a5e8abac84776d6c78b3f0a34a816e44615bc72bdaacdddc2f50ff988da380c974f0d14487be09f4e75;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1048e6215866956394fd9d5d229d9e054b60ade6c3be4658987fc9de43b9dc931161b0bc0db39f7a59ff13c8f9ec555299955c99d3ff5089b66cb9850647d950603cd86ec332f3a1af408b8e2af79301617619f05841db99573b6ea69e122c4cd4adceccc362ad8fad2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h168256255dbd93b2c1456e67dc906e8961cba246685031e084f5239164e2c14913560dbed3b7125ca4e676a808dca96679ee0c681ecd58a4b8c69364315820303c5ecdaa3385f563aa4d078f7bf2d30e667322094a027e6ac3729de03214b535e40decb70df9f3dd660;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbb08d57aa0da33dbe08ae02ff5abd0c6085be41b49343a3f16e31f5e6fd1c588d8f5bc3f27d049c928148a3540eec7ce4dc1a2de39d5612b9e81d10d97607fe060c4bf2e01f956828272cd344198e98bb965ec78e7e18d41d9e1a871ba4573ff74bf271587195547dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h91b1bae409a57c661d0c9390a6882e68591fe758bc1729c90bb91393c51ac967e465b42f36f23e930e272f5a020d995d208be7fb9d54c63f8efc60a450593ffe4645463a1bc4e6610663140d54ced4e6d93fbd5bfeb95004f6a11b3a4fd41363b7aa368dd151189c49;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2e069d63e39d6596690c219f65be86ca621b6f7afb242fbe709f2b28273defe6084af3750081308b772b47313b46a5398ec0cd7a72eeb6fe639a646ac614c60078ce90dfb25e361a315e29540ca01ef25de71a2f2fa4541f8e0ca7c9922c7537c4bd7745e2d1f4206;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38210571e82ffc9e91a8452cfaeec23438f0f6b83441bf8fd20e1a992cc92e13cb3abf8996df135d1ef955a8271d64cbd2c54dcb9e00d456038d1b3eaa4164035f52aa4e3eb0a4b4470b4b7b60a61943e6f51adbfc5485f50b4418525db9681b9c1239c1b5bd1491a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcff492642e55e22275d9a7891a21c8b6022aacc6636dec54f960640e1c888f7d8eec28966000ecb6a543d42eb336ebececd826dcec177d96fcc0053e920824884897f8c509344f0dd6977b3f5635ae5e07415a38c8cd6f87622c9211a905f8f111954040346699910e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h88c2e336fccf7e5111e42e7a635ebc7365bf8962b3abd41d220ae4698c6d7359538cadd128386c1d6b4d2e0ea6d10f0eadf194d9803d1a292b5a0deb982436499e6dbac727eb5d5acd349d8ff4b80a708599bd1d7193f79144c10378cfdbbf81d8c5ee1ff1e743b077;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca5328e1525400f6a5519b345f5421c5e4a455006c4cb811b4888fac3c1b4c93487df45f44937246c8d27692b7ae2d4bdde40fcafd25a233a76ba1a18026b83606e3c54f4a22ac43b0556d39d4e1187ae81cf123fcb1297cc053637b1094b44ed9fcc89e7586dc3953;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7895032297d9f851effe0bc8d33c4cc59d207537ae7e46b89d163971a88b5e8c16b0e5894c6031d2edd397593fae1775cd323596c69c0ce866ffa47b7958f7de23d0be08712d7dda3fb7db9365faffb628e043ca459a895cbd53e5a558e2b9c8a352a221427137f73a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haf69d89ec872dfc10942ca41b0f36c76c9c466d026be62fe15c060c2ab2b221e0d2a5e21d762b4b2f45b4f5691c840c2bcc7da021db0562ae16bee3a8324d618c913eecce745d35cd34d283e13ec012846bbbe00e7d53737e06bee9f278a0d412c257da3dda19e9fb0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38d58137bea25a1c1cbc2aeb6c58da7d4190d40de3bb68444a57c4e1f3136fb13befc477bc66f1ee0583944e9def98ec0737c9614650b98f5c02440600349bda09dbc88829c4a22b3fadfaf56e7daed597d52f9875f27da3162b1c0c2ab5cc672189b0b1937979a89f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4a9c37e6b030f2ba92ec2dd79c5487cecba5865a672b0b923650acedc6ca63df5d102762288e8dc9c4af22478c47c7c37dd53d6520817ab60588ccfbe3c5af38b636a42cf5e72641339c89dae76579f2eb425d2fcf37e3c9fa78784db9d9f1c9d25c11c1250f3dbcb8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he7414f18da0805e7039d49c230a46a29ce53d029a0c7c0aac2c9eb40657423e7e3b7907ecbcabb619f99bfb3f9b3a63e74ca8c411cedf8158e07e1663f018a3568bede06bd232c0f2b6d15a74e12b683dab81df422fa459a6759aec9e1254de285026b072644909c2c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4bde14f101aefd37879c0784af3c536836fcca668863c9825b5331a5be1517b6f2faf97dc51f2e2f0f6066a625051a7c4a1e017cc1b7b819b55de10b6d33cb195a7593100ad1825d0b195b04a0517604b61ca8cdcdcbe8d46c838c94637ca1e62467dd15239c0fffb5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee3af41eccbeea4a7350dcebbdc7781a75d760c697164f0532b951e1ee54d429ba60ec1beeed70ef40733ef0c6fc48e7d4275e3c34a9234f6cce777b86570a163fb4ab024f8d07b6cf98aca44dd786cfe10f000085b8aa2ad68653e496dc4f78bd9f2a0748176db2ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf87f2e2b5e91cae1a13a2182c7e1541fd5984a9dce4883871d8e4cf85d82c36743a65b1d549243680b7f08dd74a7e5d84bbcb2522920aa8021065c07f9d9def92f621a708f3f49365b2aae6c0b859ca7f02f555fabd149a5f04db067e451e5c3d220da3c51b9bb39ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9ae8644f5708b9f0ada3e20c1bd7dd2e6a772b84f87e207747f074372e2da86767f52bf70794c10ff0850afda3f4485055124e80f042f797f4467ab401d38832ae6c5fe21995e16ec78c1927caaaccb0fcdd9486b2d2611a01e2af93f613a0d0e9e48a4f0e79f83335;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e058274fd013777eaf434600763ebb2301a77a3780cf130e4eae8cd67f0c7e5303e8cdf3170b3623593cfb9bba811873a112d6f1722c4bebe96f583d535b3265855f0de9b6193b35c33b90d5fc078bb9eefe31015824c010daddaf40b37603350815d34d81523d7d3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0c3308f82d1fefbf74c69f955299b5bdf8c09898f43a2dd687a355d9143c1f7bddccdb354f0b50ed626fc743bf010bb5ee9db1a2b0dbeaa4217411a5aaddea04555a6c412889c7babd2bd2f71a96b0cf5bb112bbd8dba18857dd5d5151774462d7571abf6b2ff3c21;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141ba6de0a59784e2ba5ca3c6053c793889b4a30126313cc69efd00af83c23a4a8d596d82b7dc83f6954276877f5e611d945f539515a8aa2966dacea30ad11b7973cebe7f37f1848904e8ec52f2df57e609663f7b1c891ef68d1c62622d259da2c03fb86054116c691d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4da23af6b1777719bb72ce01854dc4e2c415159e3955fa184c1a7608550f32c2d8aade2a1e8872424d25fbf0013140d01ba751b33a238b7655b6b0d0ef574b0291aa02d587584c177b1d75826d6d725074967decb89e2d6e146d5619cf7967a3ff8232781f3a17836;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h49a6e739fb96db022f43c380fc1c82c338416cedf043990e18fcab87517b66d231b323f074ef1175503365705c8031382b58fb5df2bd6d5aaa5a36c354fba518886057fa0f0e45a9a87a74e1f7c080c76679f3a934a68c528166f5cf03030d39f9ba9f566ae3ee73b5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe96e9a286efa7f86d9243034f39113bd9a308fe98199fc94bb27679a0ebdfea215b335b1be546768b9954e68052aabd847d891a1318e527c7f051d2c115d4e7db91d79a7d43a76754998a72b8985f1686a8eedbf780e3dbebe968fb904b6fdf8f81c1cd1f0d230592;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1010a87bd2a589ada850ea699e03a3a2ef0b7dc59462564f6882c426e20cbef32a638895ca002c3c6cab8e96f27862e512ffa10b6547f96b267612b32c0a5c44ec9e61ed406994ccf1c2ac2015ed8e71c196b88f67480e90577fc4e5940922b5cfa1eb45fc75e6ca91f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h94af82f9cbd3252210b5b450fbea26b209a9d45200455eecca2d8920b8b76668f462b5b9af200337e2a854c64fccfd1e139d6f4be56ab73ede5c20b2b433c441fe5f1cd6979c91fb2b262a61f269abab461c1f39f8f00ca3ce2e55bef1ea30a4e6f59a9daebc13a60a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1f6974f76641d6992de16144ec96ec4245a3e8882c14fd020e5b092a36354548dd165fa0a6eb2db3bac50da8418a3be7061bb2c160223ae392e300bd6b0ca9345c163162605c8ea51509bb7340eae23ab180953e4b7d631fafcc333ea4891c7130027c80e6d7f61b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5fa9e017b032ce67fe4844887d8b308002b7f85ffc81153e87301c23958669439f0374d3b103605657b5d0e8885079a9216a89e8471f69c2afc358671c269f57ca26abbc90ff8ed0d3b3d04d2eca939e7eb7ebcd81f7a008af5e2dfbe52471c315259ec5784ab1d92a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14bed185a161d900e349e330d96ce826daecf63063ba32400da9d3cc936d0b83aab01dabec2fed5c752b362a7cf030708179e058def0e7c51e94648c30eb7f23d8d6cef6aa90f1989ee69cee2cc34ce8d1ca4bb92920359895beefe7d7c11152ab1af15d8e8c49ea5a8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h935b6cba19396ce883bd2f3cb3e524132cbaa5ddd023cb61806f28ae23b659a3a5304b4ada3f4662cc2a5ca083549311fe190ab1f173f1335963a648f1b52684a97147fc07256bee6754e2a2c13b871f6de41c437a31010d77e2d89d0470845596db98bc0fa3e296ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11c06dbea63062b79fcd919e718e9ae2f6c2b0449e8eb2e9ddb7031b13ee9ac896a45ec9286ed83a42f9b166a4b88a94af8c90da863602cc8db2bdc7d2421da483955a15a25992dd0eeb11469368c3cbd91fbaee7c3d267c55a49c1f33c28a889987c63c7c4cfcca98f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1804ce00893458a14e521f0d05cadf16083f206dbd2693ef2888267c10da7cea955ee2056cabf63baa902e1e3b9010cab8d9d46d492021397a1af7e329e4073207d74a30c65494e22f8a97aaaf37b8e47f206c97358e6bd24357624c09ae5805c88ad54df922ebfca3b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af9f7619e76edde11e60229a586dbe689d19d11b8e50e6cb5a218ab71495fe257ee149d22a729a61fe3406db0ad72e84ecb2fe3e8e8ba12742064172eecc5b623e8614d254df05f813b46b5205488a4561de44139e23caedd1ab7bc2b58a8e7ab917f6a16b7bf942fb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4a59cf0f0b6b74542f2ce458008213f4d8fcf5cbc2e82ec97f3c0e7ed847f86cfc650413e573dfb06626292569859a5a738258346e0f1cf9f3ae3e7e34b2a3edc9fbc9fb55510d30d0c2478148819812d4c328bff873835fdac3f4ecba19ebc9b02fd57ae8366d4132;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e616cb8a0e9f0b2b27756076b600ec757c5a340b4f6e3564c25500a1b41716202d83db262f01259f00defe217e6a902b15e9407e5824681921450c9f54f1b938eb8a5467e18abeb611a4d0b6a73852dfb66ddf714eb3364d84ac8e9e07fa55573352794d0783b10365;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8d5578dfdb8e3027548e3fab0e89558bb3fcd784c9e81eb06f1b72aa41aa0002116aefcd97de0a5ccc8fa04159e2b17e6cabfb56d79f7b26d3dfe11ef48600b64bf6d0faa7f3f2ef8f9efe6c31801ba2e24f05a70a62e3d31e82dcd070e56d230ae598f165fafc54c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h73f80a7c4af022ccefe173102b16f85e608619e2675323dae4db490cb37cdfc1d7ff8a9ea3efa07311b9010a806f36f77d30bee439e202e59a16cd181b7d8dff6b216be06480d2808ea96fe69dcafb3e66ce433ca3123c0d2418e7a86bbf91f8899f60b69a32843bb5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h184a8533e46e1a40194d70161093e8aa31c7110d834fcb773869adf5ac90d9eecd328cb7e7c953ee9755bee04106e58da0bcb9ce93dfdca3df2e35f9bdc4723e58b215107c05484c10681eeb0dc772c1a95659f359cef24398795001929d0e86286e0593a47f04f0785;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150d8074bd72dc5b89128c161272beb68b9d359c5a4304742b1ad2d36a7eb7d656658cb47e350f0c76995cda3f09ab1862f18f6c3ef4f5ee514e447e4434d6d608168181e0600e514fa996eaf49230bbe510da6691dcc6baf75a68a09233a2d7a2eda8b3aaf7fbfd54a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2e2a61836ec8a6eb77904456c716b4849b26fd49167a16dea4b76f71212912a02025f3e1ec40e7fa091a532424435ba6e085ef31f8da7aced143b0082180823b1922d81679f5c98753c359a19e61c880653f5fb4f3fdd230dfe58f8bf6264740649105a48a6a6593eb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d7c1c8413b2ae5cb845153d602dab5e4c4706cd40981d9322b637c2f48086bbf29322dac6d52905a8d937fb659ce2dcad6920ae18afd546ce754449c40125182c740d7f1a19c2fcb27673af93120c837905171d34aa5bdbf0d96cbd58a9e30b18a1c0b4e63c65bd9f1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h199d4769d69fbbb2d36dfccfd91c9091f23a43d827be08b0357b73f2a66825e09e29a22df521537bb95a4c23965ec1b74a6cbb8a9cd9e0582bbbb17c5989a3f5301f6ff806362b06ef55d26416cc34aed821e611b8967c3f535ec8aede734e71355fed7e2abe03863b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ce4054ea7ef58b5ebc90e995637544e16295ccb268c36c92847d05e0cfbda1f8e801a5f00ee2312227e300298c5bcd196fdf71d9b946f7d3b66df32e6184fa0910f0519305411427e71a74879b068569043fe8655c030e08e9f66280888c0db7462029817ad38071f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1516f1f12ffe36b717cde062b436e4d00f9ed282725d07045b79a12196bd4b761730823a5404d9651e3e5717ed9e8e417e141192350d9c36949c402f5cad32c5892b6da5f878289165cfc0589969a9403b8c69ec3112e5f64be67cac0e6562157803a2451dd2d6cccd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec3090a051fba66bd1e15d4cd1ae4260f91de45658ddb0f6b8aebd2ebf16765a87d6bc94816f8038ece956896f5afcd99b44dab64627297576644ddcdc0a54febc20048ef12ab45ddb273f48deabb9b189893d7b5ad6180863f74916e32f72fbb3b220083102f5af98;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hded8653c65d70c51ce0cbd94e3feb5f04a66c40012bc59eccb86017b8bec47bf3c3ba3884067235d132bdbd04f0da470ffc30448b063b98849d71a1025744d8f7e6a53c96d2890b2c52866c3cbce1edeb7840b399dcc7053e71b88a644fb21e4f9e7633297c0cc62ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h767293560785b56f6155ce480ce61c7c5df3564f989207811c7dff6a686d36b40cc5cc398dbee4da1a9a54f6cf5a8677afe82ff20b16ef3d2a4469c2207e2ac097c572135aaf1b7e66148f7eec006b42b288b546e697a21ad65c98eaa8929d448f6685f6ed394e586e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122cdcd46a35650fe46550f88c3f79803ffb867cf1d82d78139eb5770ec22ab69f81327a5cb99fa18fef03ba2c42134db105b0f9d03943879407591bb025009bc3a94ea6a29e910a2b4b2b0da1ed921bd346ed7583ba0f703b7c4ff4edd3acde7d01949a109912c9a15;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4a691cd3f58696220b8705cf5e542c4b343cfd3eed861be8a543bbd6e18b9854e0539e3d2b3ca5e77146f0682ae3d5b913f0765769ec852fc609cc676d113290fd9f379f578efbe7c6be6ed3f0b899128c65398079bd66ddfd01eae6856859a58f3ecdb36888bed851;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3393e58ad20f03f8fa79e22c582aa0ebee0dc086097d7660633d601a37d918cb4d595282982c4da1603ec074b8373a5ee9fcd91f0f98d764f9ed9dac448bd09f5a7eb9c2a10f8d8dab35668b2bfe248c7d3c76d615fca6956f304d691be24358c4f11a23b2e5d4457;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6cedd3407ddbfca9e59f6908965690d14f755fce0562a063c3353268898a822c6ecf77b9e956f0e1a2dc8681f9fc57486cf73983966fdb4ee88974458f74b4281e13d4b4533b9870a9cda2312691a7d05bfb6ee3c87d91dca90a87012181b2c47abab430015e401689;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16b1784be79abc4f627101d7e7d8975668c1d89d7b90d5c113bc12d0a3bd2309576a65dc6c814de586f4360b3e2869477c00c15827b263f11cfd0656a1a927123c4cc4091db9c43f66af1b6deec95e2fc4306b39a8a452726f3b5cbcc448c1ef68014deca0e87e0df76;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177ebe58bd5e833f510d3073cde117c3d13b463371c6fc93a9d8db24c5eb7852ddfdc19956f41fbe575806c7a4c8d4f61bc953fae7739324156ab8594ee00a898f1d7142003fad6d816876e0744e3ba2c2e17a9104695b90a3891553d508b1c3f90a06dcb4fd95d54f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d9be37b7ca6fbc835ffd276c16d5548ed1cf070c8d9711a0c5777dcbbaedb2efd9f060b3ef7a6e27420b4bdc94f0c37e7389a7394fbfbcb8940626c2326837d5dcff5aa143d0ba1f68326eea62c0bf57931657c9761d04aa453176031d7a6fff2dfab0ff41fce7e22;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha6098559ef93e0b23ab61cf669a305e4d41b28471d29cec50d1e2cfda6a015152aef60e6cb5143ea44bcc9dc9800351f1010a2e79064c2e0f6d331172629ed0eaeee16da8e4840947a433fced2cd4e68e53179fe4d53b9a265c30c2a0b087c046a72f00f053fd796de;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1310244395b238be2e6b13f701e8dc31c94473b9b532cd242a9ec9dd4400ddb575a90911c03539306c0b6a31a6a92560430537b8b68b0c9137d37c2938b14339ac7d13c1c3a622600876b692b41c2dcbec7caaed0bda358e0861a87e805a66a1970b72e50a0b9f0c09b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144d3c70037bf899bc1ada3372388f01f95231a7f525e988a9a1a8aa2b031df477196d8f351ecb2af4f0c7175044e101b423e17ac4aff3dcdc9bdc86122aa6411e36bff0ad5d59904d685b86bae358aa9c415bc4b66ce0a949fc1e61702768492698e19efa2a1e3ed1e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13273ea9c8602943cf5f54042f1d919518c06879b9eae72b797392d6cb5650910831f742e5032d4ea43ad8990f24ad4be403a9294c65da909cee37cb40661f379d0382c0dbd3b41215b5de85e8aa02ff4f631ad3cd4760b301dc67d0f37658da60a929f39015feb46e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18c814067fb10f2864a5c2a8d347ae68a6b45d4f28f02f660164c0be81b60bd1e162bb21fec8b592eccf48df4d906bf1cefe5f135d926245505f8a2ab4554e72666c547bb541e72ad55c349843d7e9b0c79551b67bc7c3cde569c4333a2c539b1caee8377dd8c8a59c7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9c71fd348b069d15bc0d65b33fea8b998bec77d01a6247c0b511f3b6871881145ac6a51345677c7b39239b3a97b970de932e3aab7477b52d465be2ebe452de18096b801bb546482c338d5e665e929ee7ad0ee8d38882e0bf57ba7151954bbe78d7ff0d640a45530b29;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10d9aff3d641efc1ec98325ddab74e5fa406b56794f4b23403dc135b4b3ade56af42f4334c95facb634444092074d367c12fc92e1d7395d20d479400b39051c9e9a758cc3bc9efe4e82a027863399d40727f423f64ca572bbc1adac5b536e9254e07d81996f16ba7bd5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a1ea9aabd20d3909eaf67f6c622ddcc4704f02dc69faf801378070529d36918b0230ccd074cc603e595b7de03120ef247541df37228de0a1e005b9279b5452d07c4e2dd40c24c2ac8481ea7e5d4d92629b517bda0b708886012766160f50cba427f7148b943c1f037;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18efa479e7497b07103fba68208c555f0a1d282c1a1d32217a95bfa67c30d08d0d7ef15bb6451dcb9f655444b7ed4afe50576e0e7b2d2af95feb20379fd63327a60846b81d2db90ab97dae2ac5732441480fd2b8224ee1b43fb8a32a9789d435afa3a3f6ca1e8a9d5aa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141448f4369b19180a8564363754c109b89248d3ae769e1cac7f9c1b05126baa8626c50f051d3ad1fff256df8d5cfb9d4dfebff79efc5aaf5e254c3f32b8efab8d65757ada25c50212436bbd7f5d2f213cb54d756b2ddffa76314af245893fe66ef2f3591d35401bcf8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd0d0a49b837d98e831cc9d2abff4fc7b145157569497cfee6f3d89dc4ef7ebbf3d35cd9074cf46daf7c96c887c78adfddbdec018974831b173861ec62dc68d73cbcb38f1414c98dc5e33fab661f75a370b74a026f55f36e9bee0a698b6ee6676fcc4f8ba5397d63b5c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc372e8d18cf89ad1eadc9ea9ce71e6884733eb3cc3a2c7173420cac13a490d83a814352030392641ae05e958de95c581f88fa3f48df692479ce848fca5670346b110a2916f0af4eb37f1d36b93828c9b80011971802d6842024469f7fc1782e0501786d803706ba60;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155a14a303e9f28fa5f8020efc3635ff9b157904d39fc3ed551bc7a697bc2b1be32c26b8e8f8763ba68c4033881881c367cecc4930721344aa911ccc331b9d2b3fc2b618a9c1d51ee528b8f9949b29439be3e8869df9647c24cc49299903e999e0f52eb0cd062a74028;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf51a5d2d1e8c528334724e74f8c9f29a735a63fcb8e13709666af9291bacc0233e2ca8d5fe3c811282c022516a1e8866a09d09ae8aa9690963a90fc1a627e20746f8766f8fb3991271ca43a6b467fd80107915b4d4b8f3452aed24a04be788207286bba6f084260314;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haf274be1f8d2ddf15eddd271194548169851d95740a5d5ed73d234c17981efd72d4ad46533dd859b8a224570048016c4b0cfa90c56e9a2f1335231b89ed0439533c2f2cf127759160f272e67d3b56d0323c9d8033830c77ad68802d4c71b12d37798a5eb10edd70b7e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4b453ef827dd80517240bb80db3a4f4adbe22891e0b10923d118025699c23ddcce188cfeee2b46d5eb9c9a6980b641432d2d35590ad81fb9bb9a7b2399c3b68bddf398a472a11bb6e7d638732b6daf01566bf12d92f17cd115e17833871ce6bddaa5ce862ea3721882;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha500ec3f59d71931b785b14d11cc3a389cee89fe2499b5eab475122aa666604174bd2643a8e7a902d9224fae9640c23eb4a43d117938d31d57181970fc8f3b20ac0adad68a6d49db7d72ae01c5b2f7960006237262d5215950ceb5b4fda36c8d9c62097412411017fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5eb73b7513d319ced232c6bf675eaaf7185a7fa21dbb7898312fd39aabcfa6f0c0976d05f72489372fccc27e9b1b18296cf53cc26ee777d3aac5c88cda79e501090e81dfc8a0f958b41977abb9e90112634dc1a55a1f795224facee8a2ece7211c1fd74576b4ae13b5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40435d12a87637566a9113315eb0eae330271727373d1186e885ae3ea3074c1cf5afeee0ddec1ce284c374719092475ec28b24b123011cb6fce9cf74617fb177f19fb109127f1187e60ba63ba402149fb4e0fd3bcd59d1f8e0d39385aee2b4083c7ea0b61d83d5e1a6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e1a1aee3211cbcb55d655f350d38cfaba6f61cd644aebcbb94d18ba49b0b2a6b4880ee8a2cec89673ac7b8cdfe1609a7f789be441efa8592e7005a3befff7db1f2336d09e92762f0478e84d04bf7217bcefa03ede475a6aced62a3c918ca369a155ea08bcfa245033a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14339c4c3b44a5b2ec6ec320e7de125173911c2af1998126161fc039ee5be6dedca592eb67ba4f14d9892110b4428ffc1714a30b8920c95d82a15fa317293acbc46ab334abeaffd9200397f3c38368867df57a2aac795a653f17922f3ee501b585a734fa7b95c0caee9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b0823845a3f3a45f6bca81a2352a9f66e31ab148f0ce4a1afaa3c82098e54c97a0283234de613d253b623a844699890c8de62bcec11bfbd2038057082bdf752c5f296b2c084f59e72ccf15dd9f2e2fe98721064ca505f5b12efca92a40c734d0d8a0f90690d4032d2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ba3a728dd6c8b9c973ba9572b941e2dd283e4ea936d5f5f3140ad93974c7667031acbbc606a47bdcf129dec6c2c091dbf90dea98b2d0fdc3ec6ccc06563786de7476a6c7a4bbe8b2acc69cc54f04681eb899436656d84fe27bf71eaf818e6c3dcca634fd50a180e81;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146342a40665da8337b933619f8ae15a81a162e2f7a218b490d5f1b8c604797dee322173b21f86486e363da67715635bdc6c3bd92d761c365947b2575679bb4e93ba3c0e04f47380e8cce78e148efef4079c418f89b1ceb622c82b143aa6416b2d479f4f1efd5301538;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a5b483eacb0c03fc55a25fb60ca14b2ef36725d9ab127c4bdeb8537651cf6ecc8e09003ccce7bc096eb122e491ad1ad27f3625baef812237f89a5ac7c878d3625113e2ae9c532931d72cdeac672bdfb4da3d02afa59cfeb3ea50009f4736f44d37df044dcf1f2cafb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e56eddd95659c83a5bb4bc6ae77286abd01a449a2e06d7f5607829e2abae4388172cda2b97e9307ab665822725b161b9f21b120716ceb9855a0a199fd31d72e12ec028af4bd9566aa699571bfcd56e22fe26d070fedd2bac866ca689907526c9e8baedbadc92abb6e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10d221d55a193afd744acc11d91d29f5f1d63ff95f399e3e0aa022fac7988d2f10d3438502a4f728d4e061836b6a29cfb6fd235acc2c723d8b20964bfc92d8ce925327826a95e4835f99127447f9a62c43e47c9f72bad260114770fda33f105ed8958b9968aae7b3337;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11d2879a5a2af9132f4ad756fc90a35fc042b4547dcf1fc041d805e3fe35c3144100db320ade2b99e6eb9595d40b27f2e6b060e2960694424d52f2dcbf5e9865bab467af6296806edf89ec26b874a11b8ecf737a11a8a87471cc32b5c0311ba46b8bea0065bc2af5308;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he3c0fc521afc1e0f96a12fe81b63e22a00717d1d8c7e4d1f300cebe0e50d50d64336a03848ccdad28b650313426331a3afec1bf007bba44cc3ead742867c77b21b2b3ef2f159a7e28373481764caeb915f755ea73f15e0285a889156358aab93f646c4e66084623f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d0080e22ee24890f1d93806f91f0fe954f376bac2480baceb7278450c9ac472c3d7c2b0aaab49dcc223109a5fd41b1c1a900900a9812a586384bb5563da64cad719821e91acb5cc6d84b583bdfe00cdcd91a50bbcdc34452dd23390120d23bb4142db9b50844fd9bec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c6bb9edc88b37f025bd57860a31559e269a910009b16eba39bcb7d880b109624c553eed84d1b5b84be2e47e0539afb51fc109e4269bbc1b4e0d1320c75bbb568b3b688fc1e5655de06b70d10a6f7c217930626452238096cb2b03bbcbe3d80c93f8e03664b3847ba28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf85e0c670a83e428434b22d23aebe94641ce5c6ffda73ac8f0b74598b6771aab5359d293d9a817df804d6749131e9367c7b7cc29a2b8e7d9b3c7567aef6afa78de4b407a0b4cb21a5961b0ed82763d75e27c66f69d3b6768cba96f7528066f65c1e3e2068a349ba9dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7c0399ae3f59263d2837522f160591587ff1443c95afc2fa0c2548a1b893c78f10e8d741e9eb054eb5bcf4da22df4e6459c1d282416fb1ad5bc59ab573906132588958d223ef4004cefbe815efbf68e8f146d1181eea1d375c4e1014a40c527df42ed7c7b868d0d3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13481fd711add40eddce4e8202860d11430d8cd00491c077977b857a9fc8be23d8b181f4be0f06fe3f104eaf15670b9c934118e941748aba9917a161d7c5f90082dd018a4f138f786813141e34fb30fb4ccea248585ea6c0983bb7e8b61adeb5f8b76cd559124fb384b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f5c6da65e680d2c112d80cd5963325749e506d139946017c78f35882c9293f3c1362b400288bb0ade1f6fe7a07602fd0e3c59838f5aeaaf1683eaefe075c6ce2d6d73e6899ee4dc68abeb2a0c6a7fbb20b0a5be7693e6844c4c623adfd586c22d11036b835ec8694c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72fe8b7c16f038e5bc25b2acfb38223a82c8a1c31a6ca8686a77a9a261d7dfe8694b1e9bd53c2af8163c83e9ac1ada24d7045d9ccfbae6e033fbe507fc8d5db691d3206c22ec7aef87cb9a3543e0ee281e94776774edc7dd4691e310f30e927677c4f85a4c648a0f0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h70f7ae324f7a877322ec454c82fe45d48b0fb0e420f1f88cc8d55f12c8c1a2d5d717cde45b2511cf23232e8e250032e677169d951e4d9b594eedd0876fa2bc699b4c7a8144a1a9c4bd3c591b60934c4d4aa442d18913bdb3cc07263eb578c79f19763acb9a9c79946b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he121ab28b13b9cb2aac3c834aa4a0789340f26a4567dfaa808043ae97da382798ad362ae0c0b1b4b28c80e10625768bd4a156652454c7de1f49b0cf646f238a13de6a41fe7ff18c85d1ae05807769310aba127b776071ff87dff8d3b3e017eceed71dba344761f607a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13d587dafa0caf96c45e0bbcc670232245d5856ccaf4c01889d0bb227e8099a3d88429698cf1167b4e95935b3b07b8c95e9c72baf00f8e57af798898ce30ff523e0d025dd8949e5a5e213fef98cb827fb38986cdba135ac5a37e4cd1dc1914a50156e26b2427b750b24;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c5106871559161ed3b9c44bac5471d638ed984c69c4d4bfaac8c9ec786a18afc42661d6245ecd61097c1462ac77bf2693877f0ac4f296410d5f7700bcfd6bc7bbfc8432af68c2c8b4dc6cdace7ce6317fa1ccee0a6215b212847c60f665770b1449a575a120315afc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac3532e497df27aaa1d8d99a1467aa8f00492c1cd523de21c32ab5ca10ccabe39d1826e00d4b69cff5a92fff5a3fc956c7360cc4947c67aa84522cbb3a55405c4fa42e5e34ca8c5a89d3be271814e11012d52c3520e84da4c83e7034e48e245b266fe49dab94a2a727;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a27779d53ea5244a253adcf14c6f68b16336055dcc63b0b523cb68d688b9068a54802d1c07606e92305ac12814207939d373eb09127b1d22ddfb02edcac30ea7ba1dab93e79b48ce9e5ac5ed8731fd0082efdcc4829b6d185aa5a7d5648113b9df6543cbd2c21b9c6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e3017120ef3f143632dcf2c77aaec9d60527f7af53ccaac475332e324eacccdf636f510034161598c43db729c171a2aefb109e49a4cdb298887d424dd2b519af8e093b066a1d09016a2cd4cd191336007236ca9db9e41cef3749600b475c0dacf9bf1c854ebfd12de1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5a4889455b9b36b20df2f52644e62a135de24687f566735b60db883c5b5ebf62b9863fb47bab7d9c6dd69719554eca40a6ccc213229eae8da59b8e59f44a3d6b08e8b40852a9ed36608c0466dbb39bd6dc612b83a4583599bd6e8d7586bc3cef80056a9062db15de9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a8f07230cb8ddef98c40729e3e47830ea4d07eb83be13476438b6519e8c4e746f4cbd4a531bedbf327c32a989e426c7795a452d1f3192f0c7d553c11baeff730270272ed013c39fc27a4584e9c75517bec077ba654682aebb67e9d44a002064e32e2f2f056ea755cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h884cb060d5967274089d18ec7619b29eb64f8489cb1167dda9c398ded73848a39ea1b03f816ef7a5bdc6f6c87d71218c837c19a418acb1d931247184532d61505ccc7171ac8447d251ab823194aa06f2eab18e7357fb4777e99a89a75ec611b5782986f43c07bf60f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h705b6cff269892dee9a5a6b12c90fa32cd34e5fe338a6ee39ca941d5998aa2ca98ffb07e57d230e4506b4acba326292bc92341019113db6d353a2fac38f945f29720938d7882d0e673de608a144b23729ec84dac0a22524320055298881352c49360adb1c3adc2d265;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee7498e7bc35fdc7fecf07cad15b0933b23925c27c0983a074076a2d8895b6a17dac659bd9bde2117ea17eab556b6447925da2f12e5461357c4f90444a7a0abfb7df971d7fe39b50a9a66fd494f5d63e92d818f122f6bd0aacbbc046532cc435fdde5e2a9b317ae2eb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h106c20ce1bca03d0b26c8910ecad056fdd1a682cd06fa1072c979daeea2fa92957f34abd3f48ee36d5257fe46914eed0f6c840571dca1795102177b0b7f839978f89a71bbd41e79763ff242e570d42040ec6425fa8450d8c9cfa4c225ddad5808b0c47413f9f9ea72c9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7cd1c0e9642318b02ae3ec605b7572f4377282fec4f32bf741594ff8d3ec008bec254a448c25ad4046bd2b05565b08311d96baba6e8703297de846d89a5481678aaaf95c09163db510d23b976cb17c40ba658c031a4f87ce0298698ea3fabfc5d2a08e1eccb18f3b2c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h168b7567e7b510afa8f91efc06914fe5b02f8922dd9a0601a9ddefe69dc06e4c7bab50e0911e9bbc05baff6d9025070a11c8a86cf5f9b4b0fdff4a45e92fcef70d7701e1f730d6dc71da8a5865122347ab0d6ed5ec16c58e9f7bd10b04bab1177fda0e5ddec72ab8be7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h149f94b033cb4fc225612a9f9fd52bfebdbd01dab43d6add68012ee4b80594f5f8717bcea07ec767548991592142141026bf28bec8c394212f6a9d247a1141e5d2f5b3eb206435212d192f728993d79e92aba9e1a74dd03e5533fde30aa95418b29114cec28abc6105c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1555b84a92d1604e0cf530dc741d83125b31f51aca67ba9560cce8882954434e1421613742d005914764aa8a8adb9122151ea60e4221e09e5ddbab1f2fc245c98c8fb36cbdc104c3daf5dc8b9a9b995bb6e8e3ce7290ad9987ec11d0fab9387521883d3516e3de8f5d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha6dea59999b29301a21463f34a765651bb6b87bd5acb1da5ae01d1264281486e6ffd8fe95a04e2f742d026cdf4302356317f73cfca2d5bcd82b2d307401963f1b92eb9d29edb45faf311c5a21d8edb0304fdb45ea5a5a03218390f34bc351dc9660b9fb0dcb5dc71c8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbc2af61a6c076f1545d4ceb6b80e47369287f0505f72c891a81ed13b4bafd6e4c4434ca69496b6a0b608502d433efd569063d0162da5e5846718709b0e0e7876574862b015ebdba0f4b5501e868c2bdf959f0f9e47139acaa86af269e197dea8b5ad037193637da496;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h377751ad6e1becf2bfd0c1fac8f3477aa14a2ba5ce81bc5d177f9c3357f308568f6eb73414c839bb03a575e059fb7786fa1f130bfac5f8edcc93d9c66afba84888a586a8fb91ce5a4539ba8b2e89eef52ab0b58f863392e8d221c694464adb1d84c4a6df2bc0701169;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h194415b05e415c4d68f28eb5b19ea4218c6d87f899d2c4652aa4391cfe1ace01f26f1a90fd4312f85f1e51b655241be6cdf181d58b1fd62c7b3592d999e01991944e66888b8895b7c0309b9f1f12e8a3df4b763f39c6f7e1461c446e9ae97b5e1f5b8e8b0fed6c7b30;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5334dadfd6b5c4f9eec2eafa4073993ed4affadcb25759cccc104b24542e9e0ea0181473caef67ead354bfe2bb57a4ef179d5ffecf4dddd89f0c76d94d63605ec50e9bc98b9d04a2b84d3dbe9cc994d6de465db9a336f7b708ec2778710dd5e7a1cd4da72d43f610e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c90ab9542130ac953472b772a5f96126718308eedb42133677804c3091fc3c62f98ba66a829186370ab228a9170457d0f9e2eded093cb32dd1277ad6b25785e65d3ca17024c761b72be9fe1511fde94819d1e2cc52087dbfc3f2a87c12d65e1152bc2c26a077d1c8f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17a18dd2482b8491cb2f5462e2c0ea194c22f2528c2a81ecc6d17a44858b464a7c4e3d0c10cd557f3b500a5468c604d2404272101e633cc71e946b002b13d7f751f565aa243306713912b07abfdb99131f52fd4a90df90fa6da0a79bba76630263c28583eb83eda907a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144a71fec82e115f68b0f6db3253107ef9e1d12de8243fe3c340b6210f3e73034ab90efe7929f6ef0d861bfddf01bd17ee20c08d1a91ad8ea1e7b9ca83c8028f5bc48a950a28abc5ce668e88f37daf1e04a925ea5fabf6447d70b509f352b3ba26b6cc7ef174360827c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcbec3989b85f192f631b258e45511f35ae5e8c25cb496f0ec6ad05c938670e2ec8201c330b388caa8fc1a07823e77331bc46b9ef2f856bb881e3a90f399e3a6964cf6c2fc7623f07695741a6b9e43d630510e32423fdf4a1994283811a0695030f62ba82215fa5ee4c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fa3ff0e93eb10d2df054f1b0373eee2e586b247fca283ddcec54c553f3af7bcfdc69c3761963b9ce3316c6a9e3961c739942ba570c8dac3ea361dc09e3e9e7c2043736300d0dc1f0c7796ee41bd40a161157d618b98b9006528c5414471a17e3f7db308bf7f0e9009e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1e1eacb07af7f8e87e06a9f59563def48d00e7fa1e23e7ea4a46858a76ecb499ca9d0c7a32c37f6f415d88cef689d755cc865f9160bc5078afc77ef9d703f557ead6e56a300a166db595741557ba3a08e9859a5cd5cd2bfdfdb80f3a844b112c530f2c7c62210eca8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1403e254960f8445b2990cee291dadccea8c82f80d4b39ba14cdaaba842a194a4c3e6769c23d117c4156147ecbeeb09920e77df84977a681e99ce23ea31615454067aff73e3cc74877c3e4c35b13750c7c8cce4b7aac767c763d0a3ec5cc8731a13eceef8f451080476;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1420753a736990b4198be5fba4fa9deaa18511e62d1b6fa78b8da21d0de483c922f2018886994d72f80979b36a37f8683b15f1777bc88bfa74e49fdaed3b14a840d67942c0394147854487944e81a789cb4f84880956fc1c0d00b0ccac1d29f9c29486e87b680dba6be;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113dd65f688f38f3b29abff45f92c1a75cf9948641332068234f1bf227fa4835cc683a7bc52f283a92822f2084e8afa872de611dd99917b65c5b149bc9512f6f0dfd290001db5a918e6d76ef0a21e1a3b4e65489b08113b430b2987b0ef29037e952e1ab1fdd38a05f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h82dced6f104c123ed7c810a56e6e83bdc1cc1ff12258b12f8a79a3e30abb497154628b9e334c093ed43e4975f28171809e0af63381b0bcb2a5ee69f63a65b5dc7e1ee2911b43a56c6e96a5e3050b90bb79b2f15fec7cf3937f2f3eff6d4a72e00734ff28476acbace2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h137b2f351d9abe9ccc100ec5f97cbd3e2fe391ae3316491bb11cfbffa2764ce92009eb2cdd7ceda15c078f0e657a3e154cc39cbd7552d911d0ec1ec185eeee7bc29a0332071e2019da7b0839f0b05019a65ae0fda1a62a84dce72eb05bbf7ffff3814db33a296dea96a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h238db54ce7ddf93aa5020bd525c0fa45a0c256f98ac489972fb3b762e66243be4e539081148c06094255c43383c2a2a99b904dc7f76f5e41e026fc62bf85ffa64f826fc84e05bfa5c41e5ce6da7460e3d051f9bbfd20eb8b570bca7df855fc1f9f3dee6bb04f8f5508;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1df5663e3552594c9d7475057bacaa0414b43782faf04ab3d170a2996ab3c2395a27f83eba59f89608f71afca4dd007d6331f3d879f562ab5300fcf16f33a80914a661b01530d1994726b6935e7ff3b57e0ec13e443d8cd750762cb241e7b4f53e5dfae6cb9a13b725d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e829a659b30a8993991fea7960874c91835d4e9b38621c85841d5102f38f2c3d19f923976b646e74a79aff3bdc0cf4f8c65f0a44aee39cce4f328de975417ffb73c9b74fd380d08846f21f0cec4288761d5369bd941a97cda0a16c5bedbe15df4f07f858dac3c8eeb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae53301cb9345ea16c63882a6c7a6b8f461a73a034735b6b4bf9782118941c30cf0b51b310a09f8d4e3f467a8e025eb8002b5150046a5377670942c50ad9a6e21650caf547b76248064ee41a86ba32c5e61e5da4312793d6fbf4d635736e49188dc3c8235f9ab04dd1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155f30fe39ec2439e27294216167186c1c7ce37756a6880549726fde3b80c9795db6cbfa16e1fb52865ceade8c0c84ea318e986d095521777970819deca69d8a904e046bc57505bb928c3ca72eacd94b76c688c0b808f4b0acbff20be85d269a65702852d740514363f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h176f7a6cd72fdfd6b9e71347dedbc720b022b3a16c62f3482ea066db92e30be8eab036d568e7d45f7da25911df9ba955c734cb867f7c068cbf3ef30b473f0740e6da815d122c94e0dd5b4c7aac922ced17163a5f6fb3a043dc842e6300a3eab2187cad52694ef121b60;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e3f27cd88f7ecead9dda38adc553b300b70e6c9bd7fe8e104a1ebf590771f7bfa74f909007e93a3108665b6807d5ee43a5cd04807974280af8eb5f99fa67c84b26df65a1efb4b99327788d10eb20d7f0cfc3c74ac485f6b8fcd1a922cbc92514894a7d0c5dc2a4c9e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h179430740b69b353be5a06f0fa9d481d391c9823e6b01c13f6d85eded72d5a8e47926b6232a7140ed98a3e7f5d5dd2f7503ac9c0bdb566d5afe081a36f59afc28cdf0b0cf6f27e1f52b59ffc985fd7cb0a4ce514dabbf2f0e0353dbe57d50ca98179d8841fab7be0a63;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9082027c5eb022a8d422dcb28cac6817db05894b0776b013a91bb22340a43bb5fdeaca8c55163660647a6f232537a834ac3252afd872ee7dd175ba2f3fb3f24d8aa3c7e0f5e339eb869caf2121660b26d45788183759d3f3fd14095d17b61acc3a524bca60d4313180;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h471bf1f5bab7cffba51881a77ce45d50186e69389116538b32ac8c71a2b7d3c8e3a0dff5a33dca49b266d6521a1fba2f699159529cc7b3e5e18650a947f482f3d743f640516937ef508a5f32bef1032098bca5ef9c0454884bb3e4c9cdd07bfce96dea7af9a716e7e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7539fd2198e198ab654beaba6ac92a50cc96b570748570ed0a73b11d6c890ee841d05f9db56576879f4adb629a2858e4e24313a016f448a46139388f0e36adeaa5694130bbcaf8e0e80b8fc3f27b66dd3034936ab7ba9af2d46a98c74ea403e191806d436df3396353;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b9deaecce332fc13e6527b46785d709075bc1b18298e88ee3c9b64a25dc3d077b060006e27bf30de1516eca67472ee1a1acffc4d3283c8a7f88cecf5f1f93293609c7e8bd0e24e30d680ec3509225232780d3322ac4a0ec59c40a8c79bf281a5fce7b3989ecce3ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1964de5eadfae7bd47129a0e2bc5ef83a5d42acf4bbccf5d478466b83235df71d29112576fb7ec98ae149e1eef2e598c166ae9cef332f7b67c1a568a13e9266edd6a4ff128378ccff5817fcafd51e6bde93ea42e594cd62e0a50c6cf2dd70b6d5012ef01eb72e1062ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h132104f556ee3f22639df5c65a99d31e6ec6d40665aa2e0c0f1c2280b510e843f30614a32998ab9bc70fa4e9f8cdad7a8fbec6beca6a2a11d30869090f076ae6d740ce3de6670b407c8de58b2c3cc2735e416265795bd9a795c7787dbfe2e4177ccc611a2d120fdb9c5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf1d6788e864ddf58712cd1d44282ba816eb8df74247df8b3c27688a1424568da8137868085624a6b3dc5cde837286c7c9a9609056eb90de808bf9058bf01c5d058892c1a89139924e81f470166272546bab3f95f12680931ed9f6abc3ca2dbe76b54e538903d199b72;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1edd5f773ba85bbd716a1b5c7233f81b122de9eb948a6a4bcd98e7c97711f3f8ed03b458397109cc99fe949fa0b055b355e030afc67266fc15d103f48ee73e091f05f44d82b8587edfc48fe6c0aca5e473a41339993425c6dff69873515f1c97c433cceaaaebfaf7b90;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1759694c9354750abf0a688a4f607fa073d610a77735026a5b94bacef9fe0e22485df26655b39a5b654af5759841e0ccf21721cc79e50ea0d5baa1b0e4ea1dfaba80878f40741a218873d20ae81296ccb3b33c572c0ce7ba2e869b1a29ebd2968304220008e30a57b5a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d1d563c93f43379ead4559efefed8aa8becdaebb06ee12afeec1aeb503ff3a9ce66a28f2326e611bd63c9a9b02ddcec41ff960dca4e0d6a72fb60dee47610793fcd2f92dd68ee428820c970f46971832dc062c2a9974f65a0d40c94589920da2b13b0d32668c07cd75;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be2b121b0f8ee83573415bba1e4797950cf21bc833a33c6184f5b6ac6c0fefc7bee097bb7a5b3bb6d4a7da6c3855fec9ec2e5b7ca8025f58b3ac2386a620cb0511bcfdc2547686fb18fd2bd567be1f64680fe86b53e09934207e72b19833db7899415eb85646ee15f2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e3e75b4455bbf6d113ada07d9c64081bff8b97ea329c245d72b8fb017b89420d046b2f2ad340b8805e9fbaa8ece2af169e438d8edd29de96554e21f68ebd9769a51c7665937f55c5b428e1da6690a55a9f950d9f66ec3f0d423613ae38ca1c87df3da50d244aaad61a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ebfb6aa28c966dedbed10fdd1c2589be233c4101c39efe288ec68d6758abea54a91b54b57337e23ad3ad69df3390571177ca45b7b506e01723064abf1836f1747f3ec5b5e2d6c7a0ec52a9ad853a3aa8ff6704fce0e95b1427f8d1795960cb1c955efbd74c92cd20d4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25fe9b669b0da17458ce339aed1e4e91a78c20d662c9f1485c2ef1b386b96ed7167a8739596141b0337d5598b6b09d9c2cbfbd0b294c5714e6f7bc38f0c850228cd788c70592da98ed324597f09fc30763bcc7f4d9d9e32d2b9c11b2609f8d9d4949d8642986509a78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e37a4c1600c419f54cde995fb619937d07d5c6591a8f6a651eca5d1b3135ae6371a71c8f14fa3d1c6193c6dbf18d5c799a1441af6d331d53b1ac46e1fc50f78a86ed55ef97a2925194e09e7efb6e307eca1492baa3c0e2bf7be00f60e2582a68214735881eca2deffb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5516528d3be63417225c953ce09a8a85843c57b7592d0070385bfe22140fc73aa728c2f127e2c192c5975d1b4709310278410cfce536cdd8e7904cbc5a63443f173ef9d8d60047cf5ada91ba0193c805a3f105a2e8c708fa620b93ed097b54c9588ebf8359ad7144f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e5cd8a315272efcdd46c69406939c8a57ae40e4feb8962e192192d70eb46062fbe111e99768f5e16767d41783ce068abd24b96326b0d1ab54dd6b4a2a0cb934465f5bda70300a5380b91c63279e2628a3a41ad3f6aefd014bc6d31035bda32cc4c466df441d695a916;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h58c24bb942e490638acea9f06220a598e30c369e79f0f7e623e51cf7e3f9c5a18033a4ddf9bdc44d269b5862333153d5f36adb8d84500f23d8ff60d34cf87b5fd015d40d424308397173ea32fb3cdc3426b640a1022aa2b351ed041b6424277523a8208e19b3a869ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9bbe4907e65cb8006d1813dfc42108e0ead501475353ee20a981fc457cf5d53e253fde443da15d2a9cfed78939a8be32fa4bb6a3092769d441620195207a7dcfdb43a0341cd3e81f1f2cc9a01df4eee2bf8a5efa45791510cb025ce179d0cfc9cc846bffeaac1958c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c765f4f67dd57aa1dba883b27b6102f9a0da71afb1646df7d35a8a55b9028185fa6d8b22734b1f10010e35b1c7ce175cec7c6fce7c4737f81c16c3bc5924e49c6e2f0503035021e5cb01d454ffa01755687986adc4c512c7a1600a29f374456cb55c4cd9ab9467bb06;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d9b7110472fcfb6b98f33957e6d92a85d3d76552329cadebb3c8e3e71095518700a714446884c4b75b642f06036d9f4030ee94461b915da3866b4f52491a8d328002d4c9a2cd6eaa0cd380db7405c41c1700bb18eb6c1f09eee72404bdd27dee9aa6b8d6bee393397;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb14edcc851a29f857d12eafdc33f5583882b0ce82cb48e4b7da8fb9dd700b1ff3be24e355ff19e5eef632301900051a76b4bae5c176d9783bcfacb5db21f04cb99e1d99940e6a5f1dc4a14251f2cbce4ca503de0ecf3dde845894089dba08b2cc2692b89ce2b8b73a1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13c3e1c9373b3e2ae522aab256b3ba0f003666ac6c2bdb385392a1cacbb5ac855f5e3055697ab9ebb4d9241c489f53c61ea909fb1b185d6451907dbd30ea19097cd678135c7123bf328a7967af4c616324dde5bcfc256b2ecb17fc1118be13edae4a0b7af2ac4ddf22f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11564fb06d5cc34653dc205d6f5d46d76645350a4385a813178617072f66a06164e31021c7404a1d243bbdf14d159c0842027aa95fd09896068493f8a2a00ca6253142f300897295bdd6e7a857c5a5435383458d0af7bf892975e101bc60546dcae7c04ff2743f752ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18230b7339c339fdac1b36818134083ffe9f8e9c1f3a0a3c412a560e3da41bf1b429c4e97b907a0d92f9d695268c45fa91fca4621ffe9aedf1ed53dcd345d427580fb19027c30fc70422465cc533a62318eac17937808ebf65615555ed293ff762e36ad79fd5e00a491;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e92a4e701c5acff9721b296efca701be2b74494f8a4f4231a9283c31362d9d60b86adf0efc63400756bf2bdc89ade47ee910b4b0240b383dee3c8bd7d2ffc7f1a6abd1b3c68c3004499b41c857799f623651ca9fa0a7193cd4793dddf1bea3fb6c7f6cb18336e9fea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb6cc172c828c713b15ff284879da075666aa96bdec0e6d4d6615edf3ccb0a3a8b236bdcb70ba55bd3e36c15ee6668dd1c22e51ba5ec36caffe112e91366f43b9d522e476442905246a8c4abb53a6e802a4256e3a1848e5dbb00aa70794f5051d841c4e3d12ef41f66b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h344a5ca2ff4adcd5e5f3191aee18be43a4c6c10cbee61d2a4559da87f06cd961588ebb205a19bd716f481b4aadfbe239c4a4c0a13ea7d69ed3dbc3149aa477119286a3b154f405782f2f252dac4a476ddd1fa91df1a04021025a33463d62b488a41da7d388196b7ec2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc33aadc61b37597865d734d35a52a68420c98143cd83565fdaf6755ae216fcad7962b27fc7c82b7d004f06df0cdc255b2614996e3d00416b267422cd817641f2f089e20d86ee50e24f30d9f34acded45ae09b4c4143c29c097d9021191e9826c765f3d33688e47296b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14bcc51a269bbff9e125ce3c83a491b80578e9e65337370a7b99233246934d70873297e16c903f808eeb6d967fe9d8878af6d57b10a7a5c308eb31ebf66bfd13997bd93c726b3723d802fbc26d8b3b16791a23ac2fdd58b2b60523c5b8315516933ad48d349ef1a299f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heda38d927ba9acd990f8c2ebfa62d74fa3e4c117c9d53778ec6ea0f0388418897f6052e0b3ca643b7e887cf417a16561e91320f554ce016cf764bfdd7f4d7adbcb7ad7087f8dc1deba700bc2a392f5e62c4b1746cfda8e4eb97cc304078a3a3c48ebe9774a9c05aab0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb5a6d212456834d18c2a2b35d8f5b0f3fe6b2c748a1ef15cdd941ae697f3b2e38f6055b20f5e3ab44de9c5ee3e691a5605d106b81d2536cea433473f94b91bc3740735dd6d585133adc26a5b9c6177959bc885e5740fb6a04cae0ea5bcdb608d063733f56f9ebac79;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd9d9bb6a1edf3d12c2ee91552e7db03834a1954f4fd62bed17eb0b8e5a383f4932b75074342605fe00674551a8f78201ff82a05e812341f1b634923aa4067d2f90ebca3b15ab7d60c9f227c4aeb795265c8392d77181489ba041beb430ca69f0a5b8ef110e1c71bb11;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1174bd011f9073bd56415fcb2be85ae9395083dab3056e803ba0a497aa6fa5b8ab01b730e234b4d86984ac15d1b3812ee3c69c31e45b71c27f2935c414247548dc354c6918e7cc891d9df5cda0f65c55e08e12de314c5ae8b7dcfdc5261176c53f1124be3d56ed1c2ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h78263f11e9f586b8e8c726ec485f64ddf24f25e3134241e9cf3bbefcf5a4888c073d3ec83a42b804ce8b3bde2f1ccd57702a4a3852df9898218a802f41350a368a60a40b809fc06959d57282838f66608598ec8f2df0b06f600f3902b6c572215b235a929b4d7569c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e9a18fd7044e0cf47ce314c17305b9c080e3e06c671c0963ba26a950161e09ce456268cacd4658850e5986a1901a2a68c8ac9a9eec9500095b2597d439a62e84cb815b28284cf60e95d92e458644966fc4e280fc9c937f3f86e6759d022d41e2ca65c7bdc79f303581;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h945c23903c8fdec0fadc43c8c09d931cb596aadca9810220f8da944912ef4ab9825e641680b4bb9f96c3d2c6605e0925420630023ddf2db9e4871ad2a21ba43bed542ddeca8af2bca5dd0c021f82a3167d8f2db2cc13140f6dc1f0fb035f44ec9baacbc48a636eaee4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1960b2d259184b8ba5ddef476d75689a27dd83e2e1595b605400ccbbb34928fc72042c47a8f3788788400c8fb1b2223fa6bdfc7c541c84a581d8f307b6f0d850369980dd4739f0634aeb4ed20812cb98b904d00bf5cd251f31ffca95d0bee75ba3de25ae860dce04df4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16abac66afa39eb45cf52dc6b0e57e56d9380dbd34da797528ef2f43c9831540b4512249033fa7c304f251ed3a26c8f2847e2cdabfdb2d96d3e7df71674b51ff42a9ddc7aaec158accac17543de81259660b9c53d46f81d7434d056f63aaa4b8fe13de90e9e4fc11215;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13db3ef8604072e7ddcd8811ddf7d7ea58c2153ed74b2c0f5e81211fdbc70bf311476b99b29b740e65f078cf8b9fa14a1c4073822917dfabe9827385ceeaad3ae2d9a47ea60c69708098cff721f40863c94443867523303a37502cd4268d06c7554284e3ee8f66bdb5a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a35524ce2dfb7ee2a7b5bc077ffcd82744f42e2a3b2cf1acfa384e30024d104e04ed1ffab4894fe6fb5aaa0d9800e188219e24e8880c1f7af48d4be1cdd59d83a6f7dcc66615c4b82e32321395b45e7ef7762466e7ff21cfafb51ea0a2c435821f15565c82eb3177b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff590973644213a59826d898ac982542ed1d0b2c4f8c00cae7c71ba310ccf785072c8ac6a97e1e88548b03f21f8c7ae40c741b322fc0a08350ff7bc968e7bbc1031a5aacc5d55fab078cef7341814d1f9bcf9ae0bb54243ecb411f784727d13fee51d2836de6b7d474;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h160b061311c71edef7626584e570c51ecbc33e8fb3b6162437883fa2f8c5660f7af3017d69144c84b53cbcf1cc1d685b800fcce7ff681fa57366a67dafb3f80d23ce865c20b358b488e1d74c358a1a8ab1e1826168d2e01c65954e4a8abe49094c5fc691fe0b8543c02;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h535f36184c32c832c20cf770c31948f580398debf87ca4e520481099151b89a05fe7994e8928d21eaa32590ede6f7676754c9a3b8ac8e7843b7fdaffc0ecbbb15f1ef99450a70dbd8ad92dd19dc14ac5fa9a5080a454e6988e9938a4082c43bd3f33b17db1b80e8ec5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f4e549f6e44c04b5ae3e15edd284fba5cf46e0922dc0a7207bcaa0f13825c4ce11cf52ff140267dc00efc13f7f33a5939a02b6131dc7004a85a7b602fd835e8ff55d8d6c2ebba672a36b7d8abb259342d5de039f8d7d27008f4323ae178ec1cdc83b797274bb4051a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd48a7888187386cab04919821a3c8f5abc4433775a4d0cbbeb5018379bc88a97a1fb608c49c5880a1c4fb8f1f0936619b8ced3edc974806295e8119d4e57d8ff3a29bdadb94f0c57f4aec7478a1dc405b2508a8a6d0086b1e76b3a846325b355d483ae24d8c168bff0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1156b5a9bbd7b2ae475ef137579f3aa5fb4b3c227f3694975e196c116cf538755ed759211aaa5aaece9d810f6c898d4555d90764a44ac5dd2093dd09f6e98e96541101c4561faa9e29083bf66e17ad5ecced6855656fb08ea04e9408975c0bf82931af63f14d9f775a6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h139d3bfe2a625116a53deb27e12c4cc8c9090c81d01809aea1fee0ef938e8df04019e0a1ff2afc20a458d26f7a7c1c16abd323a54735af0524cf8dd4a51ffdc649c3d74264d07d12a4a9b26977633739dfe4caae09f20b67b555cba2314decfd74859136d392bdfa647;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a33b5dfedf9366269f74d56da41c52906462a6b0439f3760fa8ad0b0b602afc1a9cc4fa0f5d857bccd93db60efe016cc555ac9838a527837842cf624d5488768115822fe817e73ecfbea8c2ba269d00976f03fdfb00d8c4f41cc06efaa5b5e9880b1dbaa5983237ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17ea33444d15cafc91428530185d6fd4d8df7d2fe34c6c81558362e792ed3b8f5d1c4d668eda157dcec6c06a0a82be0bd93f2e7382444f08b987d6f1897ab1cbe71384d769153ec6a9faaf9647bed0f3f98e372c2a380f4ee42c781035ede1d554a38e9c41bca74e666;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3eada7d37935687aff063a14ade8cb3ce6842b0178b83e116a4311ddfa75ddadfe0892b9c3cfc2eac85f2cb4340e59bd53bf9195d28b3d359c35265c355b4b5af4bc845f6f8ea46682516d90da53f3dbc663a877a30169ff0eb91110a650f5877c2a4953ae699afacc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e2f4927574b74bca4a24fb34d41c845be30b6a0a6a74f7fa7f12c5c70dcce744011400982589560eedd3fbbef205c13e8ad89c6f712c10f46b6c578b1cb851c468cda44c44b4d3047923d6b2154510432b014ddafd6bf8397b29784e514b8c71e564002431d19637;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h119f861d85bc5a799675596e61d67692b980bdb32190fa08ad702aa9483ade16df2fa316008fd7c7901393b2b4ce827feebcd298345b98c877e66dca6a03bb9dd8e48d3fa5a08d54a81b9332fdfcd8af5c428dbc50b6d308b37587ec94bcfdaf722131c283f559e111d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dca8050ecba8011666dfe9eeadddc2c07aa036a566cbba3881cd476f3cc5baa0b98e9ccee547a8a9cbb1e8392684390f7723d79060382e0c1ee5905c464df07148f044aedf50e6493c5871be0fe2a41bde4b59ddab14328d4c335fa20fee68b90a418ba938c2e5d43;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1a3b6beded5d9f52b05317d9b297d7982cf6b6b9a9625be62d9b38260a1d551917e061f0416a9e46ef8d45d6dbce77f05d48508acf06f2508df2da2276890a20c4710a03166a75770aba4c75436ea7cba66350cf7a0b4c578ec204c1f93bc5489fa01eb78c03d5be4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h182e46660cc683c3f3ace7820b4c65b339d1e04a35e3b4c583e9d3464e05ec220dd847f31750592a7646ea929cf36b34808513a2c1220deffbd94a7b7569187d748e6569524a10f6bb0022549244bbef7c7b9d54c5be53aef71cd5751638b946378548fbd775a413cad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155ec11357dec468fc3f9f84d8d1131976bd39c127d2acb73a3fb80adf0b166719fee4a5209f54cb1a77ae394e3117640176b21507de3bb27dfd1e7a9f737c6a5585924d7b16c90fe101d1e31be6a44d24c78d4a164d97d6a74218ef6f28b5c1707adb1a7031ef4de0c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b373edcad9c891a5b96030380ec60f5cd51c99c1a715364ef99012db8dcb02e44d3d2724d24d8af23cc3174d8c8f06376b371cb81bfc93189250d60da0f66a8e39f6a1ca6a66978ddcc67af13a8d022ff76b52099cb479a644ddd607399995a9ed82640c10b0d3246;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cfdb6a95440f34e4ae4848d407411a25c1bf02fd555fe6bf57c21b499ad6460ddb794d68883c4a3a6e5597f372526e01658b59cb214efe9e62a7e8bc4134c7d392ed491a2f4576de986832fe66906a2e1ba1fecc30260de4554752741c996da3dfa26d7ba668b9fb28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h57e89ecd62f3d86f9b0e4a55556a74a34abc22ba256a8ee948ed74ac77f9eb6c50cfb30472790f756bf640acdc9cfc70d4b1fcd881eaba484ca6ebba0e020ff1aeddd7e067370340de957bdbc348d64c777224e46eca114aa98bbdca6bc7d3492233662d9f222746fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aca8229307996b0963f13ab1f12e3fceaac4a67ec531f9f125e7e223e3ebba0b32427cb7d3eea56c3b98b0511fc3b006e0d96c174039a83b5b0030b48399f1190eca61bd636fc0216bb78f1b3524f516711979555254fbdf75c2bfafbcd5000d99af0ae840f9ad2974;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cb28d36a0f61c44d1c7c3bba7999521ec6a53cc767df222a3e27fc674a15cb10005b3ff2d0b1261fc0683de098962cf94a879f9c0bb9ddab85f57c046b5a2b6ca5b0d54f3e6f93b8b6f46fa03306d8870c97b540abda21970c4cbde950f819a8ba29538f4fc0d8997f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha5e1973e1a58a329f99f088d889b20f65f8e55c8624c5cb14994fce44f1a1b6373bfd572db8ee4e977740db74f3078eefd25215562a5ce99388515fc19972db939a82bc2fccdc933038cf73cb171729f72d69e8cd587d514260f6908481895a9b3949e8c831bbdbd4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h840406c28c9c50acf22357aa6217e01655862061e7a3d5888491edd8968c98e85abbee2b28cf022a0ebf1689f4ef2c60b7276c1db6da08319c7eb8ab0d91e6fe8833f547c770f234aacbbb2cb6ff1aaca0fe30feac5a84df0ba644c13147ee4c914bb0a3b399e59471;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b5982c80c4db02e62a9396ed7976f39a61ad0d32adf30b41f9f81d568155bbdd2ea6fe9a363d1e97cad5abf4f66f2fb319287d01f273009d7c15e7aa977152d1fb45b5c42910d2727c507ddf5a46694f848ce98d55788ef739e7054b366963af51a7d04938c5977b56;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16ad8956cdb76ac20dae2e1e9caa2109c220d8f974b18c5f902d3ffe3e457d4bdb1bca704534b3e356f190eb14216bed4d4494c9de6a96f099966bb987f8dc654a48d6c77f8015e455b27768ca364865a125c8dc9d44247db3b25891cfa1450aa1738516a6dcde16823;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd74d9d19072fbecfc35447ef7692bcf06c759717531234988f73d67dcf8082d81fe9bcf5b28097cfca00a9ba1c3a226ac8c19fbd268d3dc9efba3a5ffe93546711e139cf18786f8ce0bb10929bd0a52ced5d90783a193221ed2e6c211ad64bafa32c0b2587ea37f0e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd2678ea12a6e196c55a8db91e3db118f2fa20eeddc29cf69b27ecf1edb54539cf66da876537b23e925a7e0beeecd9d6b0af38cbc4d1e55c7bed03245de4c4352cbe244a167230e4be5754068b63de3b728ea08aa12832f5dc72646da72f974aa4465e36d96f1f774bd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12fb7fd136e1c398190e850ef49312cacafb18b8deb8cd6034aa1ed467118fcab9c9a10a958561c6d0c0ef48fe8a8abeb0aa3b0233579683ebc78613f033287e5b2035990648a4b6391f02393d463520fbc2e6c4053fb240afea3bb24d47baf1a7f40feced13f2f5657;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc74e1ee4edbc7c09b44c5b8cc4571a8dcb69c68fe14eb6c237e095184359e61d7944ad7101f6247df8afe3fd2a2ce1e9b886b5da9db816d2990e2f5365ed75243ddeb973dbe146fabb39ce00f5426909545f87f1e4161b15dc2ae4fec50dd553876d1b6eaadbc5771;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125c9674d86faf70fd0ebf1c3707f0bb9984651d5b8330580952cc53eedbbdfc0ea24e063836daca2c312882b70b17222c0424656d3fe81b6828ccb7f3602b1d2541d426ecf89771bd6def1f4c00faf47a642ef6d9e21e4be3cbdfd5e1ed044706506fae4a5cbc3f13;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140088235c6260035d43274a22311a1073be8b2ea199213a5aa3b74823e02075426a1e1fd6362b19625bc7452ae74a49af903623ae9b8abaa63f05ffbab0cf4cdf902d5376cc88cabcc9c972e1066fb768b750e3f1f05296d2cc08c2d844c532f530ca780bc2f487b74;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b11fecb3d9eab56ae84e213c43d6ee145e39e41f653d0723d3af0d266f9782013a6335164e293523a4308213dc736f4e1e57e3519ae29359ed5896164d15e3170fed50c54463d48b4a7899b9adc0b6908882890d5815763411ea6cbceff9fb1280aaed7e5d13a5a53;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h185138edcfe007278e82760f85e96719a73f1682a5cb2e97ba89a692dfc40d7ab56588aeb51e450b6e31437aebe55493799203d52ae52396c40472d05a6492a81fcfbdaaf862ba6f1a70fa3f91a56a9fcb62cd76a67f6f6419511d8a20f4f97e8c1d1456a032e40da7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1587596c125446ed50144df44f8d2706a0727f52665648e25db79a4e110f790b99af5957c0a0003ba9c2c770884db86e4289cd60d8c0f357a5cfafdd637c3acb8015bb316c8375bbc73564b041f047e6172cb2d5da8cb9e0635f00f602be6eaddd437b3faccbff207ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2124e2e5b7a0af9d1652ff01cf8409d4d8a96acdde1ad880dafa09625ef420fdf78db88357ba9f1bb555a4fa4651a5d4dcc0424c710738a59ecf1ac1890cf3a3d978811be49cb39f3476b44d678c221cc14474c006cc3b191118fbd9a922a334b0f84007bf74bcc44;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79cbfb9349541ba67b678d728977374e2feaaee170c3d85793bd7a75d85e1a2acebaba8a1713ef4a56196a62931ec02a9a53d9c8d741abb04df7e508e7a9d9a1e47d2c3542f056886c2bc80e4ac0032a024e9051d5570420f22387a41ff5dca025c3b5ff454d127f66;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h137f5a28626a87e5c8f861f56b3bce2adcd44261c9fc8249c36d1a9ec54f2c48edd38879a3f1906597f9f9f4626be75e222279e0fadb07f7d299d92d3fded98027cd2255878bf1b79270f29eae7524d0051e5b4de24343e5f49235bee67c5f36da710eb8374281d6a28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc6e26c57ca2426c397a04660d2f51f67bc50d9089e3b212a889c5c99f14a2801edbff7cd1be9bcc21649180b24f7bdd1a70b8b0dfb0fa376409540e96c68235e24074287b9666393ebc48eef954af01c91e0f460583cce9966936eaf92f3c1695599efcb1ce43cc408;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174a84687d40d367a361978efe2d311c9c249324a2200a859bbb5fddda5b0d8ecbee1346dda232d532d928f128c3f95674731be30e698f788902b80fdc791059599046c6320c8e1a5593fb66b01b54a8b1781fb94193fc4f62ebb5b4a21294489175e6dae64e9898145;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7b5579c4df132354f55069b348356b327fbbe6001f7eca41882514310fb0d2a6bcfd1c79abd34ca81acbe171f8b4f8ede112ddcea3881432e0b0ddced9bc3354045c67a633ea84d8820cdaebac35bfb7066cd497cbca02fb8f508a3129aba58af833feec64c341660e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187a6f191f185eebc1fb32549e126d76b0c1587fd00752d3dcf9c8df83e31f2547554a6ccbc531c8f1421cde72ea8b3e32a9ac13c7ded70eed74911140d7c3aac3987331b53dd27b2ea59c82f4378aa2ac76cda72d1806698d989bf9e4796f8c0db441b2a75e55394c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b445d2cc8f911628d0a4065992f7c1609d830589234e860b61388b3f55d9585a681a55eb5128bf4690567193a66a894f8625babd8fc161f9b019b9e74e5992fea40147b1258f0287beffd4dc19690bf608df5628ab4fed1a1df9cb9361823ba31127a62c55240e0c8a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a3aa29ec6cbf8542fbd5db1bf00fd9ce8328bad752267f0bef6893b1c8c56932af78078b745db3dd29020f1e823a0f8cb4fb3f5834eceeca8d1b43a0b76f582b8ef36cb9c80459582e77f6f7c37ed6dc5a7c1bf23c85649edcebbebb03f084c479f1e729ede5ed6e35;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc0a3b2ad5641186c717ad60950eda883ffd90c00b3f1fad2758e2c8c7a11f31dd09ecfc5421a667be9ceec873292da6014877b23c830975cceb35670eebcf61d15738bf5a9db0f257b0a2c8259fd7d99059d89f8e08dcb89a775bf1c33deb9f622ced4e48e14143a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h86d947758fd7981adfd7c0d04b3fa04ac33bdb146b03b0251693ff20c11f4bcb29aab45699df258d0d9c7655597a1cb2e33963d5237901700c7bedf919284175249f7e754b0a1b7b85f81d4d1d11b2fc63e89ca5ebc749e547a47f75abbf018c7fb4b6d7d640267755;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf0b134c8ecc19d88fc875d69fa769a0925479ae54ac2576a90fd37591af37444882156f70379feb917627ec6337a0e64cbd1303fdeea88b16aa7946bc28f4abd0a7eae7752c97e31e88a2987994eb8df6b588211bd9a337cf3cc53f8e940cac2f4d561c530270c7420;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h826c2c626261de8752d5b3ef103013096636ad10690a9517b95d5bad60ee0350a56584dc54f068902144c47de9dec2b06a047cc401d06eddf58b99ebdf451342c68228db37ab3304cbb2377297002c131761928c289605cc6a3c3b23200fe4c0b4f4fe9565f54996ba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc67db46f87235c96b58596216206e7c062591ea93bf71dba541896aaccd351526aa59acbf767b2673ba5f6113d5928cc11c2c6c6659c09c89fcfedbdbe4e149a3a0fd4c0c7d677de3fbddd65cecfa84c4207c1821075225a10983fc4ac96681b240b2cd9e831a1ff12;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb485f0061c2d8adf9bcd0250d183f071514c8ee43a365e0179768c7529fef6186a2acfeee975bc22814c08c488bad8d7821bbdc37e3604fbc0a2cfcb51304ab4f7ea363d9212790d43defb2858b938d52ff3628ed80790624fcc6f235e518ff3e8b181b51ced62a0a0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5a1d948d4425e1ffbf52671d581cd399e7b545252ddb065d3007793ce48bb2761fb2ef268bc7c4194084dda8b54c5c26a7e28b4a08328402ab7ec491389cc80b3a203a1c62a78e1c0279aa91067e71b62c928716f30c20ddfb8b538de56830c8084cdc4c42084e57;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hded8b2309dcb61d328a21c4f1c382e06811a578ff8ea58faec87aee42dbecdf2414df8c4d2fa407d5071e95abb13260bccf722a95e6d5a3d8b7988baa4f36253da498fc80da1dc275bd56768f5cf71fa4f0444a04877ea1c5ff21eead4721cf99908a5c00359296cc3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1174d1480ba537f02b41773dde858f513f18a9371f01cb8dce9e041af11fd62c66dc60cdcf649d3f8f28ec5ce471cbab9ce33a4a4747aaf2d2d343102e04a22087f7af449883882c9cdd0682657ce5295e672b1ea918a1d2db21b8333026dcf9b8e6e4c972504625d0e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec0423fbef7de7115e2e8adb08faabad7767691ae79ea8c1acad7f4e79b388e7e91473f90590f0f5c9a9756ab0b1a22d152d28d33539400dd3ad1ea3da088584a460bfcbe030a2441b9f3f8d60121f93068b88f038d121e7a1595eee2a18902425d6ffb733ef31655;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1930227b1478e6f254892e928acd77bd70701901e3763d2550edba672b2725b35908858b160adf7b135189b90f97da89a42f207602b0e39e3c59990ffabb94b36a923706d67607637fbcbe49153022a2f4d801c37b341102a71640f2bb3f48305b43ac465ced311d244;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e738082114d855a3be1ebc96eb8d7c4c4cd9de2f30af53bab74ce13d6466fed5886eb37d2966aee4e8742b93f37d3de5e6c54f213b4848ca44698f4e921097493d3e210806dd4822d03af8e8c18dfee3a65abfcd6b09aa2e408bbbf617184613aa0a1311053b67ef93;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16d950602222ceb1082a58f68e4131c8694a834c8d2c5b949d7bb89bb618b491af506e838fba7e3917cf570d6262c3856694f8bfbacd33689c81b781509d0c2daf5aff335b9c047a3502c2cb9baa59354e828da221e423b9263d59bef4deb7bc57cad7f586bb97c33fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5588d911ba9a5eb0beda82bc0c047999b8356d526b6f74fa2ce662641ffc501c6e4fbac0a9c711730f37b74e7856338a6202f85d30a5e6af33d0b01e56f994ca084dd2d7cbb16a21d1f74d95f5c2536538d5737967d8f74f5815d2ad49992ca872b015a51ea8e28240;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h434733cca621f0ee5268dacf47821567184cf8a53f08f25cfa55a3b036e712ffeb0bcf0bc112dccb18317eacd7503934b7769777ab307359cf48a8687555884b062abe7481b044209f1c780fd11097122d29866fb37db362731ee82db61ef5f521a8ec1b64e67f4862;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h65d18b5a1e6400dab691734c1913a3661358e65414f60ba28451acdddeb2656351b517ffe9c3a6bd264dd06d75b20b6d5dfc3d8cea01fb999b4b03f80a3b541a56c610c327a5ec385eebbd9103808c835d0a71d8bc5b2718b6e9c548d749b6dc737319dbbc1cccbec1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfaadb4ff5ef1a7370347c493d5466aecccf0def92eda73d66d2a15730394c1d21d94ee3f131f743be24d5d2022c26c7d505da7c6de403efd06ba76a730be34f7178509bbd2d3a0f51577722e800174ef57b0a28a8912a002cf119e5cb197f4a3bab1784a6372b1231d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h48f51048bf4ee1725b310b1bc397abf43c634d0ec7676dae9beef76e7d3cde6fafbb437e63b1d2b3ae000273a62c3d3b2e5bfabe473f6ea2b7637e4b2ecb9cce9b1749eb743a8a82f5f40fb09cce0f35f55b20db680c2fb37a03de284ce5e4b7d248dbf9f2c5b022d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dcc39fe8560745c936c0e7d717ca2e6661f490c428eadfd6736f5125e69b0a0f53636502d34dabd1fb6fd3eb2986109b236a4fb67a6a3fb7e5fbe3b9e87d457a23a45a2aa33e6c2142a353f24a58e05f7a3baca88260e8eeb31c4967634fba48f9ef193ce32cc84778;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d0b8a77fad37c67649b8621622e2f5a0df336ffa5d7ed23192bbbd11d60d483b7c3e040fe9c9f127c515b2f51aee7962f16dd0797fc9cd362348fab8e94d1e89fe088880bfe048561ae8d5106517b857f5b2282d27870f2be3f3ed9f35601454f71e8b39c128bf16f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22bef70ea5fa60ada29711df538cc9f8769f9a58e65896502d4decd9a079515b1c306e6c4128d22f0af688642bb3df45d38c2a95c5fdc7dd6b02fa63de61aa5471d1efe3aef9f9bc3c58701c7bbecedc3bc433069da457e2c7bbbbfab389dbefb0d53995f9336a1496;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbddace17bea4e01822766d3f009b8af4a125dd308b6fa09de0e847046ffa048ef6bd3fa8404491fec5844fc1d3321deb323f4d0a046e7d873575d469b1e1d7ddcde0852fc73d9671faae365f3610bb7f2eecd89f653d22a7e04d1094d6e71a1a5fb1decca6ecd78eef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16270c7a8a1214880c848b4ae5935ecfa4fb9954921d2d3c45a5508c124463be36b79ffd89877356df50554a775ecfb278778fbcc3874128473f6e094a4b0ca8b51a1b03fe054ca993788e005ad677a9c324d0fdef3ee1465a4fa7287e9d8647b522bbc82e708aa7553;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1dce28861a14a68ec07446cd4ccfc6ea674ec2551e60b2053f84fa116527e89b1879038fbd2a15cf41a1124f844a896ec3dda351046d0ea906fd98aa147c7fd2e2f12267d5effeba01cc05ab9f539bb91aff3d9c4aba3861f670b176a6baebee8873f1d2d6052ec72;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74e06f9b1e3e20256180942565d4b2024d0d32e4106f5586f205849dba60eeccc482e4678eb0b7aa192650ba60f31a251c32c1e19f2e5b3b76383675499cc423c32b0931c62a15ca03f4d7b65661230242ef0cdbebf33d18dbd95eaa17bb0a3b36102b3a0a90a348ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1235dc0f0c218a80ca2be59e9f79397eba8c307fbb45f5af1a862665fc509102575e07c616557c2c3451fc6ad78db844e00875a5100039dc655cb690220e8ba889e8885af88bf2738e84c08e83872ba907248bf2ef6da379851aeec345ae1975666ce0865418677644e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13fffce068817b190e79b7ecae01d8d7663f35f99afcd1becae0731615a14cd6b57cb017407931eb1bdbd8b844ca88bf60245042f00ea43103e6489eaa1a89d24facfd5534a9dbfffd0523e802ce839b0c7a241fffe8492eb888d9095f859c1bd054b990a2135c2c0ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha65f565b4770de638c1ee096995699e7f084947a953b3f1beef457a40f6e67fe62340f42e6bdff17e02703d753950c0984f927b6e7cfe9643ae3f23e14ca93889fda0bbb7906c33c95f26ffb10bbce464fc85e9b386213294aaab7abee6aa35fefdc55b4a9f370a9e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d676cf6df673dca4ec846817bef83338103e8da7ecb69c0460a1af21ed8628295e5988fdcc81ac10e2684ffa5ec739d8c502454de47bf5534dbf066009b41d1983306abeb476df224d2fda9a9e85191b7d0b3fbdee310b6f16d4e01e6188ac5e1d62a29d4777f812b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf606d5870bf0e3ab6a729ddad39eb72d368ffba5d130670bdcbf923701aaa9785db8d0bf06055774b33925b344391a25d4a5d99f5dbfc7e76b4d26a85a981e3c5493ae160d2047205eafeef748e9c18879b919e08dbdcb9121650c2461222c6ec411d77a80bbc1db0b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd2b9102e1745ebbbc04c850a75121b05be3acb6c6b397db16d620552b43c3bdf9ffbaed7eb25da11e5e12670aa81a8105c17950b5ff513b9a6bdb236d61e3d7095f8fbe08ae6b374fb7ce7f7f520ff3edc6bb4d68982ee47592d500b2d2b973c3ae2dc8617117aabf8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4d896867a19aec63b90069f94ae0aa2ff3c32188780f969caa775055297f109a68f033903c274788239a6c379ad1b89585ccf11b4e5f302fdeddfb678fc0d2de1c272697b1fd12dbb809466220aa1d589d8b1fe89ccad0c470bfe99a6167c177b9563a10aa83f2ce5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdbcfff16fcaadc10f8a7ee04e91c40305e5e503558924e93d553ccbfaf5a018c6c28ac9322302df8a021a9dad1b7c04d71c0c44f49da1574f5f78a8e2f192b9a4036c85bb64b76bb76436d4aa8ddd89456a906b7add7a11cfa4f261214b6c9f4e982ecb064b09e143b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h32b921c90fe2a8f82697d529761ffb5fff4648714958c08f87b301603578cf379c29b1e7ca6bc7d6c705686888c0abbedfd83fd3b9963b1045db08a864af19562cdf97ebb85d3a9933b011aad506c13abdc1782efc78b506ba6705b9d252b2d7ed10eaddd31c2ed9c9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d6f32cba9e57259f000511a43b627d457c9cfb8023bad619da90279676c99b4606d9f23420efe30503c1a69d09be8a5f87bd6601ae47cbaf6df9efa8e7339e70f960af493f75fc16e5bd91007841624c43c8b4e5e5eb2d67a1dd5591d4b659fec8cae6938c640347a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d675b43d53ebdabac02aef0ac5c090442bdece1ba545d83d6382fdd61b3732e60130b04805455018f358f6e24fd4db7df1d7b301dbe0faccc62564255bcf4c3b1767fa6c706d765043ee45d375260333e3f043996f79d05faf308c10c284bae277381f3af5e6a1242;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8d19d3819497f9d65ff0f0ebd2d3c9808991220258543fa1a3ea5e89b75c9efc44acca58027eaf072719300402d5e9fd61b2378e260d622730d965272a8c087bf37a5466e8905cea1413c1d08a6c1000cb967a3c1d2f6247386a92c0710462807e097005305da0b95;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1afaa49796e6d13bae1632b037ff099dd105dcd5818647408d41fb71361b90fcf9e500166a2686bdd3422d53d430b15e59b888322e821df472917b55be8312a272d13c966f376efe41cc87fc80518f1b9b1e1a7c8c4d6df9519fb5bb7088fc374f0aee93a66e46db722;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc12393c818a80e692d71ec20d334247395833bfd52c33372a9d618f0112989aaed078392b5153f2c5fb624f93662dd668dfbab84f6e47e2a6f44e7ced601bb7c41bcde9b26669dfe580a47ec89847a2feab79956d3d456aeed9403d977fb22b1673c59775c82f12b7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a44d946858b116a985de0f065198b17d9df0c79f9ef51894cbf652c414da1947bc266258f04642e706408eece82c967fadb6cb76c7688ac651e83096973ecd09a875c10718f7d3102f0fee617ddfed1623debb717371456cab1b5c51a4695e1c3dca9e563318ae3ad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c9d9f27af9314e9dcb0de1b7298a45e8406498416ef53047438aad879a5ace3af1e6133d89a0fe3562262a34e22b9315fff86eb13f6d17532d226d677da498eb766ea3cefb43a3dbaabadb680642e09feb6b841c66f9c2f94fa55b93e9374853b4581bd940ab998de5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140a59039128ea707d7ca1dc8f12978ba54f1aa5758752455a10ba9d2b785178987a1c2989dae591a44d456121a94c24312e6f6bc264e1ccd2d78de689a6c607dd795a6b1ffcba274d04ffef4d7e340caf5d9d5c300b195c31a931fd558cf53ddfd4141a0511727c772;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b66153be87e0b7c0093cebd09b9e2ce6f6ceec7b77698e608e0d82f3d71dca1231904fccc9649900fbc1442e2c31e21e44e26f43691d37513052366eb9abc27bfbfdf80c71074a2ca41ce3103a673a8f5ecb2769d571da4c921a5f9bf199d36b35284381399c0fef73;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h622abbf26584641f681ff472e6e91e6ac5dab501b79e061c453eff46af8f21942c9cc957ffd7367a7f0efbcb6fbab33d94b919b051a724c9a2af2eece2fd472bf256b47b4a26a77fd7934e3741deb09a4bff41bae9bc8323c4a0f16d34a1e2a9baa353fa919d0457ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc13bc7e54ca202e4d4d3910bdfb765e0c55027b7348b48acdb8b1d3aa91d7cf5cc180750742d3eee798c6b2869259daf0123e43fa49fa3c939f708a4e8fa9d98d186af1301e430f7baa7911bae703eb3f81939c9c837bc70a25028f3d23f9605f9c4997fee0cf04246;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a3a23ee82878a69b5e313ed38b57f373365dd3eb57c70affb41b49692dfdb52a5917b4dbd609cc04bdb7f140c2f12e3a6a92b05c2778d2eca9c0cf6351775333d89005aef85f35b72fd391762932743721f6f01e572a389983be2f17c60a710c163e26f2d980200686;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1729f4ac7715216c81746db3ef8f7f14a4a0248082e842a688bb439f4657ae2120b6e0d7c86dc98cd20c8d8975b6de220c2318c849970a76a5d65430085965e5b045bfe8d52f6a285bf50b052e598efb02862f161745e56a93338429f95181375a783c4953838d1e128;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12057179584e044139dabf094b95178231bf5e1c2fec5e9849e68675ea5337ee34a44482b25570c8ded702aea942652712b923788057c703a8d9f2ddb4e2381edbcbc9920591353a7d51b0bd2f5f64d5a3f1352f78a1814e051525df09f4371f4a07db70f81fc610cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db91d78826dce6c294aa48894d30b02955745147c95d7ed2415cfdd9b70d8bf0ca4fb541e22ad523026c0c1b5adbb8635f09094ffce8a1c640d614d181b3f3d0e8688debddea957fe0324d667915677323eb81ecc2c61117cf3a43d6aaa3b89883afcf94854024d2b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hda4d7e7031a54d4a0ec38adff4e02be390ad15de6f95bc32cec010f484f3399318e749edf325abc8f10949f20627ac4911cc3ebe54596fc8c1ff7fa9601ad0f9229d8f09b97874e14a3c3295abbdc61ced44327809f5469f87eef56e6e5f34aeb59dd9977c7b01696b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb3848b2f9b3c4e9bc6efab39b8534b189f0769e9cf281a321f930e52a082052389d12701cc38005a7916aa6a5ea7a7ca4cc673061007c6ce3684efee4da473964cddc428701a3be02299a3ce276009eeb0779c94ece1e6b0f6a701820c046f544cfe672feaf0db285f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12bec424e183b750e4a64fb6bf48acfa878bebed81e4fded9cc938b4fcac96244966b3c5b14ba14a958de66460b8eb931a8077d5ff8440756e51e90ca8d2a5602c3b44c304a54a9195d2c65f6d4dde1b4d3af57e21db995d2f724ee4117d170c511d3f627c18a8ab754;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17340a1484d8b16d6e3b5c26855afef9b9e88692db2a80bd7d8b8995cd7b7eeca51342e5617f33b8af9ac915b0835771082396541fe8b5bd40416304a869a07ae4edcfba4f25670aa3686bd173e48ea09b8bf87d9a645766e4a31b85b42352d57b36a7f3b4e07bbf58f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd13a877903fa1770e69418bb47004099a3f8bdd5d2a83c1348a24978e43bd7204b9b46eb7567f1d7d471acdd7384300692d1124fb2dfe0beadca1a0c568eb1bbc610a7ff74e770432bca828138d40e8b274a713411ac4e8daf72b4d40326030abd432b6bc553508a32;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1483628f153c9a06423c10921e677f86777d49b17e8558b4bb9bc66abc13e995b54d083f5613665f1871c6a20fc09d5d665e3ca456b9fd041b56ec41d8de7f9d44a3b3342fef479b1d4f068a76fc290a5958c0262f46420229682aa994151200af35f5047061dc3ce4b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ce9b17f2e482e8a8c6b98b959141a06c880a209eab4cdb04f62631027061cd4c7488bc8a7289cf4fafba0daaeccb20dcdece7e1b78462f393e44fe805f4cef2995ddfac68df888f8cdba784d2b231dd3b493486060c9a1a9a4e31b6ef096aaa40dd7bb30ffa7299956;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1415beb304082070ecfc04524c1b47c0f09e5bc0246a40491a25874b1d8b8f65afeca9bceefa00ac7d6067202bee2bed726130f2651528344492ab4acc66ff39b26af1776fb3f856967914cada7104e24216cbf3e23d29959e83212a16f904dd78095b3c038d6dfdd0d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8dbdcf79b3e34fac1e4f3d595324fe325243087838035ef259f104022a9e742e9d33dbf1fbbb4062c01e0e8e981c357b200efd3ab08b58a01ce6eb58f28cab3c64d0b6f46924f7841d4da418057b1fab2665e3e5629568225e83264b3b05e59e9b836a3b4a8a0bf46;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc0c72334bee411ff283dcfd11c1a11f2fee412c6bd2ce903957f75ce99896d603502157491c1e2171402cbf0739c57ad83a71b447f0b1ea91f775784d8b581aadbe2c6245e27766cbc21e10ea8003fb023d1557f91a3aa37f1b7bc448daf93328cff88df708946f027;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d033888c8771d4bcbcabf3b4e56b3cfeb01a2063f4eb157e2d6d81462e4b41dcabe154dee9105b4c4543b3d1d5cf83eb25c7e7bd16e669e7bfa6f43f1a4af98aa8e06a60711362c2e2e1ef8d852300e6805d16e1e874b5159ee1584def9249376bfd4a65e69186230a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5210b1b32e671aa4a495f3aa7d28e5ff82b4bf312a07dcf4e68a9aee11b534328d9bd4ae88bda6157b26d5f8e3e35b95c60aa6326edc816b82a13ce292aa3c861d0fafc9f488fc7a0b35a8f2f5a81ca8940384b4113a43033d269bdf89c9ae322aa3a680f079e2191;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8d5353f3645ff01786851704b3ef415c27e2665e44473c1852b5673f77c23873e6b3e6e300b7af86d4fd484445bdce03ef601e305f5adb8376da5af99d86f2b0f7a160684a71e99628ada30b852fd12a292310ad68a08e5eeada4a3ffe95afae23d936d321be41a28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8bde6d3b0550adc221ddb8f3c71cf2b96c9c221c4734e161681dff71776df441c4fd981b9abf7796df7316384ae57474fd7997d68f2589d55e84034a1cf7dd8aa3bdacfc40e61332581e33edee1adcf4e9bb7f13000c14465d4ae9b21036f34fc39b03da7ffb91780;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a21042e6ca2f06e807f4582072321e8d2b803b5587c446de4f49a801bc757f0eb160ce4997d6118f45287359029c12693a878c8c99a8bb6754f9dff0cd3cf1a05e60dabc270a6257584cc101bf9d3bcbde240dae5a59e720d08b4209cf6a7f2a354316faa037db29c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7e74e26ec6eb2143aff12901fedcc9a329151755743c4cd9af04482f2187ac3fb28cdf0e56917e913ef22de15c8846d60471bb295d8175d3fef2953352453c527d87cb7547c998267e80083bb11095d2905f26f4211c9106f63cf44b2d2ca7f9023fc5f611e32b4f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12bc82a32111e7ca3289b1f41bb732c87f112474471b05c0e5dd52d77be882db74985c8783208d3690468a405ef2cdd28322f0de7e851c9fd070fab6c58d412e9f2eb646f48e41b7670ffa7e16e91c8609e2882dbe84636eebb0de11f4ec2972d92b6b97bc96b9663dc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h152059b1e87f1be38b779cd656f0c3536e1c1ae9a5ecb4c7f8d20452af5c8b8c8ec80ea1f954d7680f373004af0db20618983d28c2c0b4be761ab617dbda1c568b56d14660897fa8d0a499f1932a18f13511d151977d457b96e2e8818240266acf235cd0cfab77dca41;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174b0c6a47ab6f00fb6acaaa3355d8d4a7b1f16ee208b38f24a1cb2aa0d54e42904788b87676c16f1b1dc8b9fa5dcff632f6bd04f8e34b6fbefc6f34fcdcca213b37d7193249d610c86fbe209a2e265dcc044868a77f3c54adc86a5848370b14ee95cf668a3882bd170;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h394a5bfcac0fe90834b5a3ad47f48b2f01d609df1b894d845a0433b70d99a769f50bada51b87656ada1d94b1fa0f0cee85a0ace7927c14c4d9f484d62fd8f6221422cde14de416f1d96331925f0f773df0fe634dbb82296ff3ab9a0a38b0b2095e16bd1b25014efcf8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e01e318004fb6cc3e19a0e311d139b641836078420bb2d31d5ad86a431289ce055717fd7f9d01fe746ec53a57035c2106ab573e88225d3ca231adc1f878f1d2c2867238e6ece101c9cde03381fba0714200cac2fa7727c1d87613d60d224f0c2c47c8d27ce0222838;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha6611c6f510beaec3cddd836a34e0e9116db6eaedb00be9d5b284fca937a7c2f1d3a13ae74496daf3cc9f722e0247e7e4799d669442fbe57e23953e608a00443992d30f3c315bc6ceb1f83ee3cfb849b812f4a4091423c3af01ca64c6ed7e3211ae95d5033def48f74;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5285f10f0e0ad119e972c4317fc4f46213a27484fc789836b864a40939b26b7c935670e359498708eceb53f23d204e36edd6720a7a3ab64cb77eff007d3bebb42d55bcbca7f79c0829c0d75990a9e70da53317eabe0bc029a9e0f349487a3ba3cb8fde92cd2155061a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19b71e1f600563481356972994a3224f3203f06f8b1c86d418b6c8efe994a68272a6d03634124dc70ac5d2901e7a65c3c89dd04db3860db934512e8c19638876eb51dbdf43dd8c2fb38e51b91dc69b51defd0fa457706a124b69821a3464686e6f7f2e04c6cdd140ce2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha16f1f89e6c29e9469b0fadc5a6faff509cbd56ff0c64585127093ca2cf756038d101fa99d28a92d6f0ec77c66a0272b5b8ac46cb384c82c1cc20f041c305af400024e9f0391c0711cc2ba2e58d580304017671bea23f29f07cbb8401a29dd257d3cd021e3ca1767ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f6ccf395cb123dea8c455e3f5a7b269e892ed84aeb40a598670fe99c4a007b70710c276f3b6a9dae0308bffe6460afbe714c07900ec447782d8aa31adfe6865a8d09f6d75015fda8f9fb5a6694788688c871a72270c91a4d0092435c82c66e577bf2775e617eb45af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5acb8ea7e60b7af8c9590504c5957b55732344a2817355814751a81b0264adc4b20f8908a892bcaa684901e9386fb2ed459044f6040b7436fd9b157a36e63beb87da9c520023a42e49aca99565dee7949dda273e596b560546092a83434a69a980127b166d65d3398;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1258025407509c45a8ea3d9001cb80fbecf2c00048a8d681a6a946f0e7cae8b0da3f9293f7dad868169ea471b913ef5431606e34cebdc5aead11ded48401b7539aeb13efc26f5c761de3bc27d33daade9eeec6100cd5a298b0bf9d22be7e6f0a6026b049483dc134597;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a28fd3169c15cd638fcfffab29628641c43a4a1a53e1d74e3add9165e6c5138d3a239386116811180c659c7cea37ae5ed07315486414d06d7e1ab90b7892b4420044002c2cbc71c1e1ac128f8eab787fba40a278bcd4efa3be7c7628521739b34cc795f2eab586e254;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8aaa46a1167b61022ce4bbc971fd2fb9d45fe05fadadcd137a9a0c0dff970e75f97ccf0a0139bcbc200251e5ccad2205459dfd2106858a148e6852e467ed1a905200f47a0a73c760e63efa0f3ec7b887c4c2e0334e337c8f77c3edb931a17ddc331cbcb486230d20c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8d3428dafdeb1d633e8294495135032dfda59ab7894ed36831ab55875ea2edfb850e956ce8293d43d80e5511a9aa438d0cdcd3132687de52930f99afdfd0568f2b0e7c9a7de354ebf60c3c3eb73c4967d1e4244cb59603e5c3433ebc50cf685e94617b56724310d0a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc035da317755164995c6acb5792eb5cf1642000d03daac810279e1d902decb1a1d53844a21195a0a57b177fb892666124ca31aba5e5277512241a5605979430d87fed824dbb84182aac797d483320825b0709e1b7b9a89de2f14edcb666d097a131dfc6e917961913f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h180e4a8995637bffc2c8b8237822f4a99e688dbb4c7daf936363790a80f968b35bf205fc7cf4d0d95176b2b609d1342510cd1bf4e3600cbf4b642aa139e356473a32c9c15e94615f6d9be07208727e01cd7e4221af2574310c6426ea9e6eebfe0e6f2a8096796753cf5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8d190b3c94a01f48ebb97f161b504b056259b802a04913dfc15f8cf53d2c042353b6e80d7588a7f0df498b6f8972a739d56e0594cbb600f6b0692127477f823c4a8c7db3894b5a4e79d5824b5a354db22bb1aa9eeae13ebac356362b274970a2123f8f4fa04e19d91e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17425043bb5145a6e7203579064a1b3b9b1f35764a8cffae8c5a987797e929ed87764694cb493de372234cc38c29b728f3b0d59e3e57a28c908131011cde266793d0e62da33b9ed969c543dc3de3e0e05fff3cdd69497d9ebe200a5d02bfef44ffc1a482b8bfef91414;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e383de87a2075e47396ff5992e1bed183cb41e9b7bd668fbef797f72cd7a11e4e7b318be53d4cd17f425fb50a6e56531510f96deed4e8eb968e28a402a20f463154e9bb8afbec0707a70b1b4f7eeacf597a2a33c4150238a62fcb35b78c738508cad75f521717a661;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d13cec6663d20f63b74d59af7ec567486b735d0fbb1f6629ffeb2d42b586dfe97a6c3ebce2c8bee3d3ff4d46721bd3f3756187b8981a5e53db583f0f5356390298a56337daf4a72b855d792fce9e36cd784096fe07a78608b2bff882321478d2380744d67dc6e683b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h771e389cb85598c3f46b6a136513cab231bee4fc2e6a9e798b4b4b87592bcd9dafacc95a47beaa9213087b640216b9c4b5331f8cb826d031961b3521645e0a6ab80d4169a3c431cd964641addab67f2f5e72dfd54d7aa8da55403795d53d14a7c02c4e8a992573e23e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h106a1699bd518cbc205b8fb3c0ec306388db95020951b6787cfefcd737a465f60ab71c799e2c9682495222888a59fb45b14f0b5758f5f48d981b94aeddc68b6dd12ac8db1c0f62e5126e239a7a0e601be0ecfb07c8832b1251279d002147fa075e209556909ee084289;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2339f044737313838baa6a23fc73c3ad8b38f9c635c8abcdacabc613f1c1636ea702b2c0ef1e9b5f65e7bb2b7510e4e52215cfc23b9becb7ec08a201ed0c60c7e0db1ad75c00ee83942ef457e93f53d7bb86f1a19272c8f3ae45d6076f2df8c6ebbca3a52fd36f7c8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7bc10a64b4507ac2fb56f03064daf0af17f732a543173c18f7e2756d3e605afeb26b9fae44f55748a9979dc7dbe2d1cd4840342a2090bc20632a2785bbe2e485778082605ea83143f0d6aa6b5db7f0004c8ed83b239d729f5ea897271c99947af6c7b7177ef0e74d1b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h173dfa0f851ddfa2addaaf099ed9135b10e48aef8ce561d0694fba07665f26337e3f45b41035118a2dfbeab17f7f092dbbf8e5158af45375d8bf17571cc3c486517106eb3158c601c89d43e0e1a9ef0bdd7e7c040cfbb95bb67c419d5082686be57631e9db1624419ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc83c89378af4bd99aaaf94bc7796e3841ffab5af16d63244d52edbeca42ed3d9d70aa9005456852a21ee647467ae61cfd7bc702e2d597e8353f8eb25eb67979e50d8993c5fce90956b34b77f80e17cf53686b52ddb868de9f7a0c8a28342d4c7daafc8f0e683d089c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h39b310a29ddca4cca15db680bb9b6a293d7e860b9ce2e03155231eb1816c6d029b8f3941826469f8c8846af8f06001693e9ed36b9197c822a078ce4d6eb125328d0544da20f5509f2a674dd78c3737e443c8577c6c9b206465f38b0bb90d328af6ccde184203ed3bd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc947cc366c0f78d011d837845aa0ef8235ed410cac21192dae75ed64db0ecd4775fc761df6308b33654b409c84a6895c663f3e57c18124d9140a25c8c8fa70bbf27cc2eae339249029f93457cd4c1f1ed84e3c8753d94c970b09785907ccdb3595b8500628e0b49587;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec7f41b96fe8c4d9c3b6f489c38e20aaf2a785fb1834cab693ea72d8f8b095a84e7fdf57efa032f54b59ff5f341a95f7f0298c502dbda7292421d9d1b949ced8ab3fec8611249f46de57068a62c5cbdd8db14ddec60fdbc142ca3ad8acd81a3281632d9a26eb81f5d5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b011b08f71030c169f9bc3f4f093db43c450c1a7d0e097cdaa3567690417f2879e46e7b7f3401b8dfe2b52390ee273263f0768dd03d0a6df3fefcf628e646f55543a9af3deff4800da67e42f9276ff7be439365d4079e3ed4ebfabf867cbb02ee3dd4bd6cc1d02834;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1721ca320847a935cd33e15dcd5a9dc8170bd2d2d8bbd1c3aa18c86d25e8933f2795f66f1b9ab807531053cc018b848fd430c790c25befbadf88dc296930fe13dd575400f7abba085925f77529f440b3eeb7d22f9323ff96083f195123a0cd5bce66c65e8959be9fd0a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15a1944efda9c51b24f3ddd3e83eec223149135f21d1014d6aff6deb6878fbb84e26040d23b9ee67d7d0a0a11bd956e0cfddac07a5db87a014b7eee6ffa3844382c0b80e8543ed049a3bce72f2c504744a85e8b23f945291faa90527dbf837e47b642965496c4de44ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7161b9d906a796d74008b4e1d9c89b2a6257b7ffe625bd072c202ee0630efbc7c90f08d608c8ed9196abc1db5998688526c2f97b53bc4f41168fabce2a6c2ca945999168edfccc7803754745eb6612d70d73e8a89c569e7ae189d9a1a246e5c1a97bbea31a8419bec4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbba37ccb6ab1fe3b1fd0037ec333212e81eb3343f3c35771aeac8e42ac90a75ea61a2cafb111c1aab4f19c56e3bcd535366c0854085b500ed3f3bf74801171488022d4946fab443834b837c2935bf56dfa4485ed0cd4f407a3fbb6f01b90d22ce6edea67c184c070da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ace143fd1bc69a9b7108c5ec75d5fd6f62ca302326d17b69dddafc1fa3924bceacb0aaeb44f852c94f1bad6936909399e1d7381ac1513eb860f3b0398c90398b280c41d8d68c08072d9f046b5dc829e9348031b094ec28dc39dfa3e0c19e78e12f050ae2127b487a7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2b111996d82a453094036f2b9fb902de7331235e114106d89c500bc2f97376f3f1534642fa0f44f80ca0d758f251de3dd4bdda2eefe60243c3236f34a28a8259123c92d650ba0757f2d8715d0a11da2c8189771b5335c15fb419d6702afb3ea0d866a905cd2d2c5797;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h205904e8f85104745264a82217ff07b222c89dfc45ce300d92b495c85cecf72173ddc9b1f52eb7dada2c0060695fe5ae45c2516dcf43d52272d1a820d4a9f90d96019b701d39a56bb05a849397d930ff377c79e7a79400a96ab9346f33cc09775976554d6a22fe7fd2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had496fc1fdc1ef30cc7364b791dee4de5d79424a2d10093f479e6e083aa997d5b06485c6aec8d2c5882f0569f9f6d3bad010a5bae844d8db9fe684f520eea125234a41852a5d909eae4f9f8e4508328d68aa4f614b30170b94fc5de6e2b1fce5d05b51267e1ed1a6b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he70ade9b52c7277af78b7d3598a597662421d768c2367bbb6085c57618f1de1553c649e1f016b2c04dd6e5937c7767050cf9aa79fdced38a0b0bcd4e9b53ca2bff757fb5d6d6f79312f137afe0f97435d256f03287b2f865ad7fe97606c7ffcc385ce447c33a00010d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd54309ec07784ae66417097d4abdd124b1907319101777b844c1b8fef19cad0c6badd12b61f1ec37fa2e1dee53901c2d80f45e5dddd89134653cd22abb1bd90b48f404dfff54cf8ed43d5ba52e401200b4412dd46af3fccf40025e026809c90d6628737168a0f99ba7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19da36c9c2e65a0b44a4261666f606c45de27fb41266ea8d525f44038d744a2eae0fd3525fd2284de3e24a419a26aecc8f34bce9a8a7f9da0a4072c92f26682cac75f6ed846e85d45e07a3eac5c33150e07cdf2262fd0222a5313033b014b2e80e9edad2a9ac370410d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1faae28f7618937f9d46574a353598d6ffba726fa61afa8fab3ad0c35192c9c5d775f5ee46df679f0300aef9aeb8a8fbb1f9dec487a40330468ab66a6dd177db49946e7597333ac50963a0884092ee4819c63ff4f60f311a1167464cf2e85bb47bb1ad5d667fdce4b89;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbca594ba14a5b784d30547f62c893d125056cea57698a1eb6a6ab62146d6a180b37db00ef087d5bd7784f63b6c6e837e70a1769a6e2b85f5b0acca7197fabc9be72b08417f731dbc46f651039034ff8e24a7a7e1868c9f965aac5aa4493531aeb28cc48de098958882;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b04e30e9da3fffad4caecb093abfeb35ffc2a3d0ce74db8c88f12e33f855228b1a1022d9dc11575f7174df66a83baaa55e0cb3c5c07e40dc61ed1faa5604d5a6bdb90a5798d9894b96d04020b23004ab25866fc2ecc8476873c73921d4ac7adc87ed4a3354b389900;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha65672f66e81b3664eea6b0928b01bee9c79b9c4514c6072d3f29513f51618f9172659e7d5655efd3adc9de30c304db9f3c2e0eb15040f6b38b57be59898505779fc115b3011de975e157addbb8a6bb59232addf96a81153cf0f0f04539c12c23cfafa69d5e08dab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5ddbf961dd98405c2500fa3773949f0909b65742c79006b6b9e7e84cbc4e4279389fadd8f67aa8d948d4107e8cc91b19a4f8fc728a263d71003f44aa9cb335dc5aa6ab0e273eaedb8c82e47286ffbf72d37f762916f578ef030d7f660feaa66ad96f860dd740aba14;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h158b0df98e19d832c9ba6854b5966558aa2767ab81b7d984dd067daee9dffd4681daf6679e5252e19320e80515206a9ac721b68becb971b7b1e64d575e22c376dae1e88e7ba9e0de97967be37a5525b132f672ab17315cd136262e64901775c86a1a71831a0a8eaff3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6381b143494968bc1425f8563f8c66a04a647c26f40cc243648c6450a7aaf3af0119c7877f1983f91131edbfd05e86ade5b46ed407203a25e6dbf6bc6644a4ad6aee0bcdeafed48a69c566273d1e72e1e1df0a69fc5d0baeb51980900c09e8b25142ab5b022f50ae31;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13c5a1c1a2c049be1ba8105194ab05c06187a3dd51ec169720fa8fb34f01cfc8403d291500bb2367c35329894ab3db5f493a284141c398f3335e35e132374cf1e04baef77abf9fef70c84df1a7d1fb85284bcd6eccd0cbdc85feee9cb2d6632d6e47650f00932989e4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha319a72a9958371cec15724b947f57e8dbba81aa9f96e6dce217d1e4a4bae4729bf7fe214ac2567418efe0f88a85b8ebd331274522703e4a1bb7a5ee28b481532214f42fe93708a3746ebda4a07a30ff0c26374b2e6cca30b2e3b68cae174a59e0c9b36be861ea81fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c14c9f1e73018ce2e76006f8b3ac85f7a53b281eecfb8150a204dd8f4c3335cd4d843c45c7e58744a82bef486c648dee3854dedcf3e9cee3f1514b1ed1dfe5d636621460a5ce56a545c9e40546b7d04a74f0f1aed602f3e19594a9de3906f62e76b6e17fbf3125b624;
        #1
        $finish();
    end
endmodule
