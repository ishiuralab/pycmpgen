module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [14:0] src16;
    reg [13:0] src17;
    reg [12:0] src18;
    reg [11:0] src19;
    reg [10:0] src20;
    reg [9:0] src21;
    reg [8:0] src22;
    reg [7:0] src23;
    reg [6:0] src24;
    reg [5:0] src25;
    reg [4:0] src26;
    reg [3:0] src27;
    reg [2:0] src28;
    reg [1:0] src29;
    reg [0:0] src30;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [31:0] srcsum;
    wire [31:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3])<<27) + ((src28[0] + src28[1] + src28[2])<<28) + ((src29[0] + src29[1])<<29) + ((src30[0])<<30);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6677c2efacada86875acc5784d44505bb8b86ddad3d7724ec2187cbe8c265034;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3376db151103e591e90826b2facbc0b227c9d9564412cdcbe7afced4a6cba084;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2006d7a5acade56b6314fd2a0317327bde147fb8a8e2d8987616deca9afa3f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4ac403973de07f510727fdf0c63adc9a6bc1bb28432ee6433d2f5c7d6e644e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d1b70420d5fdf7f70c975fd45fc09ef3477f63a5a2edf6acab9af3e91a7787b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee43e1ba562a8d11ae880b64a75a0a13bd6220d456b5356a05582fb2694c165b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17f24bff135fe7f0ba58e7159d835a8a53b23e73c747caf168e20435f26c159b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c036019cdcf8baaeeb5d1f195f98f5b6b823ecc0125a9eb413eaa91c1fa1e23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9805abe3ee81a3c9f1449e2067e00b3027fbc69f1c9e84f3f934fdd7af535426;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a225ce9987e74ab30b9a02ca8a4c7b36a6b7c30c345149be64641e5c71fc231;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb824bd573fd92bc56f30fd7b22dd52a9d104d6cbd10252fcd6092212911e85da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f9c2a8f1ab3d7d150b2de37da5ff042fbe937d0dd4450fe8fbe3175e14ee42f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h27dc2fa6923d00ad392ccc65359e3cb1ac3a748c798d57158a93a25e1f3e5501;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda16635801960d27886bc6c0a0399f7677bc272ff04289a6e82fb9ecdbc00bdf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h29ae68e8f413c85bef2b9cb7dee96ef53d26b6589c487a886c91a8d6381c10a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he496a0c27c615462c08a3f26d64d9cdf0f47aeef3fe011f473f83427ea0b61fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24f4fc48271ec74eb595a51afe5e7a3551f5a80ec6f903d1b34ce3301761b6b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c6cb29f9acdeba22f45f523787cf730171cea7f5311a76dba583c7a62040b4a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71a396a77a5036222e705676a9117142f1672a520fc8efd744294073f0da0919;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe8e0c241d46895556bf40fe899c701c8548eae7f81fffe51314e1dc465fc987;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f3ef15286b0e5522e5d2d30460f72c8132a5b0c83a0e3aebedb66fdb35c9698;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ff2f400d4ec0eb4846524e0fd73a7fc9c2d9b966f7d63ae4448b102c1ee82ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99437616e0fa8884f37da424fb2c19273299d8bff8629b988e58882bdd9762ed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha66620eaf9fdee467a1463313856a27899939946c47733fa7a44cc4ed55d6d7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62311edbee4d63eca6e4e7efb2bf491e755a7a45784e3c9c734acb705776de81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc56cb297fba36b0d6e05e464f30ac7c2bc58b6c32ad0e195eca7e06dc0ce784c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b30d3b3981d0a801e430077061fea5c9fc3f81f6a6e4a7a85760747f03b244b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b5cc08f2067c02518eb9106b274e6c20ee7f4970d0320387bcf5a3df6520beb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfabab2b3b55eac1d251b7494b969b10c0929b6fbc9e143323af3cd20e517f71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e1933319558a1f6e83ca131092f32388b460656fbbc364c6f5c2bf39b58387f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffc3c13abe3841c6e88f844e32b6c2660076d32dc7777b76a8ccbf5337790fb1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8897dc3fad577d0e51411b28e02133dbebe956ef9231fce84030e4da47d34fab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc7409a339d08302c67631ed9fb9bd0cf525e206d66dcabfc2f063a8d6947066;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h812f7aa1db33c741e390e2e34c0a4ed6980436e1cb1a94e021e2f621b00b3b43;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78616b89fb2c193034dde675116385bb2d9428b0df4dc47c6cace5381c4ee32;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfaf6649470622f08f5f7734a658e41edb937fc84d85b99f09b60d8a9df9b2d68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b922134fc2883effa4b245dfa00dac98b2c25c6055852ee923ef4ad012dde82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h592c4d1cb98319a83c716cdba7bab50bcc931e2184bef4265bf123caff1aa5c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8eaf6316e7525206f8aa8c99ce3d50c423613c99a2b13f77824ee6b2426d7a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc92e973d89495e17cf3bde977578aca6b3f3662944abacea333a516641f22ce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0b902ae6f4fd913a183ec9914a6e999f23e727abac6c1d371f753458a63b5d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbff0afe9b48ab69a684f2a8d73e37000921b3185728c31749bfb9ac2d90c426a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6da60b780e6735a4eaba05c0d58a68cc204fa6cb67c081e812208a1e1f38ba7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc519b0272cb9ad962240e8a73a720e229a8bb813f0aa3d705f1eeaf06ea4f74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h76caabc44cbc0669ed6a2017733ebf60b0be2ac1f640ef08534c1c89f4a62ad2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he916b43081c20c782dab0b8aa6bf9cc60f2629ceb75b2b0b05eab8d3e270acb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83560d94a446afb108a2871b8443f673d918ee71ab36b0ce76d8a4645c6158d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9ae4ceb6f49d9721b0a13217e318873a2a05ef190516c1a382057398b7fe965;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d464221493385ecea3ee1d21d515a26fbb651a4f7b1cc7006cf7757c05d1adf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9fa95a4888c8068b2c70cce1108457c1fafbad7d524f4697e0116b2af85dc4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h951722d6a0de2b7f206d6b3179fcff8a2b74267656fce234f5fb31dcf0882b4d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89ccc0d27cdbdc53537d30e97aa894661500b86fc087b723fe3f89747e6c26f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h817b8b7858d202d7b4390a8660e1f5c80a8c297b9dffaa8581a0ad25418cdcff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2e5c7eb8c8811c5e15aa921fc9813cb30fcfaeddffd7f2a6df81dde97b073fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff3f88838bb44ab0f79a54db4265a28b971c821a7806a335d71e0456eff8c054;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45118eddc51440f53a3feee9f6277949deaa33c09ea981ecf9c0307dcfd703c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41c9c615d43d02d556b9c12ad2a81f04e723d9f92b823b05e5fe5fb27eb32dac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed65dcc1993773c319834293b7d742dea9a82e6b50cddbcbaef808db6d0ef759;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c6df5a27e48bcb4398d892400b6cb551ae21490a1e02922ef0c8287ac3e965d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb32529ce1b2adfd1c4e9d8f86e4334b131bcaa0c50e9b4eb232609725559669;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2741fc8f3e3b4621412cdc26a8021e6874bafe66716f59656a053f2372e00854;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h48fc7f2bab9b47f8483a6c7cd769713b12c8c6cb177ac514bd7e453f6a68d3d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b2d05b32fac60d4327a54e9737703640b4a7dfc531d56b5dfa391b779efe2a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha216f3e0ee812e6cc8b100ce5ce6bbdfeac7a144411504a4444a42573cc81f5d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11dc4b449c1e07d69ee0f4ccffa4dcc24936a47cfb2dcb50ccee8bdb07df256d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd4cdeb73cc034dba69fc3572c24cd45baeb5f939a54c60d337bf95896b12fbc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac84d60d0ce281c31ba7616358447fb885244bbddb4ce1ca7d5535d952f730eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5470f181ead6663b17f3d784ccffdf67cb8a8b7098089535daf2506b42ef79b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha04a4be6bf893478193d4f83b88964962d793ce607bc88e149ece8aabddd1433;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ff95f3f2090dbc987ba920ba921c9d2a3274655fccc256a75b8f80278f3aca1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c0e0f3e33a42b9da0a4b77301574b2bd4515cb299ec0a63b3513a6122fb2d86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2dbe9e2e3d1eea2908b3f77172148ba4259c5742b83530d6c94721fd6c83db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffe6a9dd4fe076cf8c417b67ffc5d10c404b1b3bd10c91fcd5a1d9e975172834;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6cdb84ebfef5907359b628d745918d4a589d476123db1dffd247f8de39cba020;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha267aab68c66b7957d3e53abfa648f097de213885fd78c801251eaca79c91e2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h76e0de0584a13afc4582ec1120c45e99e8248377627916ccc44c2133bbcc378e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf7bfcd7bb597638e4647012f4d3374a01ecc4eff5ea06726244d3b005310912;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a6a28d4ec430e744df188038e8b7650013305fd747cb2207848b9d332fdeec6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbdc33ae463c7d06fde1a796fc2d7d8ad007369056e1d736c1a9bf53afe8a2fd7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5411982bd1e979f2049ee1b0c0b25f57447720a8d39eb92be2cd943185c60b8b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h656cfdccbe4f9088eec357632a21853d8b12e01e8ff67867dcd0f009b0545b54;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb0fb6384fafbb4f71a7270b42b3bd76af01da3aab504dbfa21ef18f464788185;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb2ccfc3223b20c23802e62fb1f0385bb0d5bfa04332a9c2f726c4f655bd641c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heceb9c73711a4bcb9d4d2f44ec5a713b26b2248c9618af8bfab638185fefd505;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he68faf669933aa12c3fd95dc4d354ff6f7cdf06a934fd2af30c8b4d80936f22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a8f9797c294eb4939ae237d151df009f28e010b7d07054a659bdf537f4d1b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37c1befc2eccdf9b732261dd2646d557686e613e6cfc6843bef85305409db95b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c2eebf0157e1e2b5d1ab4121b5581a23b260aca4bf274011c6b118ba1380c03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc38b498e88bab891c9f7167311c97c0abb1441aa32911f0ed956a975461090d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60519b63e78cc01e8ed0a91f86d4426feacc402180aeb1ebae8aff9d04d18eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h927430f3ea6765da246de17528549e64d386e31bbc2098ed8b68b5e4558516af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h423bdb38ea46e031e3ed46420eb517e67276702a0f69aeace3e88d3da5147a79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4b03645c2a3b9cee887f172a0d9e943fe594535082d85009db1698a43858215;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h543fe5a05406c6117cccc618220dec801c872560eda83fb7c71b334730091776;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1626855b34adeb21df8aeaab4c27cc6fdfac2f600d56779dd82a4dc1c13067eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a9c42051eab9b1b3311508d0ae0462e124a38cd7877f23509dfad65d510ebc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf4c95da584851c0d683aca79b247a922f2c925a9d171048f86ed57eee10fa31;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c3a9afd8890ee30bd90d5e4caabdc496a63443e51fc31ef9306f8f7e7403ba0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae2fb22cc0d8d95616cde3cdd32d533d52b4afd687bdcedc27945b0c78955de2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37776a3bc54875b954506700b920f50ccad81781ca59fcf784f6c0f07ba0de6e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6365c015d01f09543f4660f4355d7eacf9a9f8e1779b413bd0e151787229f484;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h520129ee14f883bdff2099725ef27855ea8c06ed1465549d423b81d80ed4b1a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd918fd2e587d64244b83cef271475700f622ab45864185ddecd2390e14e24902;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1655eeb38718029fa0426afa52cb72ab18aabb2e8d61442a03e0a31197d50c9c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf79b1ba7e03b9c8506e312a489568987de1fc3cd2377c221ba3b5405e927870f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfeea6b8c92e29885741e4aff1c3e8876c4d31c8b963f8963c858786a3172b39e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4f1c030430b4bfcdb6c6291e876b09de8cb8a74596de1f03d9cab4f7ad95b6b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb410a71fccb1fff0d3f86b28927d8b21d17b7cc690bc889eccc8f8729ed7b0b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9b7dd75db86751adb2b54b70c2e90eead61120c0de8871afa180f40088c7011;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heaf497a7ef9a3ff5fd445b933ad9ccc114d0f64214e1604370b2aa40cf120963;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9ef113622e18dcf202fa5671e52db8a8a37fb315e97c747e092a341a2a95022;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef1c457c6bcf0e7106f817d70ac33af9e3973401ebc83d28d0e300d317e3a59e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h264d28ceb62d661ec7d610c4761b95cd44a8b1945d12ef94154cef480c646ab3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5cb62b534ab6c814c4a3e2d5f3518675c7777b0690f9fec9e56629440e1f131;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3eda3cecddcf75e442afd30f90e11446fbeffa07cbe32805a17b95d904bb26bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb349d8c34e9d770ab780bedd9df454518332e1225b671af811973a1ee491d3f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe58f1b2ffc28281104c0eb699a2716a914c57556283db3cdb50dbb2c8290c02;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7576f62bc6084e57ddf7dcc9903e5854bdc88ebe0057b76c53fed90fc262519;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6bc9e62a0a6454aa5464b25dd5729ce46b695196f0cafdf32ad33c3070447e33;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h846f8d4d91c64cdf1af5aaf21ee007df5bb9b7d6e9db0d66cd98564f8ad754ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h907a0a0bff90a11fb81dc593dfcca4812164f23a080f552ee195626cc8005530;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f1d6794b86ab635e308d75e7fd7e779c1de359a6132ff7a64eda6fa6affb0c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2d41e36774516b2aca83fb6b4c21bcfeb5fb2ad4d2f45c919712d9c8921f892;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54b92afb526cffaa048b78500d19f1f2633c4ab84c851898785c6e99d6dbec73;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b9546f59513eff9a442008c24d8383c09c9be88c5b4739d46f57986cc15b3f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h171c845c02fbe8f13b5af78e6b2a7e5de1d31ed3b2789ad5122c06200ddb9333;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h233be813a63e90b54f215b68ca62236edd32b8b687d4ab00093e2c088521c419;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82d00e3676ae4e10ae48ebb1b3f760d0c77ade94916355b15e48b6c8b6f299bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h27857bca2d0ddc1f33371f2d7016d8fcfde35f5df5acfe6d36ca03fcc61ab1d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff1e198091509de6803e57addbc4d83b6752e505a025d51fdc39f420e0882df9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h746832bea135632e8ba48cf309d09e127030b6469be3a29029896bab2070682d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71dc11ef834662867d4bb655bfd183c0d18507e023ccc40c8417792f373a4544;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d5cefd798c6a4bf6dc1553a167f262ac9304c8ba911673b34c4201598f91250;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdfd31b2b413f898394ed8df27f27b06f1c2c0666edbc7983825792598f0dbf07;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d3becaba4294ee893724bb20c5a3dfa68feda45c785117cd7b19dff0ec1359b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h571a8c93842d0e64cc95363f5e8cafb7fa50b624ab7aedcf8a531cce7a5bd87e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6295349f87520496f1fa634b39381ef8e75dc846991e73d77dbd4195e898caf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62fe63a6effeba888226b606f7cb4fc0210e75c65aa202587c8211ca387d77bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99730948ece6652bbbd3d946349bfb4be40fc0b13b6f357b905b6a65e5da5e7d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hded75795686942fa8a8cef824679a03de941f0053317a3bb04f4da7b4667f54f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf5098b0f33cc0fe694f0470e04078b94c8b041d8f34a223ac7b90ed1eab33ce8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha22bf16eaf1d93ca788d1bcca7c0552eb130e5dade1dd9ea2d174d58a0fe8108;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c92925e02c33dff233d4b680015875b582926a4c49f17b9424d8d3c51269ef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb008d7eeb2fdfc7f32b4836cde282f0c8d79b51ee6afa2dc333acaf6535bcd9b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h372ec16263ac36d520e4b6eba8875705bfc5c892590d089c3c67a544a6cfc42e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1d3e5806ba50da8193ba08d5444a1cb0fbf5991538c117cefdc81e5e99f8a79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd47dbd1f87dad23c5112d1f4535e4d4b791207ecbfa6505855adb349e31206b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5df0207d26b12f688b50c17620abbc758352ce18f25bf862763c316601d5f9f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c511285038455828a62633c5b9933c3ca4bae7393b78e82ab177d94748b26d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d9884577772d0bad3d7095a9e3f1d4f5d8be8c9c936e9399a5c53f694c0f37a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6ea4c786b7b562fbdc60f57047d8e66770ca71df99c7193dc209ff132d23e34;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63348a4d70f45f44da166e81a24a77c4ea51b842fb8b95f269dfbb0e342171b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c0d5f414bc1dc41e12bf367721b25cd8f6a9c597093e338263661c6aae209c6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4573888a9a6dd3ba3ccc277e85f45d5126bb6a14106103c53cde94b297cbc03f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc382b1ce94f7e225c02918967129c861ed210bc864310a77c45b63cb89ef39;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6564a82139dd9f8455089bd1e72e9a54ee0110f506f5aa34d8380319073d4e03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h127bd68f21d62159d76524f20a340e16131e1b8940a5c739d5afd093e02e879f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c30ec19fe3097a8bfb8f1a09177b61864e5f1e7535911dacfdc4a45ded67930;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1549fa2f2641d50695d73c452d80f4f7829a8c0c1ab5d759f1bf54496ec9938c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c95ca773d390331ec79f38ce3ca64fd5cef394170521041e452c345fe59d19c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h690807875a9c85f79401bba2b90a4eee73f20d219fdb56ad220c4ef45e5d0296;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha83087b4586fb17141a17aeeffd689848e46d5f237020698ba8bc2cc81b62f3d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2821cda0fd24d67f37c22ae614de80cb0d414698d81639a214409436310acea2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4ca386474639372a148533e106757387c6fae25a424a62bed9e7a6130908894;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf993605b3633c739235792d5397bbd31980369b3dc069ea3574b746e9fea1972;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1f7b7aabc062870afd6b194d21837f5cb4f9973eae1d7e54879fe8344c64dc6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4a08b5850468ae987d272ac5a967bf4e8a1d4ad00a983dc46f00ee6ade65798;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd58489c910c637a06f62c63db318744c8c97f5f1ecf3cc6574d68948c60a44a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94a378054bf520d6ffcacf347e9b796712e53d7dfeed35f54756ba63b20d41a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98a3fb3c2cc84af6da0236951ad51a7e36058dc1b15c5b0bd844b966ed0fb0e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha337661d22f02bd9cd266a295e98abcc620a1a6e0ae4de416a369d2f7c4763c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf63c2f9e984c5fa2d0b491a54d649cdf51e889776a6063014a4796d1e2ea4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb63ce4d870bb25133e6b4d0a23cccdac6a287160465a7cd0b04ee5257713af7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5437bea96af1b710eeced8cb8ff8d6a7cf0eb5f57c6ccd55fa5fb597db0c81b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d451165a46c6c4cf9f1a000194d8bf43f7a5fca5a43fb136882c7866f55d2f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h508fba548f2c03be360287ee30c7ebb42189410951405f46c390369eb34ce66d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31303d4cc47f7666eddb0644f1420940a270f19f46b7df72a8f3f821079c255d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77593fed1d997378e3bd445b47bc90f314db5c6b282b3f6e67ac593150ac8df8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83f20cd97a9b37c81b29d7ecb8d8b5a679498916a621d8a86713aa3ab2904c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdeb2a31da1fb6e558a5f8c146c1aa92da478f9a030309710cbee3e63a1e1e39b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3d3b75c2ee7e73fa7de625d68664a611a192203e724038d62565e175d84e539;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28f192fd1b8321e83aa2cde3d558525c025550d1ef12b146460dd9e9111ef129;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ecb99c6234b846ec772bcbdac5d15731cfab7a31ad2ed6b344389a0ea7a12f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c90c0a07a429edcbe3ecb1bbaaeff267ffa4b18659e45b4452c6ab1ed342458;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc076c1e6dd7efd91280d6a8d8e4d69b0599cf0556345238e95d41504dc1e73d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haec61fded05d6c2e358ee909d8d70188d471fcece08321bbef6c0bf6a7f8d2aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64c53355edaf4a413ab3c110ca2b451a8036ad37c84ef42084f66d0e4506221;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f111909d4fdf429cca5a0066e145cced19e003037eb9727d8246ca3489a0058;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3ae7beaf69af9d12f77be5b8847bfa29a0f74327c7f801137613d98e024e1ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58c2b7f9938b36d450238ded3f4d5ffe0b2245dba1a9dedd847743da16eb4066;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b021a83e3489ef6f66705ddda4038083338aa540d541e501c3f893aa0dbe27a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4dcab8ff743b3eb51029adc4bdaca9298385322fb8c1b8d4709f46820b34d68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c34b4f2808da79fc4c29edb3642985cd09a2911d70cfd515fb282a7b1ba292d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9c025524c1f81338b2156f1a0b5c71528307b9a4864298892b8d60aa84a78f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5412c54a1fc50f55ac58f2cae96d58552ddf77e66fa470f0dea2008f8eb7719f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64207c3d827a35bab1145ecce2261e84a0bc626a764192f1442dc2e85c302c12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc31d1ae46d84b510f7c39ee35c743ad9b9ae083e8d7ab69810dcddc139582003;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1c6db0a9f16c30ff0e56d1666f587c7fea7cbffc031d3e135159c4b7c481bbd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf6a9b4464090f9723eea6a8a984b84642c68465fb38737abc8ce0c710619970;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a08ca3c48fb24cf70d3517aede5483fef3e64890378a35a81b15f7f787e3e24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e7b2ad098aadc802f5644b95d3b02f3b472bc250072d9a094a942f49c7a7feb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he11c640aa1115eed10460494366327a30d510694969bc5826ac82f02e7495320;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d317db4a0457e160c6ec6ab4127aca1bad1bfcf02d551b066ae6bbd187bdeda;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdab92311b58018e36da5214151bfddc64b42d19e18b8ec309a22212aa51fa155;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1942258133d585942db6bd8bfab1a27e0229a469a23d14ba37e0938ac159112f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0c10130a4803be5ccf65765e13fa7cadf490e3854a276c47743d8f64dba1687;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ff7ca5a70cc5c5894c208154f465af62d0a6a0fe62667d5709e9244d206b58;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h791c39d85e683b89c33600c9361c346c4b650eb3c3553958d5313af13383f32f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfcf9c23214981a3440501b780001b4338bf8b77267c559cff3a9dd9a53dbd0a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c5732164bb0934ddeef8c7b63a90b7c45b52c09e85606103d2709e27d7ece86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf34d9bc65bf2f0c76c3d67a91512c527d9e500b03aab19a78e99982136baa57;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1d014922d0b7533fbd8a2c8c5550b9a1975653962521c0d30cedd85a952899;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a14aeceb6c41d056822817302df2024b276bf5361b1c80eb9e0091398a62449;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52d7b6992605ea4e8a66fc15afd2ec4abcd0bb44afcbc1bcf206f824b9713ba3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24dac03b7e4e1693a77f14a05f794755916c0f63f79992575093cb4d0d0ab854;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h470b41fdf29dd11c75226e7879b581d469f2d2bc3cd8934a3feb4c70dcad0883;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd15ef1108565c20012c39e7e4820783b1fcbf9fa94cdcb9a36da90d5f9c1e955;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h14e2d560e4f13feb1f27d248a068c4434d00dc5b1105c0e553c1c912276c5a7c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf705711f01258f9277e8aacc5ab646612e536796a03906239d155f2952ae45e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4feb940dc99e3941b897228fad8e061346743ca7e6a3f2d3590a7044d9cf83eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a2a66d6f1cb20f6744fe065fb68133942cbdef1942e9f5d1f839bb0f9c147bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2215f94b3a862de55fd7c98a1f81cac69447332ca86500d30ca222c52165fb23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1bb8f462fe9a12743a5e13ad1386fcc8defa7d62f7b39785c26f796c67db25d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6bb0584d53ce7c246609a85769b298b2f8ddab721c5255ce490e8261d68f5715;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9b4eb31a752f0a8099f703fea435f78f31ba541399bd7dfcc2d9369b9e564ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h258302d3cb99f33a3aab5c89449b9e8ebf4d00dab80af0a31e66a5cb7329cfaf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5af0dbf198bd8da1eb9f946546719857d7c5d050ea29470136de9e16690aca0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93e3d0db09453c482cb1ef2cec254cac24d7f442982b66364b950586c4e6c2b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58fed94f9f5a5e9d22644b37f281ff817d0471d81da20cf1bbf29dc950af17e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae23eb85edf673c30e2d94b96a7f8028a415e8198940325148a4700140395821;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1290e767920d73fed0bbae98568d82783dbe231b8bd637f5d9fd71f53a1bf0d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc78cdaabf83b5ec0e72a149cf6940beb08e6fc184da28f8afaa47d3248ae130;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7552556b4bfe8db7251e34277e4a9ea7153d5d2d0eed8d54fb7a2ef3ff49f995;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1187af0d98440aab328882e24dfc9ac391258dd81b8559e6f88b76d67fee072;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ee276fea5288cd2a62c5328c77e9c1bfba36bc341d84c0d5fb4807eaac1b717;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98d041a9fa67d4db77023a87ef151b315140aabe4a264ace8bc0fc52ce05bbb5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2658ca320482be1a0c8d121983b46c7623825f2de80e9bffe803bfd1ade17dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a1d759ef377c22c6377c1620fc82af945e7442edce7d92ba93aaa56c2cf4437;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b28183fc86c7b540fe88f7549597a6a7a871177a0ad054a1464372e892ef568;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd77c5e23bdaaa6d2cb654613619ed62bd9481a203f3c7f0c903605d2917001f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3216f38ea03995f86ff32b2c0918f922b4acf13f695c91be8bea91091331424b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h312c7d7e57c50865b7ee5159b9536eb6f4cb5341db33399ccdb4b4d19f2963bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf431efdbd6fe8d4be41dfcbe6e024da9287c314c8f6dbcca5a8c37917d6559e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc49a9378248c262f99914ff8c782deeed88d77a107d86398d75f9a4ee1d2d9b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41b652911cda0ab68aead958857a319318130d135553686bbb047c42c3e8b7a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h931e1fc00bbff8cc85425d32498df3f1f38104402a13e0aeb902cc346cdab329;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6987c0fb8f66318140759796aeaf3a134695f9f33925261fc6d4eae29061253a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h43431d3d4353400ed73503a6da5d081e3534d75801cff1f4c867ca24e0b949dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4232463f70f66ae6101cd80997b91123aeeaf3a54510d8f701b768ca82b864b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce76125fa17501318ebb8374f96295dc41a5e49d39c27fa2525f9e1f9d3a9d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7d3fab62d80ff51c6fa92de0c6153b6ba6f1a4da6015121fdff8619af3892ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h857f9af5837b2f90b77be7774fa63ba1f92e2f9e8220707d1abf1339ea7c69a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41cc64995c6f3d1595966f04bcabf7c84d253fefb0653b93e53539091a1e4926;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h780f89714295fef5727c804a1b073059cf148ebb73e5c58aedb660bfb352a46d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h314e8c93e904a1524a82fe09d2089089ae330b7a6d2d756967e8583f9e8e3087;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4341da779b5487eac895710fb5bfd2e3eba79a11d18ecd0ce91620ee12cee71f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2511fa1b1820eb12a2b47db07a7c721b2203ab780c0a5298e695838d981ab376;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h892f41846c8612e413100d15a991a921ab9ed34a22269ce6882d37cf3f1991e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ec5f1162a1bd37a5b92ddbc86f3ee2b9092d63209541bbcadedb8c4a0d34eb4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54637c50ef3cc4d4189667814ff283edf6321b3379c4a6bdcbde04e846072f26;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf611befe0c0ba6a9b8b52b0efa091bfdedf0bbea02240a0459417a18e013f1b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h949a5501de474e1dd20bf2c2985c5f77617105740ad6f7ca2fc6bbc2d40ccb78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h13c46fce6668244a6bce46b2efa4b4423641e4a0e937d40fa97929adb34fe3f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2dcda083d18259f55a95c40c0b457f179900d354ba9cc504b1f5ee9e31015408;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e870c1985536cb6380da87bc7b24e2141600289af03d1fe5f0ddde9f3903ddf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8727641e84c4e774d2062ced31460352b66fb7cadb1a6d7bff3e01f425c0fed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42798eaf1d7180c0270d3a9b6328fa66f8f7bb4b17561352b38835c713385f3b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb047aef37bb034c7fae92fb6415aa84115e0c4eb3a7d3ecd2b61a549ccf80c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb81440d00424c503c10fdb0f6c6d6f765fb36a06aba8ba9526b0b8951e372073;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbdd8af3b38456808c970ff97035f335e863344e84487d848bba67c87f91e7be4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28f0618c67f87d6e4a0497f93f95498759aa6ebb2ed99145ac8f7ae81d28ce82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h207d0523c2fdd5d05f4c07d1fb3203407323a31a70b188d8528e008c72bbd4a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a6dee713aa3b8b5209389bb29773ce9e83482c1282c459334cd4262f2d378b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd3b606e39f682526f0afe1b9167de856980c86cad34f50eb19b0186c087509d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefe295345b9b2fa259ee050798f35b7ed2d201fb85c1ac23d37222fed1da4b04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h118518b98a2baf9c7cf4eb4e74c3cd1e6eea1deaf0d1ad99f4d440532c927d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h583fdad45133830097da365a67547982ae504fe9d367c6f7a005ebd315aced40;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75b68d4e01e9ca33f7523b58a2224b4f34b33dc65def3febe13c2e8733e2891;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf98f3c2e8a07058fd25d80ddf2c384d645b56173f6bd2403e9061836e37a77b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hedbbfe6f31aef23c9934d8259dac3aa83df9e2e2b99f8fc1df623c740265d0a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca03d9faf44a4f9b22c9d986b1e3cdcdb79213b06d13fa61f5cc22ce2ef5ac5f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a8d6c9428eb4ea9585d9e1b2775b061d1d048ab25c97fcfda604bb11884fa2f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h190cc68648c1f82b659571892b6fed3af3cfb943898eabf498fa166e17468074;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hddab28d9e18af572d48f95476d8229f93487b7f2235322e1555915a005b66931;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52ba47ec16462013e44ecbc1aa797f76a91cee7adc70e9713b06d56e83fdd7cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa62ee2f9280ea2f016ef647a70e8e3094566977a512f5299e54d1eb1d52b7b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5d084bcce215e7583b66f6426b0bbafea06fb95aed72212d3fa9774a04bd085;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15bce80ad1ae0c6f946aa3a587871da559e3d9a9cb6e4c0c97c0e811c49d350;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8bc54d801ad40d51493292a9218780e7bd33361dee16eb3ab30300ef1e7801b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d5140e60cbed7e71f4939bd91771e93f6b6ff974d7cb86f7f045d5d884bd56c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4680a025250869ee5d6e09331915614dcbf8d13fe906d942706dddc1b39e7fdf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88445553e58255598931fb344cddbc8e6426ad0c2e1177c6025faba7d514ce9d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h34b9756ff9c1f00a0cb4b1d9b53bcac3b094a7437683da1cd59e04da52b0ea97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf45bb2d527fe65112eaead8f6f7c7a26efd0a02ba85f2c6ccabe7d0c18a7b66d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ef05f69b785a9fff351e25fca6e750072742d8b4d85a75d4f63dfd5145d6745;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h393b70079d341eed8fe8f958d9165007003ce56f468aa54bf5827d1f433185ce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23b00a4c1ff69664741676bd8aa2a9a845fc395c97bb957dff501572806478b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h844ca5b398b74e725c186e8a3029374557b5be172398ab6b033103735ff045b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc348869474536a5b9eb268ad858c7435ff2e3760d498c212b3042e38b3c90a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h27000e66c59fd2d725c94828bf967e009067096096687801877eb88d2c6887f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58c5920d069f836935a59715d51a6f8c9f0531690c7e0b17a40b2aec579429ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb1593b76def44adeba6a1fb9f66e25d2efebd02341709e01469be09d4720222;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h249aa1b178ea32f5ef1549b5cc2fefff40ac5a8e5065d4f7e030cea7845fd948;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h905ea0c622abe3eac5145191ef6a6092149c042d0bcf96d98e0811646cee9b1a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h500e3d0c6baa1619983e11a2d8d319e92494ce60eefbc03153dd938cb56c247c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hccb139182c6646571aea1fdbacab0bb8b8dd8cc6414df727a98f1bbac51adf3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a1210d51149297c56b90f43d8feb831078bb5980566516d5d4fc6b75227416b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2a88d45df08e864e163300d7049a35e15e8c992e91a2b2029fdfe6e782c526b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba08c2ea4fa85831dadd6e92537b2cb1b495aef0e7bf2c4030a289ea970d0b73;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78ada9cbbdacd6454b2369cced9d44c83a158007851b9c3acb374bfdbd06127f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5da804367472aedaeee0b79eaeb5b0efc3ce87fbdaf63e6ed7d36e05589dba0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a17379d6315174c7c3a9f4958aa2ac14084245cf9cf92d7bd1e837499b6f8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hada12b135913efff445e378bd78f7ef91c9540a58c43d61fbb99e1afa1583e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he26a54fdc69a252c7b12aa3f655a73be25c451aba91534165591212a830f8317;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86255467068a2819dc3d45ce32a09046cbf1bd2d72b4ac2be29e008a9fb47b3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e77a9bb08e02d93bc24b3498b6f92d9da47b4beb1ec57ff2b3d689272c9fee4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7d2e48dfaba961bf46c62e8e344f370d32ac071c7ccd4efa949985659b463e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c4b13a81c42011111b2e773d98392844807ba36e24976daebfac1ae3b688d84;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdfdb00005e7985ae914707c88a5baa13a907b39378d2b56a826d99256ecdc1fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94128ecaa86fb9e4aeabde86bc871369248ca4be389ae12f659e76e5a89b9e91;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha813033320863d6958be98126fcf8aae29bba9337aa5309fb964ba99a10e6625;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0c16308686e4636e2f5a4af941b1c8181d8f4403937ad934ade08e94cffecce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92297867bfa02b9468a40553ee2f6dfb22ee4ac96a88c7a04ac3f40c7f08e5a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d5bdb18ef4677568d7eee2d6269b3fc21eeeeff73cdc59cb96068da379b6d5a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8556f3e12da8d38e3dcb236e2eb8458300dfab9b537818e42213941693c58d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5bc43188c6e7cabb1bfc7937c839ce1bbd28be6fac23d7abf9284e076db90cca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5171a0f8a0dd1825b55c417e1d1ba22b85c986c6c24c11462d3a76aeb25f87ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ce6afb25cf1d236996ffd778183ffc9f00cc4e62131e1eb93d1ef5b1fcc0f4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h458ed801a1bfaccb5f26f70260191656b49138b9d18d7f94332e2410c7dee84e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12b66be974eb0605fd72a7a042372e78e40d5343b987bc6bafaa1f58aa7b742e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ad0e8dc7beca7faa92af46037f447b17e91c9ca297653ed8aeac81b50feb0d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha1126a8b7fe83f0d085c5125a972c44c0ef7e93684ef609fe6cad6c1b8492511;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6a9e9b149a4f6ec7330c53397a9eb412e1e554d2fe52fd450f273335bd5d950f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e3d439b5617fab77e7e4b59cee90544d8de2a2053c4bce04f06fb0557044039;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h144bcb965ed5ec9c102c1796b691327d5d44b272188541cad5874b3f1327ae9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d7b432708d3bfb60c19f568f6d367f3bbba8aea29d5d5240df795949cdee48f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3597155441d8cc9c3c19a7af6fc8bc8225b9f1eab13ab40010638918bcf6937;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h58cfbf626a663f594d877ed86981923c66b281662d008085da6ab228292bae86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ecdfd973af61c2dae4c6a640c022015ae0e7efc312d2cb9e128c977f1a7539e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h845cef4b8c70a308944618203343e6135c2382460e4acc15728fce1ac879db35;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac964855e68b7be0306754c1c5256284044fadccf4f43f4c9dea9c643c88db10;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4b8bd7dba2a47fdb44641b3e686d04ba60e66eec049d39ec100b720a0ca35;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8de0d8b54a5b10e5372ec29606ca9a5a86002130be4af0ce40d836c8f84341ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haebb8a9d4da433a36c8eae93a5495278c7c27cbf4fd1662a418d388dff52ad18;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h610202086e590a0450a2569c6405fad80eb58f39d9e7cecaa81f3337942cea8c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h205969cf087e584793ece77fd4541ab7cd089fa797a83794b73aa376be6e046c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4822f36d58974fd7e5e1297758ad71b5954b9bd642b96d593cc6e7877c365820;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4489bf9b9a79f833a562db82aa3c6bb091055d02899875baac52eb904a0e2d92;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8bd3aa793e80c0117dc28840c670aaa1c3cc310cc7ae48c055437c34e52154e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6aec1d85e9649cc9e67ff1e3420d85394a2c4f2d44457148dc73df8c4a630551;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2067b5ac7785a7ad7bf5f27febf3e39a1071de2e340325755a668decbc1b7f1b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c0429cfcbb23c694a4731730461c32d9332d8ba730d0931b029658c5d20043f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h922a060b34cd3fb12c5b842df362a8d5b34496bba65759b53b327d09c9e5c6e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2498048c5ce4ade363643ff0122bfe07357e2538b13b8f061259cf1bdb850e97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8a40df3f3b150bba96bb50af8201b857d9ca3f4d86643c15e1b36ca496a687e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2fbec477c0646ef32e5db34ef0cce340d62e77630617831f0dfc63f58a24928f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc71cd44e35a639cdcf8b72999278206f058a731bbaba369d887b0e4c6f02c0a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc137b779dc514d15b57a56a35d5935482f24ea529a5e28c109171ecf3f0b00b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd927c5d6c30686c7dcce0ee9f002338bf251f88a9bb1b1ad9a0c88070eeb09e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9944f255eaf44bec53727106e89004d84ff76bbc1618fc6516ff57bc13509532;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf0fb656da0a02bf297eaa403903e2f5f45533e1157aee094fe7cb17a9bf0e5e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60d193c9926a51b807282cdfbd5fe22aefd4aba61857a5e21d6410cfe542bb07;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ccfa2077b173cc37fe08dcc801c11780791e21241258f46cbeb6d8f71431cf5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haaa0f68d1affc291fbc7a2e42352198273e9c6e7c451374078eed8dc63973f18;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha669817ed36892e99335b5ca71679f2675e9e7e87169b41aee5b93bba1f51773;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h728e33a3a32f7e4e273540dbebb886e47407e27d988b6c0e3ca8205ba948f817;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5eb5fc09ed9b694679a6e214d93514b62245182c83ac59c1f5f3ca57c5d43a08;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he390e6b5e7b1ff8752bf9909dbe0737c3e58dd8758941a9bf6e2c50a8c726c4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83f793ee42f91aa32af700ad4b89d8a39823a706410da9048e2f0f2d2fb4731f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e720b427b093a139d5c9c4314724041df879745707ef389e84fdc433e70f8e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf0710e1cc0b70610fa05996a9eee2efab5a0332ba9d7814c7bcc5db5497d7f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h380b4caa3336a9d2a729743c1329a13cbf03f15351543db818d5629fe7268554;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6734c27880dee9b0c1ebc2d3df1bd290300e51ec0bfeaeb1f21510d105abd3ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab992e3221fa1bfb4d01ace071edaa9611c783b35cc09e082256b0224bb0d143;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1c1236843a4a7d7812eac7f4a637d72fae2d3f0c7529da28c5fc0dedee11606;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf23dcbcf2680db92628363ebb57a92a1a84c66ddea06b44f332587d28228102d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h358122bd691bb5f184cc06be04715dddacd0e5803d9d2cba240fb78ad84f5d56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h613c420337a41e32b4bdab79c957e1148a5ac7fd7bbcdfa8ae07f02f95a88eb8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9fd7b3ae09e70061ce23ecf8ce4e848198eee986a54dc05f6f17e99d5180bd5a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h455e594321792e8da0a431f1c74c690aa04595ed3727c18d8bf9a5e5df9a4dc0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4351ec6be7fab11deb55b013853d4cda78f882497c0c5c45dbaf30d21bb2b307;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf71619a465445fd303f1f9e6622022444ed16794ba7ffe5203e6d05315e2f883;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96f1d22f3f78f3896fe710a0df62562fcd584926a53a3eb41c9fb2dc873c2468;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7282b186e19684f1c6eccf466caad7c27f41d7150ced7856c520cae2ef44d70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc3f33dad06df90681df907fc8cf48d943f532c00fd67b040f2919eecd931d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b82fcaf04083cfea6d7dbd998a89163ef291f9a356d3bc220973a444d7eeef9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20b1c3f7511399d934eb7bd2090aee9d96d862e50f099c9a59e3e62dfb1254a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ebcf032bbaacb05ff9a2b972f3499c25fcd1e7fef30260ccd6dea9207d15cdb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c11bf0b5dc6e6934791f4814b193a043370b9ebe637d3764cf3e41dc6a75b80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcfd2d60a666545befaf38c28951d09f1c3c585dda174de752c1891637860f4b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h529d266575d7e45855e2c5930bff622aee2e2d5b1095eaac170025bdf45acb49;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97748669c3cbcf90935164d799afd3e55f4dc27b4219f5d60db8718c9f8774;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23df6031e26188eaa166dcc62034c56ef90615e87e64b899ba379e66268b337b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87d30a246fc0dc3f5b2ba911278431517e6aba2cd0fd5e9ad8dcfe35d09fe00d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha333a4ef69e9295e07caf0d49cbe09ca05edf1ab3a4164fe977bda9d8214bc1f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f7eaeb9f8c6e7b8edf2c9fa77d3f8094755ba278808a11cc4659c7430da5b3e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8bff97170b4dd657359ddab862c01f6d8baebde4adb982931302c3a54b3f2da1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9366d9a3cdfa9d1d45036990740fecab3957ae5560e350fdd7ee9680bedcfae0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc57791182ee3ebdc01d268862c3e3278146ebe86275f5ad7a98bd0589a2ada8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb6eca75149a38d7dc8b4e284ba1b0326fb01e300f3a1a24fbf00aaf63de7c95;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82871a0b03a9736de5db98e99c31004469335ab27457e1baaa81a7a0774855ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he163f039ee4b0ca9a0e312f36afa33359c0c351f4c4fe3b2532bcf4a98c310a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h738b8c542d7e0569efd6f7db6378b86228eef0d3d387901238381b31ce5134b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3211dda8e1d247c46142cc76ab67d63fd1d219718aaedc494c07b65e8101543a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef62b4978ea5c9a29cd512e5fd9c2582a02874c13340abb8040e34bb88c5bf24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12a97cd36d23aca957285f48ac288afbd49770b2812d2ea7b502a61b2fdd4c58;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h754ff9d687e59865161505618d43e450e4cb07a0ae88db2c1092004a37ef9a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcdc2daa2d6f3b4b6768827df64d868f73782174885b5a93c0e593be68ff2d5e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha34578c1fbca870f725e1c8b07526c87e618f4aeff0c11069cce0a8a070af467;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d68cca91cc5d543241a2acb8a8ae42d7c18168066b4fb02e6c2957b598fb46c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba5044fffd335c0be3a975b1c96fed7257cd863fca6fdfda557dc2abfd9706bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1448fd836811cb3fafdd146c1a63b9bb7909a23e4b13b1bd9e1afff5f03c5f81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7fe418dbc21c24a433c05279071117331b47c4bf117cd1f390afd3d605d1430;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b0160d33e6cc3bfd1059b991e86e60198e58fb25d1f2fd1d151b878872e3aa8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e8731db269be06ca807421e0ed203846fd181560095a58c7e263af360448e2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf743e52b850c472bccf2f6a031abb1c1ebd007d9a1d497d5837287dcbacae80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba56c7856e84b761a1c79dd0052c56ee121041c716ba48521a782b75904ac213;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab392329cf2042ca75eb6af728eaa10915d35791f919443c36ec5fab17ce2d9b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1541bd88ddaed196ac86eb82ce9be5a692b387d719ecde7ee375d43161d6868;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd739fa7e67b1e1c6c2cc89e13d63259d6a06405fa67990722d6b050ceeb6ab52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10de6be2fe55e0529a2850310302d6eff66940521778134b2ce0b4b97f184db8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a5fe31987d915d1e104cd30ce789bd843a828fda7f6913a6e9ddadb8976caf0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd13367258932601173bda27532c34b124b873cd2be6aa7d5c613e3c471756a21;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb786b77a39a5db0fcfdfd218d3c5c82f892097a2dcb5b6d3f338a1689dc729c4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h409ab7d4127de107097cc4aec357fef8c020a2d1ec638c9af8071dd7d5efaa4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hccd720d53f99742ef00898950635d0381ba442cd814e84d978a205b42a19d432;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17a45fcd76b28169dbd6d4bfef025079900efd165e53a3be838b0a235c4b97a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff84b3a46ab1c1e77a2348421bee0fe52ae675eb3018f0f109c5e7af4ed53552;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb4ff6ff8eac4c8bb3343322c9611c21c72243266716765a9aeea5c28cee3798;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h409c5c11da1804b35fdacbbbcff382eb75aa3b12fde00a2498022d37bd05d667;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42f03c75d802f99710485a1594fff0b041a10c19d177e77fc5967c31c9100a04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h664906580ab3d2e388830f53e251ded190ed5a8615fc6c94859293634c0839bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57352469651ff4bae54def043bd8736d9d773cbeecac3fcfbdbbdd6b696258b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d0fe1906d1288f68dfd5bfe7ab2bd1b31eb9e86cb137fd11c099934d48a89de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb71642bc75a55b2f0de443c0b93c4a923ad023cbd987626826de4988ba9b634e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f1bbcf66786f79f1c30f696c966c195b57b9ff075f7127741ab334e8a093314;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbfb044841b7b420b781d8271c1b10b0a7634993ae48c0076e0ec49a572e51ffb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2be7c6f3caff775bf2d639be448feb289665146d7648e4a22dddeff4ac75233a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab9baa3d3521eaeb674248d34c0de0a1804f842557c6c2bec675d4941da53da4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6081e413773811303ad90d9af50cf8770a208987b6598afa50ad39c7bbdf99ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38921d6dcb47c48ad72e54ca07cc72fbd3dbfc4ed01d63191af63aac6b2483df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1411335dab9af811b699d668014d5fe86c5b3fa4d6b73591f84fc132cf70ea0d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he857bf9c939e199e25ec18add961a2e348c858f4b6b01a7bcc3403db468fb2f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9ec5d83586d51ddd7a112258f7012aa1a9eac1601fc68066744254da17ee293;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e646587c90f72baa235475369fce5b8ce209b787804f7705f71e993a0ae3460;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1e186b712c6a0ea0098cd82741617c34b18a061494f12e07ca996a9c4f16679;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90b0c27ad33b23bfe25e1e4dc4c64449aec61744e7ffff1e68b791d34ea0621;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha1a25dca601f35bf1ca8243b24cd44cf798d3f379f81c55d03c1d26889450ffe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf5aea7a7ec4583487ece6cd2af44dc61634fdde2af1cc1a6bc77041e7d21247a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h713dc89e49307520730cf54fed22e76a93c151e96cb70a351f0bdea76f247a39;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha80d4140113c935e6482d3c0b771c40092e0500ff6361e0ccd1377746cef77fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a501f8a347edc292800448875cbfb4d1075c5fedd8c67ddbe1ca8c89a71f49b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha35af63322f4fbf9d7e03de44fe67433ffb334ba13eb8c8c9b9aa5b71a05880b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h229758ca1035c4a6b7feae75f7a13dc6c1b0722787559f70fde7bfc1a4525b3e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb23761ceb796d64c4da17b04126e0b7b203da13ed1238bee79573b9a7f7b1db6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb0b5b80cff2b8c0686920d2079c2a2bff35971c476476ce8f33b4fda392c6afe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1d9903ebb0b3a17e948ce0ab08302dbdf6d92cfe43f638fd3c003614a15061f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf85bd2b623cd890192c759ffdaef788c68bad99d1ba6cd7a9ad82dd5f2503998;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3691a47f9ee999f0b1cbff01d5ba303135ca1e4b18815604f67898e8078b716;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7682bf4702f6883e0d638ea7e9b6b4d1a6229f859ec98571ab347e8cfb99f41;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1874e2acab99d27e6269ebe7a4922cb896e69291261ea1a25718cf4c0b388c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1fba1cb6037e2872311075f68c79479d8716ef111fcdcfa52ad71526a53703b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb0f9f67a786e74c92a2595eb1f55ba65d263ebdf38aafd715a45ffcd93d6321e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e67cbf6052dc04f2dbb7c0f2c496685aa76f772fc4af57600dd7d5e0fa73db7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hccf44cc2cb6d77c7e85067107b59a1ffd7eb13e87077cdde26a12ec05c6fefef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57338262cf9eb271dc799374b3677ba71b64d29e68e96169e86840c17b8440d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae3685cab1cd55480bb7f01b4395ae91fab3b6e9a54e6cae19cf83949cb6aad8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe1eb4dc72a3610893b247e090376d56f4a5ff32522c2f13041510a563e2c882;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6f46f65324a564aff1daed6b9c1e5e5dc480fcab994d883ca62d96d23b2f307;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97bb58e3adbc0c240154ebfe55e7f32993cdc8c0600d351fced2635b80ce2ed0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5cc0371da5b762950160a3bbd02191c93245bb9a181d5d002c93e271ac274afa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcfbb60505433306d00cb7800502ce8c9fb8c8a484085210f3320c1cffdd12bda;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e145cdf7e099b2c239d6ec9aeda5b8cf2ec530cd10cc1eb3db6891060aa087a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e15df6421a9b352f55718b9d05593d31e6a4a69ad171e4d6025e7399144ccf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdde6979114e08ef7363f8cfba11a4ebb56026021dba8ef2f850c2898bf6b4ae3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h42a4d1406a99c99e3a0f3999c36f0070e59c10a379839b2beadc4effdfdc603f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h764b6d59c41ec168eb004656151e745f721a519d730b9e0b3c9c57bf456518a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4dce0f5e641de7fb131cc4ab1664d826f5e01a47424647266ddafd5405b8842;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h154ac264ba51d035d36d7a944da3828d4a3e1be560b78528794cfcc9d498127c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7143bf573f7819a501c523f5f42cf8df7f0772fe4f8af81b89fc94d4314a4221;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc75aaaa4e479dbd9369f1851c96fac9ed1b28f7e3ba378a7570a0311df0cb0dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h642fb53ab2d9bd944980f5f845c913a59b1a9edba0569304fb5895e5d4320936;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6f287f8954f85faf21c2f422649d70bc790517ca9e58ad36f17128474f7c304;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf382e63f4adb627dac2d467e980c8d4d02eea604f2dd892ab85a185b78ce61ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6cb3ec2dc25fca1b8db8f894f9d54330071ba2aa16c80038385302cfce47eb47;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5cef3f9e41ed122bd3ce563256f3ecda3ba10f5d940a3c32ee9413372d1af276;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4309a134683fab8225a4e1b02435bed0ce497dccb7c08927a24daee6481d6981;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e861704270a601ab5d4102bcd811488e215056840bb67e8e272d694ae8beaef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6513fe06046ebe1fa6a35ea36010b1e9293d5b030f025357face350c327845b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd066f5fe52b5c38338e555135d9b7147c6d1c6c9de3c2918df4bb79302e4d8f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc3ca10a40a2a38c27c3497ae14f434a5b37779df1b129547a4b564e508fdbb6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcccd64f131b7e2f5901f509a51d6e877740971269fee7a80a00e894b25766033;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h95b870557ffb916033939ed62c6b065f8e724a1f339445e0331f65f10529e7cd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c9bf632fb30d303e9d2483b228ef74fc942ec3bbb17a4f172fc646cadebb16d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44feaeb82097a9a90fa7deabefad0aa5cc0eec22ff79e1506582f929dea749b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f6e017653776d72e368bd91b0b2d32b52d12fc5d48f6cf09029bffed2586cf1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8991051abd7c8f3d65a9eec7d983c3670a985837d13202a82704ef8a2354dae0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfbd75056bc1cf2f6a28bfc04c4e021798a29dba86077e76bc1f805ee364d767c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b6dd2c4a542311aa30d3984285b987e6f1b26b01c94541dd9465f640f89fb9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2bca25ff4327dc16baa3c33da3f34545f647aa72475aa8b5914f09bc36d5359b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h137ac99dd286baef2bfb9ea5615661ed61a0070e72c49b814b1f48e522cd2e4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb0f963215e76489d2ec864519a7aafe26a865b872ffdd0928d6a0aee5f61332e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa8103cb1e7f9747e151d9f5c70ee3397bc9c9fdbb9e871717bfcd078f1ea7c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7bd931721531743948a53c8076b3b5336899d8e56b070d64dd0b0f40eba9874a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7bf919bca7585b98caa6c5004065dd293f51a470f4825e75ffcfe89defd4d313;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h367c289b4d4f33b658d35a462f0be0e7d54bfcfa2a2fb2e4b46e509d4f6e12d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd403ecf42d8cfbc8c7b389e11adca26fec8ef321fdfd2b9410c94316fcd2521;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23ca6a18c5142bf446a8500e445032c9f2cc508f30524c05c0b1cad6fae85c17;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7f203db7e4ade8530e39903ce7cefedb8649862855ee7df5fe0defbd523d1a67;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h536c12455d0bafddd9d85fcc2a7148077cde9729fa5dd8c9f66f1f63330d421a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54761700bcdb166452d5953ee69125fb71c659ec7d55f7236df8403637abe6ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5983c19f064736a83da11d6f61e80515e8e1d49e871134b65dab447ca4883e9b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa21b4e88ea21bb0bb608b4e22a193b853f32bb064ebe4e6874af12a507e1693;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd085f7e186aee29e99be14bf77ca1a4e7de4a393b52cb4e756435bdaafdf7c89;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ce5bc7132c56f92c45178c1a980609c1338cba096f420497f8bf806d0da17b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4f81173d091d33e2a9811c8f659a1bf204d4ad67dc03a6c3d492faedc358f52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha17ef6349b374cf16edd022bd4cbde62e92a849406557285859aa8fff5d7b58d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfef0acf37b90cfc2958ceaa5c197639d1755cd83542133b0262ae0863f899025;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b5a019102a7f597b41fe9245e4879730899da862990d31177fc22968d2a9f04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfd20e64d05bb8ec13df2a6b209dd3bb839416632f185c567f2c1cdfcc8696c79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdcff78037e060d7f5e7668aedd74ee680b8ff92ba9884a438240e5cba1e9dbbd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he099a23c68b036f222bb0e63606df84f95d49fb9b1463a7c7f60b7ca7df27b21;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbbfa7662cea99839b772bbfa0a75e6636e45673ac101884b234c613156d3cdbf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb0f9f3e566d8c8e2d24284ff263adcc634d8eab4c176ff3a5ffb432a5b47f15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2a914c06ccbc69ac5edceeffc1359f2b0d9336b586416d45a2a413ab67e06ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e02daa6233c2965413db91369f0c19730f421b0d326e72dc78e9fff7f4f0311;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h191fbf69c79bd1142410c9795f386b2ed0db94e75bbcd15ed24f2d5e9f4f2c7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc8b2a06671f3d91035799fddba7c76c9982b6d63cad0f235c005968f18207ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he96691c31a354562ff7cf935e797e9b259c28e97d3d6aee65d266bc495099807;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4234f4c2ae08744421977133201ae8569e4fe7fff55800a0c1c9e260c8cd38;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7ce1e0facd2595a977c9dc2efbe0cab9bcf15443d7ef145c42bcce97fc11f36;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31bdd298e16086da1e8e3167540975dc248e058d94f86fe286583115cb37ab0a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e5f21c3745d669847eaa4c22544b9167528965a4bee7e5a6868301bf1ff8326;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8623766a42011bd13e31185c7e1502b4810e2ac9c119ccb2bd5cee45f457c70a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h479f73efb253e8dfd25ac970cabe9ade0fd93bc5f83cb4703a7bc12db4cca7c6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb36d4572e11cd9120f76994d7f4cddc94c88a8b18db4349d97cbbc3e98ad3111;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3bda378c52301f7fac7bd5cd54e2081e4657cffd2032bcf9b256534b7feeef56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf00bd60cd1d39c7acdeb199d13eedc8f54d690ae7ecd7dedbf23a2af01993bc6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d7377973fef6e90cd41cc8137d86f2cea8e23993f0f8cbff60039e966c2ef4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf512f9c1b8247556a8798dd4b877d50185db531e3f29508b48ef454517a69864;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac73084ce3eb5a2bfd9037121f91c6d938db8bda22e22e6a87832100abd196a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf96834966dd3f9e3fc86cdc86adc1bd0baef0193e29eb3366f8620081fe9fac2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8dea9697f32c8073d8ba05f509aef4354b48947ebbf6634d36dfa91e12f67c78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb2cb2e160198abf0ff7755f7af923009d86041f1106890137490610fb2611dd4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7af6a9e2c867b9939b9bf829911a1a94226a7bf4cac4261a12fa9c575079d71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce477609c47d93a17011354dbb2340b2bb6b8571fedf8a99e9669131c22e6e9c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9456276ddaacfe484af7835305217bbde7eb8f484405283d7aa604117084d5c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5dcb8211be6ef5ddd5ff16516d7951e475a7daf67ea1452d6ac3efae56c3ce4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5bf8277d01e4e90d7c196e4384d5cf90f91bdab4be7e704414ae9f489fc1fe8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6f82b7c7b98d981defd6f112b1478a91280a599bf41699d3aafa281c43740de9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45760e7d7e39cb382f3fbc6ed0bd5ef1b00b2b9b9c06ba8c6acde199ed97752b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h756e4b3b6498fa44caababbcdd6e17e0e93c328aafbd3328a1c34d7a594f69ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf722f3b0d5f5134f87040b1c15f565bc636b9329fdf7ce46fae4d5f751221ca6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3808870ac810c0240953e2d39d9083711e1aaa1804b4549451ee1f5919c32e59;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd12d8e122d55e2cb618627a6072bda91da7840b911a984b1bb21d323e8bdedd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5648dbfce50f998c18ad43ecb2378fdd2752e7f8520bc48ff46744aead8f8f72;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd61baaf5b9d1f6ff6530a53622b17e0c29869efad0c72e59208259da18a28e58;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0f7631d58c01be9f269470bb87ab1286e3ef2e8e80880226a28ee05a0227af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf876c228dcf84da1c6df2536a5cef860b232746243b99b1f14468415cdbf53a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd591b2f90428ee694fec8aaa7df3469afd3d798e5763fd8c5dea1d10045a2fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb90c6f81789c54ed19dc1df0348a342245e1ec1920e6cab1bed8364c00bc288e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4815a58169b63642ff07b2cad8deec6e09513ab211669293240f8fe37a1c5430;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3fd3b2944f503aa270b50cfd9c71261229a522843052962b94fdec14a337359;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e98cbfbcbd838cf7b9c75e937272991438dcd5779c1329912f8e9ac0569b003;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3edaf92650bcbad3ae2400ca0564f51e4ae8d32cbfc8bbe93e1e6a7459e24bd1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28985bce83a87fbe6d02c1ac4d10e22989ffb016727000aff16e0776b356d917;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdfef4197a22149b46f1285f01b3adfc66a355469af1e6ecb75913c68d0196957;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31afe0fc38360755d775a435156b34c8366c66acdccbbf0631396555cd2e768b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h343d8d4aa91beca090479f82575225dc3bea32e12e1f83aa68b4f8e0b43ea583;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6c42e182f74266bfac2688d887f5661226dad88b03ed9e80cc1a41b77c831d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c29f468512e09dd4a0de0eae7496dcdfce67fc4c547431ab4812c9b5705bb4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h29128c9e07ab2b8939fe84dea8b6a09b01bc985966b3a0a161085e27a383a4d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28598d2fae576e2aa9ac84d8e38609a41bde4a477ca8544edc4edd89592fb28d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb883b8fb7fa58b91baf39fe2b544f443a5c789cb91f9a188e1b8c00211d5c3c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed57c23de8e4b12616a80a1d134e570433e283968e98b27a46cf7ae5c77da894;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbac2b593276c5ce2a52312a464ac31afd9a18ed1abc7a9421a49981141580899;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35b5f73ace8078dd72cbfbe160da6b28a6c1dda800dd61f937c91814f23f9579;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7087238e843e54e9cffeaa03161f7bfd6f352072d424cfdfcf4d82150236a051;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20eda4242d88183cfd8c5cbba6901f39ac909249ffac79c86898badaf006a57c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b531a7dd935df9aaccde15161f31fc79eef0349606a82b02af17a6b80e6324;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62e8aa1e027d639cc80b9fb8c5914ffd2b14657111c2c1fa00582378ec997036;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc288fcaab199cec396f506361178fd53cbb3b0f1501f698c10b780b786dbd4fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h30b57a39679d1385ae68f898ed2194dfb7bd7924ba641dd421bb9bfebbd4758;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e85fd382616f5f6c0afe3b2b6f391fc1f975db64cf9111526f6ecd3d5f75d3b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbbdc8376b587372450a2aeb0a5f9ec55585ae8e61abb7ad5b563443361e6064b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39b94e4198e6f97a3346b89d0a4e2e5b2b5d625acca43c6be60e1c7404ba3d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb580d7bd7e03dd57cdf325671ace17ed174e8eb886a1c73d7e0b76ff952fbfa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hebae8fd64963406469503de3189dbe0c5d65797b0a5bfa9d8ffe5951903f0b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d5d094657c034d93d70f6b5160c04b787c8c1e645fe08fa03f1820d3cd83092;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h355c91310075a2e6fc297807feb54837e5b7bb74b1655575e7316bf9459beeab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19eb5025459b098bc5d2fbf7ff7e0a0a356ffc2d69f238b09162a25f366719d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21faa7acb3216e8c3d4692da33f5a8771baf16a330dfc4c41a5d1f0b24b09142;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcad0e7ca4253f30b8594b757029b5c546b1de67459f8e400e5613dab97e3a151;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc82a0fba83f5f9b4bb588d5fdd375b5a158ea74c6e6a273ad528a05113a14bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45db76f82ece7f7c8567e89e4cac1d4362559bdb2ca7d1f0b242b83de26c3b6f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9aab8b9cf2758c4d37014c5657441b8928ea5b2181b45f9a0bf2ec21e346716f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7d43d9eae4c7118ef01eeb5c6026a95b7f9ce757f9cc76176dd25b86b3e7593;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e3f3d64bf23ecdbc2260b09c1efd959b6d6cef13b6123008b928684de56c2d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h416dda5a90e9f6490c83c93a5289606ebe1fd7b3337a7d86ced35b6d71874345;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha593f6d9fc79abdd50707e3993dab62e5b9c19849ea734f46c5c123489750142;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h857279fb8f13a4dc4601724ebf34b87c23f3b8044d50801c9f1867d0bc313a34;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heaa85c0a7694335f0c1532f452603a5a45834d2fc0a71468c292adaa2da3a55e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3290dcfa790590161a861acad0732eb630f88f8d969100812f68cc1c99c100e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3bf7bea19bb625f968b8402baf5df4e12dccf35e40c6dadc6e22e31ee6add2b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe7fe694c69c067205da27972a6344d253a2a133ae9329b5fbbafdf8fd68f84;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9daca728a44215aea8f7ade23d252c8404de8c0a59a5d6b87e20b24976710e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec36139376c4e6bcb04d867605f43c1792253c4ba25742d69354c2e25fb544dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h27556e1f523283b67b7675031116f60b7f8cc2eac5d9fb95702f590ed324aab4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a5c0c4e8e28a377d74cec4d8e66bd9a443e6ff9fd9e6d6790340d19e4eb13df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4ebed24c25941791ff1577f975d9510e62cc8ee3ffb21cceebd7256c3f931a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb09a1066352801a70b49893ecd68e323c444d1ee9d5ff9b6dd0796c40cdbcec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86acb86263cd1f8bff94547f8fab7ce7158a5234dd4b27250719f8490e3333a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea3d3d0c3b3cc71e6316c35a78638f963a68cb434b01af26d5bf38bae773999;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32a7d32d263450d808a83f685e9a94b7d36f9687f6e706d6d491cb0715fa5c7d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h336d5646ee9ae5acf6c2603bd2809ad72191482ec19bfd2d16505eb1bf714ccf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0a8e5af895445d5307130572170664c8e51bae4110851b36eefee361bb8fe95;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4cdec9fbee629c53b76ad3c385b4c17f3073338bcf6a374927f1d6c06c5f02f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c7a88687a4787fbc1d18e30673b92d2a7aa2d38b703eb7ec4d5be0bfbb538fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf10d7bed5382901666cace86979f6b165d1b980c0bbd8e9cd16b07cfef0f4e12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab9341ded1ac9f6666467e66d7cbe9fd399fd65c4891182ba472bc58ab327fc7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf5e67e87925933d16ec242b3ec893015df81a02aba363e86b9154e923b648851;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9aeee91394c0bdb055fec4fd9c1ebb9ffcd014c38ce009143aefc5f16726dc0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d2bfad4a38e1db55b16f251b317812de9a496dfb3a87881dd56b65a2ed3a2a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4edd756988ad48e160864ad1e368be2a60006445c9c1542a2802299ef56dfafa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he182fbae6f681b7065c4406cb48dbf427b8f3e155b1b514ac32343979d622d63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ca2ba9c16e236b4837d74bd1f197d3f84a1916a57c97c355083957bdb4559a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb40c4a3d8ea04131196353afcd103678d8c26bc31c4f242064d83f8333a4a623;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h620b108315f6421a2122302f92a11367199230c96406ffc6449378a301748443;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d0260f67649d34cd9f92b14086a328afbeb4c566bddcb1a4c6221de3b93c360;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he28697035005f702528e06b65018e2215a83d98ed1b2ccde0ce5dba17781e7b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h844253c1ff21c2c9485b83ea088a0d43b3ee935dea5498481ead297653b03668;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d0a687890770e72c7af4b12ae38037885c66812325c698b453805f7e3044a32;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9fe8d0fae791fc60df56cdaf505736e41d51f61982352c090e30596cf8f1eebe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h79e7044e1bc666ef7dda32a68d801eca231bd7b227f1569605b82a071a2909d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e178819699934553b6eba82384001f94d872e574df210b84c2805f5c9f11bba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75f4ea1fc317bf3108de8c226c12d8ad7377887226028452a96d844dcda3d9b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf6c522b453bcbe2ef893495621ab5452c5ec1fbe50b18a01fa3d73d190d07f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38980afc56f0727ab9029f22d1e26b142fa433bff5156dbfd3d5b976cb6aacb7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he43c1e53177ec5c1a6d8510154a0313ec640f4befd755a46e721effe3888956;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h34209cc14184962677f470d35d0433cf8dc4fa7890d891e1824e18e2dc5de9d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcdad61885cd1937b2da155680095df8a4e9291a4f7bd34813cc08d13a125ad06;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h747d7674c90ebcc5587b1bfe79e1f6d9188d4cab81f31191321c4143547d75d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35bd37da842544ca5b98fc27764bfd242285ecd4857e401e3b7d374481c9f0fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99c64147ba6d4df7b21fb1591a1f07f0c96e20f31d16f03b9b65375016c730e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2f06ae580c996884968fe26cf5042453649228e716dd830b947ce82d56bab02;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc64949233030d74b5396d0a0f85008aacafdb2223ecdb0a615ebbca31d774a78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35bae0289f57104bc7014e83e65914a06f0b1e222f4bafa6bcd2bfa443625d80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b894cd47f64eed2003d82d59b9f367d1dd65f6853fd061068bf7622b287af33;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61b23c59b4ca273da404d26eafb12e9c836d9180e517ddad81d656bcc52fdfb9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83794385b8c24164e09cc9c2e9631f3d4a0b5c938a1a6d0a5b7874b66b5ef927;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb400b91f9374799f6fdbc07d95343591ec893c2608ad9a920bb3f83f4270f174;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54a4902f26fb2b4278a8903f50c33aabafc482313f7de7598308671980b4d31f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9546ebbdc8d46374706d862a093d0fdd65672419bf1ce1ff8eb1b1ef6641d846;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haeb2da13e4cf841778eda896f01d49646cdb9bdbd0e3f8eae211504e8a1adfd7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfe8335974f1f4ef08097c018690786e1ea3b747f1117fbb23884b0899cf7e81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ac15df0bc4f25b85e1acc7055c65e1d84d826aa0f7bef330c18b88208901454;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb647b979a8f22ac6b28a080660afd44aedebd31549df11fe7f8b5c035e25693e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h30755bf7844c5d21fe126a5635b67a9dfa8c852c8e0f8604f97c9f989febfbd9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf87674862ec2c751c7ae95ea91d4411c8449c76fba286d29e53aac79a528581;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h29209fd7438e7bd812695e09c56dda33ade08fd44cc515c685c9c5b97a0e3d56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56ee11cf87f0683aedfeb48063eed50ac08828fd684e29efb486c29f633f0290;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee7bd85a49b01b633fae72b99bf895059219ad30639aa92a85496b52714ae20c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf044d933aab24e4319e696c50f6af416559d184ebf7347771de98dcd922d0ce3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hecdfe22aa83460e3d4f2f65e10e41d884300ad5a4da7987ef23602932a4f717f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1dee861135aeb949f637bdf79c0335fea5578b7c31e41f1412f2be041e14a52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e4d66c8bff572d26dd95e19d13594a8f91d2d0d51fae9a0120185606f314b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20206b3ac1cfba7b844a670c580b88e36752969288a72a971d4fc555c2c8f32b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47297d2a4bfc9a71fdf549a7756d9cdd5f0c10098e24d3f1626cf5a7d0de06bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha873852cfbe86939ec205b55a3ec7d1dde0aaf2458e7ca3758648e28e42ecdfd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6ecbacf20fc450628c81a968f06104661e97e8b1447672be7c2e54b52e07812;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd1e2160a23fb88d128ffdba1ddaa845ddd6149bc0d36b9fde7e801c0108ae50;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h798954aad6a5a67cdb70d8e14797628e44fa4460213946d38d2f5a4d415b80b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc096932276fb20049e419521920231d9e4637dcf22b34f146d31483362220c62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h723d45cc388449e30fa1bb5113758e8ed6826a7844c387c36459c24becf8857a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h825f8e2bb53efdf012264c22fac8f9558f201656a00e593046cfef28149703ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he95f5a78bfe8b815ba4bc2270b43766e9b62ae7557bf4f000181efdb41ff5200;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46c32b45e187f140cee8da960157f5e82e4c1a2ab92a7181a9c33fcaf68c238;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4eeec66f5be4edf1328dd82b4392a2346d3d58aca34fdb4cb73e523b192a365a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd57805b80fe06fb12805a44dda8be11f8267a9713d7aac6fa7376a4cdac1b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d096484d9391d4d2ffde8b0cf156a2be4b6369a9b4674530c68775c61faf212;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha62c3c1b9de5be487641923154f4eddcf79428bba407919d354b2806cc61280b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf869ee2e420c98bea0faaaabfdd8a398eabc7a93b1c210c20811929f2382801e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2cf861a7ca9d94e808efe2476c9079c511ef0a2e069166fb5c2f68b9015ce66;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7fc7a33bebad5bf7b81dcf7ad64278c3819419cb0c6754a68218d0d5db6b181c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdae976bfa34a6c65f73ba6d6f999b43e841c44186163369c03dd844221876d96;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h558d7d7534c248849f1662dc7af73fa3615ce9fd13fc8e84953d059b359e343e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd162cefdcab6215a15dbd76de9d1d52271a45ea862618f5b6d028ebb8793db34;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h632672ab89516d9cfbd32419d662da90dc3991e47fd8d321dba93dfa67bd0dd5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c55d422c4f5821e2fe096f440897736f327969fb9ff3336ed259b978b14fbe5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'habcb61bbaab8c41bf7a5bfbd72ba130ef50dce8b37bc784f1ba08d03fb20cfd8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6cc8e2ea1742baa92bdc9cf40f8fc1ee88f2dcce4617f18a9ac2265979e50e75;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha93fd97b8e6d06c3c3e75980c8608facf7777559efbec6bb370d29877ea3114e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f2ce1d414fa3b0c5e06feec42be78095381ee01a156ca6cb93df2d7f7b93b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4165c41d71c85dda87896cbf2326b2461f428bdaa1b595e905d7d59ee5d187;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hddbb429c2e5400af28043f9d7a328dae49770afba9808ccbcd29c2571e1ab443;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24d6de8fff600df4ffff86518aa6d462cb43bd63dc99f0d0c368b6adbe0949d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ffefa71c98f3ac3493138a1f369e4a5f173aef6a06f14d91674b50d10de7e70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ff0b2807758961351c5e65b20663db34bfe94f02ad41947f3ef89a830c5af26;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32dacdf0fca7bbefa5cc3a03d047b521e1e1efae5755ea29b8bd94c3f04be7aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2349d466888fce13c7cda2f1d367986cd8d3bc68b5f7cedb3603f8066f93d96;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ecfe230ba7701110dc6c97fcfdb3f30e3ad609e9cb9b67a85faa45b96ecd0d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc658e4726f7e77a0fa12ebf043613deb796bcb033e690ad44cf2193c3a431d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17b57a2938418099cd677286627d1a686aac95fff2fe7b459b50733f84a04984;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf29ab5677fdfd532c610044ec554769f76b879f9fbf740965decf7c00397273;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf7b72236cab4fcd7f04d06b1175b0ee05b7cd819b9daed0f1ba3d0c070febd5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a2bb9c72fd09645298c629049eab208f904f479de89ead0db1f3d5751295ac3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9872ea5c45906d3c0d05b1e1bed4080e759017f40cb1234c4176e8cdd81f37d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb107b02c8bb0e8b75e65917e89312570c7f13a4808bfa150f009ba0f7e23eb24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3bc7a5c96e3784923f74c530eb72a230c445b70bd9e5e76e7defa2c59dc43259;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h421d1cfa5f852ef0be07016606b097168385d8f7325acb268dfa5e8fed5dbda9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0938c633c143845695bc7de36b9f825e2ce6823aadab354e37cfb102e28d526;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he50d1481f32e0f5d4eaffbda4204b7f1c16372dfaecfefe518973afe2dbf4a53;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c97ce8116cbcdb06f04bbbbe38552e9b04573ea080c65643bab0ffb84ab14db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5c69565ce1683e8d0d5887e9a6e5d5f5183e84d0eb27b6aa78b607370e106ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19cb096e4f5a95b6c3b2d48a6b4222197b6f7a0d9ac083edf77841d69af3afb1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35a9787843faca7a7733f67d590e0498830d1cf51d297526443244732550a384;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3cdd5cdcd62dced74ed2dca6d5e655c90c214ca3d4e834ed200af692873e36a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h972730d21be77534e649c44de126e9d3a21931b2f0edbadad3a6604601d37500;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ed659aef160919e1c44e96abde7150f26ed7f6d2d84b7b5697654cdf99a5a57;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hada2d4c32461730dcc5f0524032210d859a25d7999fc4d51cb9962ff601a51a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a29f105e349147494641a7abe89de74f5b691f0d57262d428b12dc536145107;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha450053d26d8db7607ab2aee93a971d97a5e6b9377f723a5139a25364b23c28e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab0f5c99fc6a2418b75fc015f96eb2f84545c5dafeb6e0494837c35bdd74c0d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcaf8c8738a5fdbfd6394bc5efc337f25c0ff85b268f1a04aea0dcc54900fd22c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h29cdbc3a5d48f7d64feed5dbaba7b7855b22187a3a448c72a81f03dc83ed2c2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4a469527247eec2f58bfdebdf423bce3d9ab001b5b72836679a3f7110c9a3c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f49f6665466750c4ddcb7ec5a2006a74cd7f8d350c188cedd01b01280d28781;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17896ad8196568e29803d417b047fc38a9e617227aa087e8b4dc271bfc6cb0ec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7cc84d5cd8113c9bdf6dd66ffd1f92a642f14ca7b75c7a75155382ee72d1f5c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53cbf09fcdf9c97317196e6d7db141d4e4bad1df1203b71202fa39fc29ca15aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf111a98fafba2c2aeb8a099d4a4619af1efda198c0082fa4b85317ee2c0e8b5c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41cf1fc76b191018bc2b19e13a6e8ca545f0e0690deca8862dbede4ba143607c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a1c7b10ee6ce274f19ef59ff0144fba824f6bc5166a7486d29371d35cbe821b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41de5508806086715ae02591957da11196efd6386efa84bb20ee8243cef0c632;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36a8263ac29724d83e566333d8fd5ad121a6d8f92756974c399b04b9d3aeb235;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20a565c298facb2af67f77934be39df70259191f74407c2da3053322b63cf9cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf447b4546feff5f26c9c5ed61ec745ffba73d418b16ad9a3040550d8d96e9403;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7435caf0486d4f003f4c4094fe56cf1b41584f2309ca9913717ee04342570cb8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7967b37110de2ef648b61416a33699678056e7c8513fc8384d718f1ede2cf696;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97553363f94b2e2704bd89facc72f2ee9c026a3011ec4af80b6a3677acf76cc7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9fe8f64307048526a407a0ab72d7d500b0a8dda54aa8d7181152bd486a5ee386;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1eb4c4f2f1db8d6584ec4de0a609b5caf0ee754eb54cc574a94415af3e65e7b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75ce48b9b3c819baf6d035d06f3862d801413eb09fe24f3139a7f8ab6357f966;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3acffd61850c6ef65ced35075b0232debdfd021798d7cd9adcdf29304166c05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h46aafc8d5c56ba42c48bd578cf41a403cc98e3912db91f02a8b0ba822824e1d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5c204f99613bfd92990e541b4252848b1111bc71a21bb9110d9d4dc2a688fdd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a93ac6b2b015745239f426198f1ca5d410e75372a606bbc374b1f42124896df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4454e6fe1806fd53e0706d4dd1d8ee33faf78c6bfdb9e813b9e990da7f5d4c01;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h993b0d60c0a5b66d520b511df0a6bb88dbe98c26058d0016b2355e0e16fdb901;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb60721f6f896954f779e96a30d9ebf3906a7aaefe19c2ec875b2a2e22c6f541;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45eb244d9ddf041a62199e9a0d96670814ee577a529752497dd20f4b654e064;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb7a3f924c803123592f1ff23aba646dc7d351acef975f0527d6f0f41a2c0e47;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9b7ea02a22f17dc89394ad10f2136485332bb5a47385c9f2069ba13d504b1ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d312edbe03d100e743c0d84d58de4f7859d88e491bc88d01aa6cc4716413f68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h489ff75cc0bce43783f697a09325414d721927ac857f6c6f200e40662b37def5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1610475c0798953729af801aff7c69897f04a4b825a9ac08ef46c0837f624f91;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7e0667a521892b22a001f6bc367f0d2f63fd319811fa4da81c565619a462cde;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45f05e09e18176b70604c5e5225012818592925d74cfc41e70a2b90c121972c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hafc7aeb9b2ced9c25786892f27ce7229a59ae4d68196a65758f9ba761772d3ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c5b5c4c9f35538573da304fb445970e6ffa10e5e5af42786fd15affc83f99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he487de48564e97f4a5341ddce4a0a5915a9963b2223d5598f315f5d1bd7b7602;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae4a92b5f73c104591c650d579b127f445d439760463b7cac1116d1086116468;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1f116cbccdbfa06d58cb073525d0310afdbe45ec24f97e91fc227bedc17cdf7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf27b9291a3d75041e94d393a37fc6e81e0d250d866a37bd85d098ba42bb6a94e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h491a983be864a44469e4231b77375f9be33256e4485fd108c45747e13cdf77d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1fb1db9b2481dd520818f6bc90709d7a3c392be639561dce0e4da01aa0dba4a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a23c5d13332a5f5e77e8c528347de4d36cb5157a35ac4cf38688ddf676eebd7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h100e72232ad39baf502d068ed523552e7cca4531ccd525a3b8180590f890f316;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70cebe1e038ad5e870581a1eeae3f7da9ff1908fffa6c1057f994e0ad77b21e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h27f59fa3b22a755738e2fd6460e6941a60ab7ea88c748444f1932f3fefc7eac8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98ae867ffea5ab58a0a243eb37fb62755590c2373d0a01308295eac2db2f56da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44a8c0f7c90ebf80e094cee56f8e4f7aa666dd18c893eecdf24a53ed3ddeba52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc22abe891ff88b14fcab514a107038f26114d693c286c35a44745b9bbdfffc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h296adaf892246e1fe4daddb19746ceddd26669b540362ec30fcd694142e58618;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2e0d7e7c1d62f91f9d82b9f52b54eb378d9ea0bcb337246394b5811bdf65961;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h735de52ae020be6aa4fba23592db953da0d36a73ca1241a083fafe71ffa6e3ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce1188c7ccaa8a94c10ae30e0880cb5acb14824148adbde5fb6a54cfb56a1dc1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9da96868e245ee410df029f31e644b0c9deec9fd1e8aa9c42277494976c7e411;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hddc8025598c6a1b57d7fdd8b93d4ea63f3aa3d9d125f2eef5ee40da29ba4cc8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90cf77133234b871d0da0d48fe8f408c47f626a6943bd76d5000bc70e4b0200f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72d4f5853a1df3f847391be40e540657c055e0cf9a10e86fc3fe0bc7e52f3d56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39a4dca55a80d2e03439a075a252679495ade49fb0acc6ed23e9e8e028452db0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2458b136d35501db5007770d4edd2bc93f7fe48e2dea2cb2aa01bd5a62e38506;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9638f859abcb16901bc7775d4a070587b4ec329785c4b537d0da43a8e80048a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1df0d6d82d120e36d3370e4dcde6420d4a99d57478ffa91b5b5e1276d347d9ec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd65e2e7cc796eb189e7818eb66e71ab3773852f25d9a56f165613f3f3faf053;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0ccb40b3ae6e31530cc0c5e86b5c107c1c90d355525a973810c1b739fc089fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d65eab0536e413a9b88746044e5bfa4f077edf9ba0d80296b0f329878e25354;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38be0a4e00484a0cb43fc3d57aa35a566afb4618b1e033c44b8fedaea2a63bd9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d5588fc6869c64773758000e08f57d4a0d19a35c1533517275f25f05fa00a07;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h551f85a6b68f23f0c07ae3a28255cde3478d3839b5cb26bb0479c8328417503e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa32d46977652da79e77d62656f2a474e72fe0e4cbc4ad2a70bf722121a7d4fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5c8a27c9f89b8d6bd30f9a8747e6d22cef748e467cb4a7f6b5bd19a6e12503e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haad647328520caa9f67d3b71904fdb632d2872414301049489f2fbe25012b3be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17a4b38fa0e514ab4fa01838e9ba793f4ba30125d10b04c38c9f8621a4ec266e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha1739675a2bc9f63118a241ef64938bdc0e9fec37afb37a0eed372f382d4d620;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3887716319b452ab6bdd9543ee3d9659dd1d35c9562955e65ab48b436be5282f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3575fc6dc157c4ac9cd87914c958b02615233e918422b02d5d3cd1160e0cf1d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf89f4964ed2dbb6d2cc2b5e5f320dd06a89e9f0fd5ccb7bf21983201d48a3fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71bebbf36f7b7d824d35727aec32c8de7305e46ae9499ecc50a225b4aa58c69a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hafa6c25f74299c0f1757023ff51a0e34f20e3601d4256d71d3d5c0d7efdefb3b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha26dd86210a4797997ffd9d127f52addb9143a7d3a6a9c2360c0f903307343df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f52a42576c920d6aac49af39e42a7ccdb89340dff7c4a3c8e887697d7d93803;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77f16ea327c11a8a0c9beab8519f50683509928bd7a46f19d97ef575d05a2e5e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd08659a02e3edf52bcb8edc92f795caaefca4b9d107d8612b4babe26d5af912;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h597cd6ce72b05048c3ff52e5955557d253c00bc550bab638812c94f2f213cb9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b28616cd2676160aac35372d271496d8ede9924ad49c57c176596a3241f9200;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffad60fd1914831f84806c4782833c425553c070c3ae7a57b83533e0d3b9eaf3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3bd85c69aa8f593f4498893d31bfc71a0633d946e14a4b3cb23ce4234c433797;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda36263860a7253a699ec4b7894919739e4fb6ef6922d2b3459229c6c69de025;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93e0db222d3ca819f481e22ef440c16abf8c428fef6f0035e5ef23d097304706;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83a655593137dc9559ae6d4a5d702838be34cbfb572eb85e08a825b8c0989531;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15f4032bd91ffcdae04df67d1418206dbc09bf2a645cb04a15eab9cc36a7987d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96cfc34f1c3428ed8b15334baa6d665389b89ff63944061b7b5065ce1337c6b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5039bcaf5113861ca226d82df5c673394ecf4de887505fcd6686cb3d5be7d25b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2437bc7db4dbf22676bc1d93b1088f723e8fcf0d061c0dde1993136c04c41152;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7820cfefc2b309af6b05bd2508450f34f1cd121688af3221786926f4c0de49a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h443973dd5c15318c3b17d587f7bfe2c0ec9a53ccd055471219405fe08e7c7ca1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7da72b958ff3e5601a66d4d8197fa231785c57e66eed429f5e66b375947f09e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd41a88e7f0a2a17590dda5b2b6e304e06af66d743a88a6a9c0ccfb8e62a4f207;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5d264b933750dab85e14a2d0256fd1165b48f8eb43a391a90470286f2ab37ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h130f83eb7b6fd7f55f279b642562fffca84a2ccacc576297f0325db270393e6b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h13e0f4e552b2314d9fb3fa82687cddd61e428103815843ae33e7c4c3574182c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36e54ec5c8c2e4c96cc1a25ac1b2c189fa43f9e9559b90f2da40e8359356273c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5aad14f3e43cd0209ffd2771697e2d7135c3953f547fbb2bb9cc8e5d5ef88ebe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd641f2da498de3b77b401f01b1eecf08579dba53655999d8d41c0c811c392692;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7a687ea008057c45c835efc382f9aa9bf90ab202d03309a7807d00f1f248846;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h18f639b7ed63196eafe754d34c29019af37a903b49e9bdc6cf9c784738f1ba24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h827ccbbc6cb5c1c8cd462d3a085dc0b25302555a88035a4659a69b2b47c7dc3f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94f727aeab9c42720823da82e5948f919ede35544fb1dc5c83de6cbde3f7c52f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4eee73a10fe232e9a9e711daa754354891d372107fa75265ee1084f9c9d99e5d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6bc8f02435272d805e5b4d8e084bbc38f03a7e4285bca112318d88ba354e6c01;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce36462de65bbe5d7963eb644691d9f68d1967d4d11c0b4844bd435c4d9ea6a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5826e071af8a8fbcfac58d8f8d9cf23048dec4da7434d8970919ef0d8df97959;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98a68e1b69f8a507bdd1800336e1d64e2810743d954cf39b221802be3095f0c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8587e91e56d770502c05d54fbbb8515b6872070ca686663089f44044f1f008c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h311d73fbfa41c0297d42fe59c96dfffb8e7c968b3a2e60d2dbdc41e657e43650;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ab3865cc782e0f4ae2debc2599531a24808a35d47e932e93a6bbce444ba978;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63b9cb7ddaa808aa714e0e95f190e76d46858f71c675f26053111e1838c1bdd2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d2d50483da71f5db29dd393636d17fbbd721447c34712ff0fba6e6b21f053f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h253a7953b83740353893389227c2eb3e315e7ce5f0be33df779734f0b5127b0d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc650c30be31aea4312f30bba21d12ea6ccc6ea9cd81b4a970b6073d08bca9b8c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc86b969f84f2d3b5101e34dd00cec9fddce78678f59126b2c10597672edc2056;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63e6ea8d97bd4ced9a1517638df0e489690d5eb8701f5cb161343a3c93846fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h14d6dee64a8f8028548d934d7b65e74bd2bbc684c872827e73fc332144aae82e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he337c4a0cb7bc086d76f5940134c54e9a65f205fdfaf37c25f6ea3958e8f4b0b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha68e66eefceef70e5a9461a0b9cf3256d5bccf63920e967b136ee893e77f770f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab769ca57c98a0682066281913bddacfa83d4f5e9c81a4a1aadf033cb0593b1d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5f89c7c05f7edadb0ca8f67742a78ec7b2f9f7abd3f71444faa4f53d4dd4bc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9542301fc55c5365f430110e3e872a32e51c8c8a3fd54d0b55bd90f3d1ab367d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f6f33e25ea03cfb7283ccb7c7766992dd8cf0d6634a8df4338e80bc2f4f6249;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcec8c9ff5a2812607591b4ab570a135aa49da4af2f04aabb17918c3748b06432;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ef7a7cd8c0e21b164fe924ecabf1ed4c18412011de9dbc88d97a9e8af77e9bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee3ffc408a799351e0d1c64705e5753802e9ea4c111724e1b0c1cb58cb03b463;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h115f4d057201ae9ed3eb2bec906ab71a647d61a813aae0a1c9364aea117d0ad6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51a046453b6769c6ae83ba8465a77727e1d0582dd743edd61c29ad8842eb0f2e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5ef1e57b1ac244b263c6925ec35fa87d71140a83ead84d867bf49dfc25ff067;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77fcda05a1532ef1422f6c62b1014f0157ecaa31dae9657a474a0182148fff25;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a94372bbc8d5833d464be00a8ccc7c283ac7a9dde47fd1ef76646f2fda8a235;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3db1d9f528b439a361b944e474247404afe0cd7934b8df0b06ae28d283918119;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfad4fb224d8b94cdc1db0998a9db82689fac45898f6bfa127bc335f6db01b1db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba11e8d68d1d99d34aa15ed74971000852bd3f7e52a71747237c790a790b778d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ee60ac25e288de1f2572186b6533bcf32f7c6193bb2679e9b9835ed6abcd5e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h733b303c2c9033b98a1f7da7a209d7701219353e3d8f29b47378cac5072dd544;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h495af0557716b0013b4e281ddbf6bbf2fd44e58deffd1491a10e02f21b08ac45;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf03a307ec1b856e7e601e80390ddbc1d666c49e8c1af95cda617c8b167d851a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha78386c51dd61a08178ad10bb1ece2391a13568eb30f832959a3e56a1eb8dd36;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h714ba8edc685c9d6e6f95ae20accebf6f1efe4900738591482c761f2d2357637;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4f453cc7d6080efda02430fafc4190401b31cc43738aa464457af26c1899165;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a41d4b655eb1e43eb3aab14a2c08fee35018191f22ce7aa35cbbd7c5d40346e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53624c91e2d7f4fbac45a5159f15c5411400e55eba674f1861921a583e890561;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he82765ebea76ff39a32972525a3e969d3f91e05ea39f70eef2dd7fd7626f86be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2fef415c73555dfbbc0d9f66da3d1c57fad03db167e0ecb7dc99f7e098e2925f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec72034d755549411114396cc69e6c8d097c2d4778d5ff415914037e63504131;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbcc20b3d6988325747a2512f7463e50127540291fc6621aa48a49d59faeb9b34;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6aff33c7c12f4951922c4f3163ef43b1ee156f7e40062ed95a9a23b3d66362b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e3579b0e8675d97c75cffb1ca9ea6b1ad3aa28343440f475350b0ec832477cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb3764d9c0118b35d7a4ff3c5f427bcff51a36771b110f84a1862d30efaeb95a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h34fc937381965045802cd880f2f65a37bee3b32def980ae4a848a72085de1b34;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h682a74976f7ebf39f131b996d4a0966a0787f1743d9169dd6ac7c82d726ce273;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h289b2d77a016b04a3d75b94b9a678f98d5b5a230d1d8834ff5ac2dd3490a443e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8aa49936346e89a75af9eb2859b7301b37956011f5e28864bc5edfb46adf36f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71d92e8ac6c1de2830e0ca8deb5ab01bda1916cc728ed46fa74b17bc270c238e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf1e0103e362d53b3fb2f9c32d0c91056cf0da6b38ef57fa12b3e1ce902795ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a043a08ac70384c9602e4736bbf0673e05ba4c4706c8a8c08c2e1b80f265340;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha50087b3c69c58b4b1986b3c7e46a0c9641ff8177f1fa3aab8daa2d22991ce4c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23c7c33286424e61c1c85bd82e9f6fb0dd8685aa3b43827c5f8ffc3618f885c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h76c66ac28b17f77338cf6ed77dba23203a0bbae46ec3e37a0e4d777a75464d69;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6636caa55fe7bc9b0a7eab139c4b67c0dff1e198e779c27a5f52a39de351a4e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9317c4cca4198722f3388ec1564bf2caf878c0c355002a076dc9da8ee44eff15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4961f420dac96db670e12da1663ea28bfbb56b35300764f2f909333c736f449e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h423f3b29ada4d6702d590205d39991d8899c34f9294e6731651b9c106a8ba92b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3935f0a46e229481e4a10772c748cbee02e481ddacd0641de9614b5849f09acb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51011f694397cf240488c2dec7a6405c8100ba3619a7f05cdafc760bc4747bb4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcaaa5007c330ca4b98476863e99278ce02ff84d609556ea3eed0738d8cc1efc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h76d091717ef9b90b674d8417210f0846c304c7974cb835fdcb13c609cbc0c81e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcab271004551d816f332f574647bcaeebaa015b3a22c751aaa73ca996be77ee7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e83ea6d67bdd4fc7eddaad4b5c4f24bc8e005b3fb4d1c5ec5e4616dfb85f4ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h109ef6b7841c397409a1870d688987ed09d4d9493b38bbd236b0d862ea4c562;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0c8a5784219ea1123f3b7055ff458cb40471b868401a466b3802bca6d39151b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5dcd0bf4aee834576ce5dc7f7c083b4219e892f717164b2dd1b3df090e3a4e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h322bff18a5d39bdf45b6a3742a828fb0c598e50cd74455978de07910bc058b0a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92234a9efbc3c6ef7afc8f0dc7ae6ad90795779f248760cf39994ae7cd82a962;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2159e101a8c825856761c5abd2b54496cacff351f27f903bff326cbfab657402;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdea846736c27c5c120d318e2c9f89e3fa32e218b0ff8b644763490b6b100e723;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb83d44cb3cbdcd8f04ec054ebd20eaa855c6f05d3c6e6cc7027dd5c0dc82a02;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h18b0b79db0628f64dafe60dc2a56749ac9999fd3e7485460910e5df5b0b2a24c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h547fc2619fda0eac3df5897823e4420010f279f2208209c1f3b5b1f46410b6fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h681045e3fb27b52587de9c687b3f210efb07746fec535f0c5656c470efbda8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc40eafbcfea3e9f7f3a9ba7a7cf32adbd26390d362b09b2db18d9738ca5e12d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffef45b255b2f6aa0b8ee648ddc450e0b44a61815449ba12b42e374280facc89;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h839e8b8b800ef0d9d6692cd7b2d8cf24d31dd4689b9f382a177814a49aedc55;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h554a85b73c5e21c2c3debd519391521953345e4b1fd95535d37e319df52082cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb8bfb9ad60c81dcba51b3aa5ae0f50f2d0b7763eccaa80a708a0c23cf2964f36;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17d5c6759337e17c032299d5c7a4527078c8ae8beb864abb5344cf04a514849d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hed94de72283172cebc85c7b12f6472de1cd3ae23f4b8f0ecb7a639c2658bb77a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38092ab578abdf1b6ba928e6cb9d7ac8119684f38876d29016f3f0b05dda52b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha392bebfa387d36c99d5f87ec8524e2a7e2c48f1e7199414520e64c91e0ad2e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7dae0521d2dcc6dcf1aa72f4344ff473ed7e6df7c3541d43adb866d41b6c1bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69348ebdf7fcd4db4e40962410d8967f00410fa135d9de1ffb94604903d6829f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h237a4d63490843b639e3a2533a00bbdb4adb474e31194d6ddb5118a368307f7c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf0116ff1179340e4391255a69668b1278da617253fc58577e5432155888be09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6251c9690a24f56c518cacbd038d91f16eafc82c81203fba5882cafdd46e708f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a2e56cccf75ff3852c3e69b491900ac29d7da785eca068e8bbce9d624f28060;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2799393c3ec1ad6ef39f3bfb25bd23e43bb2586fa7a559b78e76e69a6d6b522d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haec12d4c72588be272c7ac134b264daf8c59299a3bc7462dfac89bc958607c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8be2230b9a5c387418d9e0f42909cfd4fbf6da043057cc145daef93cf72b725;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h13af776ebc5c21cc100f3957aec2e8019fe7ca4d154367f8c0f897b41f58242b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h422951c963eb2df92d898d64b17f4694c8ce97f7fae129cb44734500c26905f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h788a5bc4045bfd365230a785fde00ed3bbc414193d960e5fa9d51efd720a5201;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h67fa271c79b64d0235a3b08eddde87097e86665bfa9a87f50965dbd726e707e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdf2d975fd67938c8e86dce2c05a4bc3165f4d0fa4b13092aeaec4fa5f941d5fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93af2b76ff88a5475e92bb3e5b2d9711d57301556c710b73a9a65517bb5e3d4a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ebc47fd31529912422a9ef4c87cde09f576ddbd0417e71d9b9273b498c9de08;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec8b5aa957fca97acc32c6a64e92906050647827842e52b48b37b1a0dcb3717d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70a6ce5cae0cce9aba58d33a7710059f3a9a395d1b52d2fe4865207d8c015c2c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1bc49f8c6bc495e2f1b1bc072ab96a5b134ac611f713cea4d4b27db86e9e0a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1093a8905d01f31542aa0c23573324ff074cfb3b6db7cd10166d7a0f63fa8b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7fd172b47d9b6630485d806bc9e2718ec4e99d1182bf224318ee1420ef44c199;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9378f315d5aba40921ac8f134a7cfd3f8aafa7675338ea21f859cb1f73805579;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea40d4bf0b9beac3e46b490133e33a8f3b1223915e856884ca4f56f4b76d2eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf25cb1918b99341866e7a060aeea6177a53650eee17018ded7b08444b4e20472;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdccacf991f87c1be89fa79eb839afe8f5a1314e19b6b5a4f339682587d92fdf9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9d988deeb5f5da4948b7c1209562cd92e2cd0917e52b96b7280275f8786f7cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he38cbcfc65f1164bba69097f44daa988a1602c031a60239c07fbdd3360046dec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c9daa4aab9bc4d06b0ca121ca27d6dd5ce9c11cfa24aba1642e326115471e69;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce3d0a47ff4dc0503ac30fc97a6e090058f61a1e6375fb2e68b534094efa3c8b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb696a7d9cf146a12daff37322caa635126c7b1c188cd1c8e790fefccd940f89b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac27ccf55401ed1188e57da2bf6010da54cd126781b77c7551a620799b6ea87a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba28e76e84a9f5a08cc5af0531b41c6c30c4f4ac44582b960a642b996a650d80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a4a9bbf7cad2fb3d55c670e2f039fe6b02ff86fd5166ae3e49967e6c7fd9a61;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda1237388cb9310fa6a102c176db658e53ac8ad30321fb99c3d043248cc8071b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b0e53ad0df6fd71d09aa7efd8d94d288b765ebd201eed337cedc25e6bf7cc5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdbafd573ced9380e072290c92bc28b21d82b6ffc0aaa39417c2ccff8e6d80119;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20c85b4a1b058075ea464e4e393c2da05d0d05b289947d757b0595aa802c6f22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28b5ff30db21f44d744cdab3fab8cdd06852dbb42c53bc5df04b12076080c89d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6551ec35adacd42acdb8a1b7f202369c7b10e61e6329be2674770bd9ba7208f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h18ff05f697db8458fa55f03f640ce2384b73cc9a16274399e4c314206255fda7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h203d7349e334998636a1ffdbaede5625888b2c564733bde15c05fef4d3f6eff1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5ccdd7bcb128f8daa1c30b7ddf5c64aac24365bec20746ddb21c3cf4f4afd613;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb77387c14aedcbc7fa337a6ae4ef5b4860e56cb0bf479df501b1437d1123c7b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb47cb15116702a0cc7d9b429157a2ba26d32397bbc05e0ed02c4cec0801997a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ee03cd6b1c8bcd8af24dd2a5dc4b098b623ef420b5e55eb9484c5d427da17c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ffadb4c2fb8ac33950d9e78de5338b2a26cf10d74bd711ab570cfd734d27aa1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d5109a241555ae369564ce648ef26328be1104546dee475e3e37ad11606243e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb7db49fcd86ac4106c7c1c85d576d7dd74c1aec1454bd5e614ef57c850a3a2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6bdce630097e0d0a90ac9f0a5cba36e61b77fe8a34d89bbd1435ba43c993cac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h759217a7744ab6aa94f1e38a66e6f6eb84e15773f14c522e76da9485d48e30d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5447f74e85338b498cd6f30be5087f8a9f4765d937d81b4867762210f97d9d22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e1ceb00d998cfda35bf38cee8a800600a60842e2e47521b00d813e401f56e7b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc4aaf46690d8dc2e797f5fdb1615cd365d4175a6fa26b2b943f32023230fd6f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5809050e1971361bdbbef0db4b17071a29b874ec8a1f7ff4cb8d998a24637d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90a65e616519ba66eef740ef26413c8c6eaa05b7ffe7aba3826c2368c35c4e15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h568f25e282164774869c7fb93a4789bae29933ef996ef02cf2cce9f68f486752;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6d2d2f2b0e9ed056b44fca0e76ccf66bfc0bdbb907b9a1f17108f152d3b5b303;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h421609b2247e13f195a6874a15756d5ca1b2046305950c7ce9e62a18eebaef76;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he75f1badc3403fd686d25f06e576223e68b72793443f97138c702d8fad7d2af9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heeb0291166c2e138667cb3f29836755cfc40b44b46a3eda7f5e49639023f26a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d23952bf6d1d9d1a86b6e82e95d464593c87047e1703a3960e944a82647a681;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h898dc24a2e86ca06cadeee901895b68d0386135c74420d345b4a6f0eadf19b3f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h406b64759f017e1b6ab2971737a4e4b6fb3b215c4cc37877779be9a46272b4f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f9dac9f78ae3786fb1d3a05a2187c74a8e6c68ffa47e47bf85a69b19ca882c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68c773489a28464b8f664e6ed9d5397486e44070736079fa2533566566ac57aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec5152d22f90467b0c694ac7d6804f761fd0a5f115b5acf1036a44c3534e1557;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h323526d7388d90ffc58c813861e1c7391fbeeb1b11c609c1f423940ab22d844e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e67ea8b86179bf274098530d59bf22525f25bb65f63c90d61a0eebc7008a21f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2982805dbde3135970f5d934df2c24a6b807ac860f1e30eed84664f3fb3d9502;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c803cdc56525e5e06d94ee43c6f902ee8b3eb5d0429ff355a4a26e22d845697;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20a24106718f2b63084e2dffaa4f58cfc8b93c47238793290157e715415ea940;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h370f7b479c0369d88eb1607ffac74df0fc3a2aa656a9dda2a767c517a22c11e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92fce6544aba849ec9bd5f058a089f02547acc6b75587766a9a5dcfe2d47c072;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h724841e261f8adb2c2043afa74eba000cf3d39cb184e168fb575899485e64b80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66782d009c74bfb5e3defe84f8d8120d63c7cdec256ec3ebd23b11b4ddb8c023;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b9961cd96bd3bf3a8aeb541ebe7f8d32cdc8696846d044a9b500ed272325c18;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1cb3b27c94648e6783d966e4c13a70def849dccccdbac3ad9a0aead7308f61b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6279d6276ff4dfe2ee3a83f7ce4eddf84a1f4d978659a5ad6888a113275124d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h481fb4d68f12cbef8e34c8e244a6f405276e4642119098c06b8d0bf028ef190b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h95583fe0813611b004a642907e6d417779efb352310b63941d678dace0fb1041;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4a272f24901eb932a5f4b881e8363c5c46ff0d27eeecfdf7af0d2eaa423fb22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h717889b974779dea0f90eac7a6be6f97c84819e1d763b7ca8f28904b923b3b55;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6825c43c5f535bb003c0994cf60c1ac7581953953b43b338b880680e7e35ba68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9331cc2c28bb0f7c74be5f9e984d6ed1c6908c11ac8d80586291e59e858e7911;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had41d9dea62594db21dcc1dd76f04eee1a104e86fa67ac31bbe9596d4d9a433b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h107d9ba5b2ef2b7fa030b02ea7ff49aedbdc4934dea1a19490f96ae71babf7fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87b4552261015b0bc666777ccfb6526fc4774ca792cec762d1b355474a0ae3d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc33af3171bde492ca78fee80dd8f437713d1271ef7132d7a71c3b098ef846fb0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b0944757dd79f018ba119ae414290b0e64d2dc79f34cd39f5ee6135402cc7ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee0690181137f71b6d0caabc3cbbd37a19fb93cbdbc43ef7b21b70687486f1a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7f1af0e7c24a2f77e1eda29594dfa82db00c9686a2b58bf7e58893ccb9810a81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h278654cb56eff46958b2e3528eac42ff1efc33b1877a5cba865c53fc568c6e4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha97fe5aaefdd3bb31f6284340840d5b57d81299e502440498d373a9ded147b33;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82a91cf97af22e68c6f741207c626a0c62efe49fb2a028ccce98649f057ba55c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ea68dfc9d5b02c9384d63a3fa4871d7bf9e8e30c9173bda322a327eba7a17f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb834726441921e9990b4c6bbba57d66f08e364da21520787fb02848230f65451;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31aac6822b6d82d0b19c48716af9418431d756778a3a94addd097302a848f47e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68bfd4fdd51897a9144c19b4365ce261ea0219eb541994b1642567c546d55b28;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc54da53e3e4b8afbac62873a2f4ad84f0d59017f9fd1a151b5ba60060559b5f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15d14f206f2245508305a4676c5408b424b0fee4f68005f973eee82e7544940c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75c5ce4dad208e6332a5e949398ac02d48cb8c3245400f168ba2b7e5c40af667;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1af3fd9a1af075a2fb89d66cf7adaf3a596c3da4acb404c97f848771a70f7ebc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf844cac1519ed3ea9dedfc9d67e1b8d19a47f70fc86a8bd648499f85efc20147;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1c44f1ffbb80333572297a0793162b8a6229b07073598e8849e3f9c7c29289a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b384d227a27175201da8a5e84b18d2dfddcd244bc50afb474eca30d424802c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c2054822e98f828b8ef2886ff2c31dc8d60bd52a60de542698823a978e17bf2;
        #1
        $finish();
    end
endmodule
