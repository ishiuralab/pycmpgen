module testbench();
    reg [30:0] src0;
    reg [30:0] src1;
    reg [30:0] src2;
    reg [30:0] src3;
    reg [30:0] src4;
    reg [30:0] src5;
    reg [30:0] src6;
    reg [30:0] src7;
    reg [30:0] src8;
    reg [30:0] src9;
    reg [30:0] src10;
    reg [30:0] src11;
    reg [30:0] src12;
    reg [30:0] src13;
    reg [30:0] src14;
    reg [30:0] src15;
    reg [30:0] src16;
    reg [30:0] src17;
    reg [30:0] src18;
    reg [30:0] src19;
    reg [30:0] src20;
    reg [30:0] src21;
    reg [30:0] src22;
    reg [30:0] src23;
    reg [30:0] src24;
    reg [30:0] src25;
    reg [30:0] src26;
    reg [30:0] src27;
    reg [30:0] src28;
    reg [30:0] src29;
    reg [30:0] src30;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [35:0] srcsum;
    wire [35:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12031257329357c503a754847d5ac5ab4f4cbdc8c7b9c5556f71ec5a1742ec7864fb24812de76537a2760f9c2ee27b79279585c1afda22a5b714556e98932ba2fb3661b84fed6408c7c9d03b4d668ad83c6c036f45f0595cb6510d8fcd472eef2db973692311b4c4513459d8318c24eded87329a55d870337;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hedd323c8d477d69674ca50c8a0f634f7b47022897992887f50acdd48052eb1cb7bb49ba488ee71992b365ae0635afd4626c4319b4bc63f2600970c22a8c897181c31f96c402e0fdbfabc67077baada3a64dd0e9324abbcceacf75ecf2a2b42ca0a882f11eac010b1a488d6182531b120aa53e867231c8d51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1682804ac67fc6839debdf9f5feb0b2fb58b3ac7476f9c8d708021e07e07f12054980722369031108469074d77c0047aacd18f858479f78c0e07b488d69c24ce9076b988d2991cf4fa22e11b75dc9a8fc8124ddbf4cffa34e6db0f8e390d6f812eb3f032f69d279c83b81e65dd554e4d66edcfaf25533e91c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb48218cdad2a9b6f0775b4235aa894a598853847f7ef5208422652e90dec4637015a34d081b948b48fea28a7f482187fc4a18197cb0cefef5edbc55fb3ac7718ea346458b30411cbb53c4e495039671cb980b7f603424976b40c4b4c4d74f58d7383494d58ce562e8e9bb13aa5e852e53b75855e642ba5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd2a39b367e5683b009b92a5126839cb471ea0ae13a38166219aab6316dcc79a22f5eea3edd0bf85e3667739782976503b6d9b3b13b180293afc020d846e5474643acc8d1e9ba1b90e7e5668fafca87f421d1d451e855614da3167ad9ef0889b73589c87cbb03968953f64b933cf8f473b21d52f844c4e0d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17af821b92935f7b61fc9e7bc0c29c0232f324253e84149f35efa676714e4a2e1433f43a555b528d574e5ef061581fb3ff50eefdd7df08245dddc1f6e98374e8e483b65634d4556b9a4bc9a5850393646814d33cde990ec6e53e0d20e2053879a28fadda1fd6f9a83c753ec90c5754c5504b958a7991666d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5bab58d4ca03960441641edabe6eceef234c528257d3d89b26e877b3da3c6a7f6394c6a06e7068caffc8a1538d39bfa5a37e7a2bb86d687d366743ee52162f8de03590521a180571c397b2e46f571db3499130de60e621e61b5f1102b1c9a4e7ece5ab09cc0fbb7c63ae7450929ee0cb0a28d578479efb56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b4f3f65a1d1a30a73e7c74bdb6188cf46925004e52bfac2466a1e98eeacbd64756dee2781f85968f70b74eca773de0689cadc49f090308d81fe4e4f0cbfba0074b48a3b0d1e5a54fee20dae531c869607a597758bd946a4aa480733df8f2d6f1f2f18bfc131ae8ac76006a58922742bd990a709568b120b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c6d8077a2488db67b325a4f2551cda22984087d637ebfa2cc442e80d089cf2a72c99c2cd8c1ac6bb808d7504d39ecec71acfff720adbedcdbd6e94eb63c5d92bfbf55b90b71f0e0bcaaa4fefc5e48ad9c3d5dc9201c146fa3fd664cc3d35dee70c256969cfd3a6267ed5cb9a7c9f61d833ad8c3715fcfc13;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf62b7ac8913390c611dfa1af86dd7df77ccae79f204cbf66604f3d3e43a5a377727d10667dfa96ef03aa6ab3f54937d23457a9d8e7d042c29726009eb0f013643bc8b0b7686e5da5ca3f05aa8d1987d833c33a24715ea919e7ae0aee0d43e4e03c339865ad93684b4ffe9b91020a22f0024544f2f06865;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1215cf1e62d5c35ecfad8192cfb92554d3932edfdc6a9ba34d6023cef3fca1a63c1244847de5ee7889f8ed6f15e1bc4130b6c54835368da3ea714e525f66382519d0a41bdb0d4bca025588ad899bd49c61fa9625ff7d6026350567f2a953c723a157d59653d6214bd970fa22960252aa6600a80e03ea29c2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c8b2f367d01013e4ea4d0a21e8e0f57d4603008f6b47f2b11274e91b04bcf15533eec5bde29a7810d6af9ed372f5ca981e70600a2475632770644f11d1a98025d1bd5cffaacf6446ba4709bef65300da32ac3f263a28b8846a6178a3b157ebcdd37a418181905b9fc9e21cca07cd7fa8f8734e7e4dbabbe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d5d889383083dc3560780b4704404c47a7ed2fa0f6cb59578acd66692a63f45cc7293c12c8b351b778e57f1da0075a63683b3e85ece790a49c334f04c56a28240ba82e5472aff06a639d7031292bcd0e29f296edd0daf0c8865846f15e0b73daf6c2aa0e658b27f09624233a8949610b0f46c6f1a508f62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e6c2cc5668715bf174aa1e85cf2afb36e18b64c61da3267016cc642e7dc0beca13eb2ffb503813a59470dacee4db48eeb884d7e41d4b2521d4cf6e9028c746d8d599ed3e9202867fc5148e207fa327760d8e3d3d627b6acbb4e92b28afc1eac47f2175a128dda7f300562b3e298c8942ac74143be30bd07;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9e8ab3ec6ac26fa8c11190219a43956e71fbd39acf6a0453db570e5b2f622e2558440e93b8040f54f103e543e81315e7c1018fe4304d2172a65d814507bc4cd3df14b71f8ef91adc60c6396b213ac5f27ba064faf6676769872436a1dfce16855fc4f393d20990af459246e73f5b60228ab777088fdb3bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h167bea675877f0a4ed478680493a274b8836c8b7b11b736de16134ecef820330df9deeee13073f616d921e96235b2cefbcf3058f09c69b6618775fe6eee64f0a795cc701ffeab9ea88276a46ec6aaee19dd96adfb1d3e2875612192a3f2b547e45707ffed530d0e37ad2162e59f4ce6ae723f18089fe88f03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc29664b31d0a36a02c85a51e835c1c8ab6a49881675cef26549324f69c2777651692dd2a4144d2e238c49f6f1eff232c7a53d50dd19a9b5093cbc7660deea07f4bcf02ad7b983f2befb23b18b89235f8435310746ac6be2e8d202e8258e6f7fc730d23e6c80595a187dd17329cc32aebe08ae8a94170e9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12609b21c3895aed9492721ed4f0db4c9112165d1822c627bd402dc5d65e05a56bc78ef950524008685cc947241fb354eb288e968fd516b821403559ce0ae7a2eef36673b7258f21e7d6422da48f457fc80a32e093d04bad8e1f1b4be3483996d78b33f64b5ea8efb274264884a9d76b8abeec25194176bcb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e02f2fcf188c25fd658a67322efd580b3bbe146fa7ada24beaf2160ed88294bcd30b216e18367c17b6ef771235f59f9c6da0a77ce3afd18066f24f48a82b28697a22d37a1740e5ccbcdbfada7c7785d81eb4a40cfc92fa09a4e08fc5f2bc333f64cabffdbc0eddcde70337c0418a4302133b60f44f7d9509;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6aafe37703157d4c3e664fbca5aa80862af52c5fc0bdae450c03937a60382b21370a76f013c83a32c55eb485609297af265ae3dd34db6857bd28ba2957599b2f643974d302e8094c12570302d19e98a1a121216e07f52f6c3f264ede6ee1270923cf93ef92388b0e5a7552f31c50d76d056b23dd91bef46;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h144e43ff0773648863f5a6aef5cc3310691ea0949014a26c2319237598842c943c220404f1ac9942282eacc05796ba6f12adde6c41cebac0921f4c850d16dc726f329a00cdcd6c626f54435c82b69b98bab20c7d25777f8e00991ab5c771ae417588b5eeb5c43b3c9453bbf8041ed17fb947f90aa8566b061;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c4020a6f3c84c8543351e3c88faba99cdc7ba9dc49b9fbf39290f8e268ae17475df0332427d02e2a6eda622f7b99cbaec4f7b9b8849d6ba234e5d0242e54d08b602a3ffea70cb6739cc1485b85a55cb62c5d4218d11443222d6d0850344aff7bc33c5f37652984ab70ba4be0a7486c886fe1afe912ca2a80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hecb6ce19997313740aa46469ff139b35244578c196ac9b2d06899ff7d3719561ccf2f82494cedfb45727e9468a9573d74771ffef058a854d27af3df1875a82311dead8afe3d21b421897cd4132bfcb73767a57ec18e728e508314731ab32ff4cfad94344a42cf07958ffbfaa31ba81e8a3687a45b34261a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h85b969eee20439e1e56e0bb05297eb847c0c1194902b702b1b89e1f0001db0910cbdefdc98242ea0543a8aa7fdf70be45e41cc256b9e1f93b1cc69814cd6858abedc692c902cda967dd5365f26605d8e8d6b79822fc7bea86f966c892c4a1b7e8286e38290614a698a3ca02eaae748efd2283a73b8a10d52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15712c0015fc83c98ea7903679bd61caa133854a07675b7aae3da99bc83b4a165d103cce87b0e02ee66f94335a4f571d1502876d99a073e549619c5b1475049fde221b3e5d459de438d068744df72587c237115340b1ba8f8cb58b5115cdc81c9e877863106ad81c64bfe1e5d168c3e958ebbb80488b09202;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8d8d9499b20faef2362fe7b210a8a0f2eca08f74acce833cf6aa65245cbfba8e4df1c17de16461dbe41d69e592dc2704f26276f61d08440035c3fe47f7790130e1e24f4fb4921db6517ee9a6e25201c8c220916aa986a62a66a2d9d6f4f59bb515fd17a20f27d87d82978816a5eb3e6b11791550878352f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf82eb0d57ee617db8c23de791a04749571c2f5d464520ad175fbbe6b58d0a5b6f76e42f52c7ce1ca1b471dceee6ac5230ea9bcd55bf84a9d1b5d3a92204aa3462d039cdabebe517b81ca5effce140a865383dd94a13db130d836de94c8ea55f83a64ca7bc5961a2f3822a27c188f2aba500d8d246e98c64;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c5bf312b40316fd18ac8e42a042cc2cdd6d00520c6d7521811282ab6058525640795e694aa7679606902a64713275884d436f8316ab1f571a5e1e19004d23ad693b5ebe5343fa4a4b9cbe8382c3ba45da0d586aa0ba7bf24a54a9b2168108b84ada1290d98f3aed35c053638aed9e807583bfa56e16f9f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196d7a550d6db51edd1e049e011f4bdce9a6e6eab8566871a78c3f6df611597cfa8d5dfc7e24e5c53817f0cb123383b56e52e9d1d233a4d64b5a6364a93cb23c7aac8a9a76e0c3a77434ba0a6c631fa9ab9365edf6e51166134dc1be072e942bc48172174ab147a2fc3886b98c0514f424bb5a828fa1217a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8d9da01fcf5c12850b9dde3be1b1c4a51cdbfe73d6f65be24c0c5f63be4047ac32e195fc4caaef0ab6c0faeb5802e95067aa8a0b1285a18b0e9d6b23a5009159c9824cea6ea10f3048d5d85a794ba73ae8d1fd5e00a6edb1e5142b648026ad868a338084e01840a20fbb3488c54a20897e7f95a26b50468;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h92d0e9f6578e5c20d8fbe9b2d4771900f662e8451610498c6ac3a2f73a6926e881a6220b3f1f61e252cb3574a991f80892f462fe6c96362a544be69afc2c6fd2d2b4503c57621ca23c6613e5afeacc99e553946f87fe37b1360c621f78b774fbfca88718f0583926040d11f0e42e62c733c732d2fa655cce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h131b46ee9ed21e090bca56836e980f7c1a9ddf75673d217bead5c25c89653ce969d4a53e04107acfaa1f637cddc98cbcaa912e36774aaec45a93d34bd5b4bb98ec3ba26185f287a520f714922a3c93c30d6bad7f0d7ff228f70a77e04baa63d8b39c43c940e9345bf29d3a0d07d33a45e819776c22623aa81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1003ded2ee3287770e61b289a15409e131c30d2afb537b5bc7ddbb4884bf1e24c5a8acb2e32f23e16ad802f98898c3f8b6ffd00d52dcbb605930c591620f76f532f646bb9d1f8d60d62fa91f13a59ec0e7f265857c6a5da6d699c7fe711a33d3f9dfbb0ec8db4a002db044b040bd4ad0309f9acd9624d2d57;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b4145e268ba9f8d0a6f24a644868b3e7467c41ead8cbb5bf4b89cb6fb8409d19575f29e6d62c3fd758f373957ee3916a255efbbbb235f35870396cf600073a747e7becd13e11a8962bd4ffcb061ce0c9bd8a8d28982bcf0e27ed0fb9fac594a77d42ebdeeb9bdcb8aa24ffd62d6e75df3b4a2bd88d72cbd5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c7f31ea4d183366ee3507d9d602f86895427ab2c419fe5f3f12829c4b2df510984e44c0f39aff68406264ea5f81adb62448092e13a08f899d138eec19c7e972e56f3b2831f948200dfc5ac293f5b2d5a8d1dfcef682292aef7b55ff8520ff87af359e5441f9b65caf5c22b6addd32f0038cc56a412b74f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eb553b09371cbe6fe328fc451e724d2effd6c67326f09679b79d1b6c2ccde1520d83351ab1a266f07899a0b529acd355f4442fb5d98790843871cd3e0489f89c22e50e6b24740f60db60dd34fa92d38d0824412d655acf5c5dacc0d624148925680ab9c503b5e3bfbda6f0e2102ff875b4e1eae75e741589;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8f3c372e822d157b38be76e40771511c56dccf27c3d1d1e3c9e35078ee23a34536cd2c798923877b35ccd5f178a490bc52e49fe374f200a1675f36f6862bb29631f404fa643c7f79d3f641e0c9d9cc504269fbe08ebaec4003d9ee773c18b9394fabde560b46f258ac1c7a080669336eea34f7e65698dcb1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1956946d711d614b87a03c972a74bb1647422697e808bfd02e5b584f4abcc66d92a53ac3522ffbff04725678142c40a3e2624652366961408574c595db1da10f0f9d9df44e6473bbaa8ec04cb0712c4a7da1f4f22fc71df164e421dbb08d46abfedcc122f9f0b43d361674d6704874d7545abaa15722e0985;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had5595a6b9a68964bfb4defea60ad17f3b7cf42e7afea5f34554a30ea8038ab603f6fc2aaf79869c95d2782b2413cfcaa53c183a6575031763d5d557c39ccd9bbd119343917f4f37775e145e0abf604d9f402789d468fd8e0e3678cd614b0dfbd42704edb7248fd0be7022c809e6fa67de4bfd243ac768d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b4c2cbc8e2bc814a41d6bdf9fb74a06c554cfc472b0b37659c5da4b9ff3d14faf008b8083ca3158d0443b7f40ee123bd1b4b50dd1b919b3ea3327190c70034257192c55ace00c372f91b88e5cf5fd6252467cc31fca31c5355c6ad3870cebf2033a1cff8e03313cc56474501936dd97612f041a22dfbc39;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1e1348baffded787a1be0f3e9b3aa1993ee2787ac13b87fadd41d76ddbf83e651dc7810728d74801870e836fdc62393a603c9f2eba552cfabb4fcff018be20d27a6ad1f04f1f53a40a5d93c00777c1f7041fd85437c68c889c74dfd4a396994c688be1eaa5bd842b5090509fe0bd36763899ab072eb271;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc9f89a168488f45a01f4c5772bc046a450e69e091d5cfd038c3b5e359a5cb901b11483baddc45c46c6bcf7d58886d4f133cfd21e2f4cea6d79556cd5664fa36e3ec8f4ef74ea162f2aff4ece68212d73bb93db8b2359a7b7bcc5cbadbeec8128eabf75cf510eba144b5a8809a35e7aa8fde59fc91f923b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8fb7c822f844e0352deffe53b0ab70eb81ba017945c18c064dfc10d55848a16102c0ab3a2554bc5eaed4046b6a8cd13e3d909220c3bbd7d3d965891dd8ac12515eb5485793e60d7ac892c042230bdf2ffbf9301ce53bf18532f4c8f645104f8b3f106b88662cc964e028c94d307fb02cc36f55665d607263;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f01e086eaa61ab8af36afdc73144c2e11c7cdbc01b60ff5439818a0d983fa5ad06df1859841095a0bc31c904eec9b6f796146a2a9311d0429a25ba0fb1acc5401449014fad77669667e812c47a622eeede176c4bdd5fb9661b56869993909443cffa9fa9cbe808a954b13ed0ca7afafe463bfc62686adfa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15a98b9171795fcee60d612ad2df83ce2de5d92387472720dd68f69570605d85fc63da223a73d57595d02dfe61c3069622d8a6e936194cd1fe5f27a7b235a30395145c22de6e13fe3af501fc4328cac361dffc86aea2c5f23ea1b37b7f7fdb501ef3c9d2fd9a64fb4e89be1f8db82575e23c76092bcfac423;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fffd3b735c229550064263b9ddb7d7c25fd7810ed1d559e480248a9efd0de8ba8983e8cbc4b3c7e659f64c2eac17a2660a152930cc210971c47cabab52bcb0c68e3e355ece10f6e0dc81a9cfb33aff682e1bfd7238af1221f2a8993a6acd52a1756f192a3f5336fc500b1bccd73985389c1ff260d20204e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h133f45f94ae4aacbedd9cccb0cfbc44fefe6d80abac50db61bfea11ad5cff06469312f30d5fc44bb026a1344546fd3aea48aec18a99c1e0662ab7327ebf23efd82d9197287c5518f0bb65b7ff5736381ca04f2b559a39edae3d3d65954c4f5a727b2ecb56e095ab9e7623ef061198161cdb358d9b62c963a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17a80fcf8c61126974de8da6befd18c9f0c056904f983e247a69399c95de384ba0b027e2a91813dccaaa886dad192f07b516b676da1c978804bc8940816cd0e2d3ef8d2f8498e542ce4dd60a327d7e41d789a79b1c54de3c0c35b8ed93d36883dafd1a2c97d2c3a87ca2451ea4a3469d7f1ced4442a46eb99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17120f76e9bc035d982adb0553dfd2c3ee50284d96ec454a5504831d723f461088d020202b7e489953ef10b5bad7cab0ad558872e2475c4489a65ec15046c694a4cf4c507f74841418e8ab87c0a22f3278ff0deec97bd9b20eea78b7aa7125f897dc4fc01e0845f387696def9f0ddfd57965586e5fee9cc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb2c1a3589a28f77ea8caf93463cef199ada00540d0b339dd16c71a78dd224815019ef18a5ae57e265d243f64044c4d93a8a1131a73848224b00544e9158df124c826954527b161f54c835481388ecff591c8eee178425326e67d37114acf1f3845d7b66672c06e91a22df2e3a73296ddc13dee451ed8f199;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14ba49b738b5568b8c072ef1bab17813ed8f4267cee07903a4d4f093e20ec81f8da32a8045e228aeacdbfad8c670e89fb535388f95db4a1cf92031ca9bc90f81bcc0b9d34852c075d9e9108f1edd7f88ccf4896b11ac8368537132f99e675081e90bbbd0e19a28d01f0b12fc08be755c4b217deb3355e0b93;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eda8b4a00cddf741ccabec4f25db5fc2791401ce4f939295b41828add773ab6f5c2e1d0f28b2d6c1ace41ce788a127f127a16ea94a44643ec05a8a0cf272fb74a6b0c7377b9e29f8e79d52273fed6f3b4e827cb617e63d354e589d5046e8ef4183c784b46ce8db48c780b9bb1f41542fc813e0c4dde7073f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb9c98653c0d488d6a768e4c4ca32587b1a7cb404c570a9bcbfd6872d5dd2ce3d7b3b67ac068a72f012aa8a9d5307f2f10fe8355d4482cbf072717311dc8ee6e008a4fff9cbccb66cfd8bd867a5a4edede126604db86955b7fc9c53ee1e3da3afde68c8f83c58025add406af7f66a76d1bd27b1a68cfb4c31;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13b3c30c43702176cea042a63e90d58e7569cc8a616f272cddf58fbebcbaf5d73e584ebb00ce58a09757bd73f0b6afa9ab0eb55e68aa860d1df9b97e9ded39ab965a3af8fdaa650792fa8d0ef85cb825e3881c4d689a0435dee0363ae23442ffa905cbc5c7c8b671f780c65c5d6191cdc7e55b6b4270a9b99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c1b1954d2da12771d340d439d8d512db8321bb68424f1876f95df87430069e503638a0058302b3158031fb6d8a6433db20790f7cdb910203c9c55fd9d261bc5d813ab2bf7c0f9f0d45abc07e2b9e256eb42cfb6a208c62bbe63513f21e4648e21c6cbf5d6af7134139dc246b84b3f4aadb6cfb3d6d86aab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1165d531f71ec6d9be5a219d7a413168faf507408c7f08935049b948979f0eb9904de6a94c302f64ef65ec739cf1afa65a37a3494c011c2542b92d1dcfa16600f662f621cf476860b82c7e13582b8370e138cd72dc01c5c74724ac078a6bb311d7d8e36c5607264b12ac1a66daf7dd1090fd3811a1bd0a1e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8bab6813292baba5fcbe8afed48ea53b5de14173143d4c2fc521338f7ec16f8c97c12a4f1baf1faf63fc144db9817907d4d42caff4c3b8ffc7010bac9b08110384720dd86d65f6cd9fc10c3f19944e545fd3faad948b759f7901e0ef8d9261375681b040faa042a0fab54c8eac0589493e44324d1d8ac83;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3c09ff238316572520d346caad7b8dd2aa06c7e7a5aa2d3a031d8344ed6a33fa6ca32e48250bde69cb4c66c9febe6415299acbfcb9575d8ab8ffd6091e3340ed565e062c155c073c4abcadbd6907a6ddff3e50301e1f87f45029da3238f2e8b9685b480059e58d42c5fcb337f09727ff2372a99515244bdd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf0c665ea511349a54e50c80de876fc72efb359b57b7d46a0ded4a9f41c932343837473df86c0e24b5b0451f6aea43827a6ccc05f14bc22bf7917f04d1eac67857037eb6d3fc5832c80b69a03d819ba9dd871a7adc4270fbfe928d8f374d1314df365464fb7c97829aa4dd6a4ad93f9fa01d17e5c31c9bb28;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d53a64ea38b6c510d81816dcd1c652e232f6def688bb52fdd0e061a8e2872c0919640183ef7f5cb58ae592783a5b6d4f46190fa46bb3f87e0d88685b212cab648682586bfae9f6ccb9f16c0c9d6eb9d23538e2a859424d682a6969cd9d5bc09b5ca9586a49a7b482facedbc29070143978cb52af9156fe6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc8e9b3f5800d2ebbaa1fc8d05118b4894a905aa626326b6b8001f90e883100def8de0af4ae9c2c8ecefe94ac15efdd47618318407a7aaed813b8c29305f5a5d9010b37fcf188cc886145ae33715ef9ce04516496b8a2bf0d71a17182440abb6ba7ac1ad325fd1ac7bd8e011b372e5b11703b007fc93c77be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha62af974fdd5d45e962577e15f8dcc1b226e6dd3ebeea8314e4a8cd1275f4a58b76fd86e301871d51ca3a296c2683de556a028e87c63059bf8b6a83f4b53fe8480b6b72df77a3e730a120e42df02dcbb2b65787772769e57f74a6c0b6ad6e2efae33d28a3526102134de1beb45f54d18098d5ba527834205;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c5c00d32ae62353a362651337d80df2ca3b38d1e85b2c43528ec8280eb3ca5b5d5ebb4e4956988d5408ef952e42b431f35420682c4d306d6470ff15f2ce025496d8dfc0d489ad90f9369882fc5c794f5643c542849a60b6511154b20658e940b3399eeda5cd1165f4116263ab350a0c7a015f3e16fae5f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b43a4a510f3bee90aab049d25390813095a59483a4074f40aa9bbd6f7d45e9b5d6671ef270d53195d66cc804682942807667113000e0851d7d6408da707a3f32ab64b5e82fdba73eff6d445845d8fc4725c35b66d61baa0257d434b1b2d6d8a820d50d168f803c370bc2a1dd4b950502ec27179f6cb3ef7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9944e73c9bd3af3653269494fbd05371d56818cbc8a7834c526241870dc2e1c23bca6270415e8a65dbb540823ee468826b99e3ab9340ae6d1ae0d728662d89b0229b74f10f9a763a73069ac627291d3adb2b5a2bca813ad3adbceaa1fbd5f9fbabb10758f87e83dce57265ca1921553e98f910cd5e98d145;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33b17cdba36816935b6683a2974d0fc7b564a112ce16d6db03df5c1cfc0800f35109b177c90f07a6a55e44c79ed626a89dc47a39998164002b87584622f69a73e06b535680375136929121b1181c9002a3fa47fe9947226f2ec2ada354d16c258cab6a1490f4117754d14b5f835a2a2a7161640bf5b61da1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f314e595fcea02464ce2670d4c67bf9925c65cdd58b6eb658f74dd6caf78bf74e93c6a00bc9b6d053e06fbe048e9763ef8f65db111a2d550a507fd93a3171db4dbcc5de1432310a9963bb6837678bb896b0ed78a672231abe6cfa6553672a3a820c5bd9a35172cde80d4ea76993446b273dfed3c90c36b7c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46341e941f1aa9ad2864abd714d9e504e43dfacfbaebe6cfc2b1d472ee8cd1559bd455b93a71f315aef09935635683f262627607a22c77866b7454921422ede1cd8cf4c3aa3a8091ae0cd8186141e526efcda69e8d070fa49e840c836f323b8e7bc81249281f562d7ac2df161c9dd1e1e9c81a8566c1506c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb12e351179a0fc9e29c0449f18ab72721a08beb5d9ae045f069ea679c863c73533e022f4d22a33e4268d493f089690f9f9c62363c52491780d9486f981abe39fd4fbff84ba9babad8824610efbbbb17b18e1bae0a687c0d86643f65300582e4ccbe2e894203e2285b86367e0a086c04e7847946c083b3b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d8acf5c2ec1f07f8469fe97de9a971d67a2780152fa7dd7c383d1426fed41f3b74b3e3597dad10e898c26b9e1b316a5d3d80100e332f98db25f7075111a5bd7628c2bafb6b85998e6c09b8f321494787ff131e177b279c131912da7277341a5fa32884b6601e9df988536170b694d4faa3ca0482a7432cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c8ae783a48c09978f065dcdf100f26ede3443577f52f351069e697f07713a5199b2f85affe07363723a13a08cfea046653a82165175c946b618b30153dc0b320bfda174fbe5dc2c2803db8ea2e4dbc94b266017aed79864e492a1c4ee6b4df056abd2e5b43412a16ff5af9946f0ca8b194b36eb55a09059;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37dc4d38fe395ed3383376bb10e2da3422ecbfed46fb3be7567e842337575c0eb0bd9ee92adf26c57d0cbb48998ffb1d958200fb9e6e978d293e3f01ddb0a506d3d60e1dfe62562857a41cae227c7f160952a72d3f73af4e19f94f168ea3d3f08dda769b41cf653b540bea00732831a170e4db04b99820a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1055b46d5f862b8f65b2aa2eef2d28cffad39589b6445a65ffa42953fbf5fb33ece3a24c08c5c315ba943f3307419438c7f4152b279705f8434e2d9bc39931649518c4a563a6e0c0d302539c10e4604a3ae5364494f4ef1f3720767cf9d84d3ace3400dfc4b2fd1b32d9804a0b376b73e543ffae0c160d5ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3aad8817a37b4051e7cd0b5548eb77e8d200fe32839a7c7bad280b03ba4df509912127e0143a555526366e526ecda4ae0096ac9f3a7880faa80cd64dd44362b8e4d2f2096d9d0a91d0fdbe3d38e60360d847ee66f7edc513ddc95c14875b144ce52c7407c06bda8426c28afdfed3e4c2313bc327c2d65c91;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f0faa2ecc5ce05e7581df4ba753d2a7ce9d191bdcf694ecc0a101e6ff2f6b47e49f76dc510216c91f6f5c2e2d368c88242856a698d905e8e3228561aa8ce227c749aa03f0f2b482a6ca85a76eb26161d6e5056468fffa38ba34f50e154b3f4cf0ef4e13dcb078e4b54175597327683d4dd1b07d4c4c8b88a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a855d3d25263221d677a708ee69c2c88d7c65c0bcec53547c96cf583ed4b0068586bd45f5b1519129805ac3c7cae4efe9bf54163a123a0bc55ba096d7bc5131cebf0f693c8d5004f079342f757c1500ff3fc4b20a18ec4052662397bcd215c6649eb2349633f82bd8307fa7a97b57556de4016a93ca304d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h178a8fce4565c1bc56a164955715a7e4c8276b3cc8db49393ad125d86bdaf47822856a734fae44dd1c7b531378db21201732a70365641a1608d327ce5c0c534483bb03c5c930a56b5adbfce249735bfa94b02ddebedbc8736e497b1ea06e36b1e441f5577dbbe17ca4351d42b76c0a47d6e4b7b0187ccfe97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12de21703bd702a4fa770ba37a387956292e5c3fdc2f243e89572d28c72270dce4b6d97eebd53f52a1ad22e7f26552cc1b277e0ec0db72a01c2102e66de80dfde33ee66f90ba153f24e383889456b59f30867529a66a52d298c6ff3fd9948868f8fa6610a91f494663811f800a4d3e93d27ec6e634d0afdc4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c173df6cfe5b7969cde525375dedc8f261aca257b395b422f5cf968569b4d2ddd6a5954fe410667985e8b0dda8125b60c2db783eace0cfb953404200c114c370da8a49b32ecbc1be9d78b0b9a61b2de1aabfcd6ffcf88444badfc37bbe01126d76a347d6d550e3a21dc0c224fead38968570ca5d775db4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1008f6d319515bdfd182fb361e64823360ad6b99e05c5bd5c8069490a4a5558efb80b229dea7a6d73574e5861f171fb5a39814486faa3f5604d7bf4b7dd9f5044a3dbde0120ef8b17d003f6b23b35b26fee2390a5f1c3de597667debf4c882e3d3e129c8da4b7b96845fdbd190f432efedee9122c77e319a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h96390e29cb02f91f0a309b445a884de722f97110bb52a0950c7ed2ab13d159dbe2a8099a14eb19f539362d63da9df2101fe43ac72883a868c51c96a939b6657e1cadd1ca020d48c1627a5fc8f2c71592a89108fc7a444ec16fc21ebd037f0047e46b436772727589d3907bb78ef954fcd6cc16f0a3e9881b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15325a8e15637ae39972d89b265c5acaaba512d35b1d46fbdba98dce46d445478991f672115c03ef834e1215bae62ba749941fd2936545ca5c81e052db82f7386d7a80f67f9c86b9837e77a5de1830aa0eee50e5eb09b2c78420191d88f20c9c7b91d434154f472e2d876a2c1712fad6e4b4443283315b0a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2b26405154bfdd29af119562df2a6812f2c3a2ba4bd62d51e735914a8580f58e132dd36d7a9d1b982851f33733239c9157c2acde50516766a25213ee830a9857bd4ec5d716414da1b1e70b5e66b2b3635b3fe2941cdf9ef672dbe8e79e5d583703cdf6c6ded1cdf60bcc00cffdde76809db84e0e3176f05f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8499c8b066e6ea680dd8ffae329a9948465088c4ab6402182f4197e5032360c7a6f3676537754252f637c611ee111b7e32cc0da2aa0060ec073c0a87edc47823064f470567eeec8f46a4212aea868fa4f371b6ba87d7950eb087d6e2ffd144d536135cc40148cdfccedfd0e120afe8371a8bfece54e1f416;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b6909d3e0f5600b1fbafbbf43188a80b7f742c5f22acb935d7dcf6cb3892d2339036184550ee38e19fe3c515437bc1fd03e5bb06738bba6cd231bdb9e0576dff9a5ac3fbedf2dfe86fa3a20aa777b08bc57326dcaeae6052f388f4e0edb9856be6a4c0d8eaf1cde36a7d8a9be45702d66d82881817f812;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc3dccb742a9886efa32b0f62e5671c7db30828e310c286c888b885fe91bc2f497342eb89454d43a0e2dbb11a157719c3e870aef2d6f836e7a90bee45e1cd95e62e4a495bc8d9d9c49a12902444f0632a1acd524b93fa81eb2e544738981bc69838f89def93ceb6600a8d6d495680f474356d189bef1e803;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3dcfbd1825ffeecd28b10ae12e6c7701ce0724d15581022fa918307d1fca4b66eb5f0f1349b0b792c4f8dd9a20a5a619f37b74798978687ff74927ea969eaba6f9c390589082101f0f4d05ba2c8826d3aaa94a4a9ef311fd108004af6e367cd295b0f313a232665e92112f29e8fc4891703e4b6c912adeba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c30e9ae81ff3025207d0e7859f0df09da637d1722c4f1a97100ff744a398188cfa803db5600928e1dc5ae34a6f44bd01a730a688bfcb14de2ea59bbb29b457d756c83b238e0364e70a7f1c117b975ef1f1ea32a7c0c083b3f4bf9dca855d1473ea9386636e288e3d9f249fec803cb3a73302f96fbc98f1d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186025b0e2ba03c49f3a4481bd33acf1ccb50786a60fbd76bf510784f702892462d74be9b566f1d7725c69685c9ccbacb0e91e4cb5400fd91e06eb5b93a612c830dadeb0aaa9c5b80187161e5b9dc1bf342704f277777e7a2f5321a8d1ad9b64bd8e4ccee4c3b1d8f4d7593c6d026cc1e83b7236e34eff0d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2d6dbe63ddb33d75680592189e0e86d2453877ee1bc97e5b6fe334027e68dace77732eddec885c9038328e66b74482251bd9d1f80504198f9ad5e24cba4bd7df105c6a125897756d9b254bae20758d2ab1094e1d4ffcd9ccd168220a7d296882ab4fbe5f49082a89bcbe4d72ab1684718959cd161e56e3d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a960fe3fc778eaf70e2d8cd35ba6ad25887c684011e5b6aa5f454bd6d13247e708bbe2bf2cf21bbbf941ea7e76a1824a28e0d9c548304478180fc53d29152ceb9ef6508215fc151269d0c22e6b0ee45bc1082ca8470a1298aa5de8d1f5184fa0e03533b4e8a64e44e1168c48fbf4c8e55845b9fbe54e201c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10551631a0589719a38a912d721dace9ad621c9eb2c7469a7e0c061ad952ad826e712bc965e33942d4fda7425ab43922cf74120b9919191867083487b31cee4cf2ae3c4cc9484014433a1a038853b35b749fb3aeb3d7ee335ab30b02e6d9882f7c3d375008ca8398a3519cc858239660dd6d79bbfa72a31f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha8fd69a1db8ab8a1506deb3ee6e32d6fc3458b7ff9aad45e62d700bd029963c556b1311071317a277f4cb7decc38e3f30ae0001c642c2ee4878465991df709e587b4e19ab86250a1f51a23b0227ff51aab4f8836dbbed55ac40249faf33e0f57c101483644cf9c6c857949ba3eeb52eaf57280bff658dc77;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb035baf7d7a56074fe786682b705e07f7d03316ec96e78fb530fe25e5bbe6fe927fab7b4d4f75e822a48a0d7754237b9d3c3537161f697aa3b0a0100efc191ca2238445bb5a58390c14c0eaa5a4f9a97aaef18794765c6f30bfe12059269243cce2bca876157c0c47c68585cdc862b66b0a11a5efe6754ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eb4e543c4bc27a54abd7ef853d2a17530812361b081476d8f9b671f38d42cd67ba273e3a6a7fb3e817a3cfb79ecda3315caa3ef3a17eab5042a5b7a15e69018b48bd6465498c56a270f6c6ea52b2941a48996378be1e25a8628a24d352e0dd6c64920f465d6aab9e386eb4e7365ad483141bd8da11e2cc76;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117c47115faf46c5c2b312195f7e259aeaa9158f516fcdeb3379b68a153d332d737a180a516b236e07af161bd78b719b06f0bfbee229c44eb4f77837d53ef081562e5f384975a3718163c761a2f950e47593d1baf0a272d300389b2c0a12a0fd14e81d61a17662e060b90d0c871793118b22e858774e048a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156ed2da8e6e88c92319c292a7a93f35d63a49c7f412b7c4e55e575491b4434d8cc3481ba560ea8f28aab9ac6c6561106df320329db677f21fdb31d2ff9ac448bcea62da3e262dafbc4f0d0414160cbbeb22cc1b5276e9d6983ef0f425616e6a86c77788c8f6394e2466351d31444679099791c5ce6d04f71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfa81f8b04c39d1a8d3a0eb79b7693c1646afa9c97a680d4e67ca9d29f10fbcb6c15b866bec8cbccb915b664ac1da1c585a3bd79442a5e158847c680a1588c1398037277548910842fabc5c235ecfd9d22634da5d1ac5a3159dd99f4867d09e1bfef174b5c620949b6f80b40860591ae8ddd5b40fc47f92b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3bab6d019c55bb169894fa94d2f3fc72484a8975a05b3f76dda585a047a5ddd90f68b72cb9b8f17c3983c57e138a5c43a9e43396f974a7321c477cd6526f0ad13fe3cf9b55773f665bf518160e7341bc35629c386e122a9a6683140be2fdcdead864c4b1558020402d1ab935a47bc778878e70ec66252727;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h417b58df34250e2fc4ebb3f2022c7db045fa4df656c7a53c0450fde5245dc8ee7028a479ad62ad5d01e7f5fc0bf84b30ccf7ed6a8585281245a529b50e1316e909858dc8f3ef0f68191dbdfbc9e2a82ea4bcf5749a132514e44d7807ad0a1fb860bfc8531d49989ac1bcdbb77af2fabf9b4ea25bb02036a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1845d2c35a0d67d420a2fa9df16ba580ec001a3fbe26d5546221b390c261c4cebfefb10608d839e779b623223c1a40a9dce189ecffaf5d3b34aab4d49ccc1fcc32ea87cf45abed0d27d7093fa45ea23fb42f72a0eb5873dd6e2b3b342f8d8d329ecbb7f62b5f15990cc57207a46654c7f92ae0a65c5cc90d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb4efbc5329f8942ea7ba2ddc7923eea91af68f858b022aa3267a406d7cf18767365c374bf7565c48336dea83b50857f89b74a761ba3b21e12ba806791f4ed09b722338c7c9294d26d8c3098aaeef60e44795922e86227085fe8d8d1ea187bec3db1cf5d7879af1413ed7acdebd7cc3309cdc1e7e57997acf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h43fa3a3532b6932ff87a0a65b1a236c97265f46b1b730ce8337290c61e11a23c1b9994430e730ad9543d2bd5a06faf7b66201c4b537dde98c0039875cfbd14a5d96436bd2c72f1d6c16da76d8cddcc71dcbbfaa776eb0aa3bd5ad573b194a8ef62182ae01739989891f8cee7806b21377ac3a76eb617c846;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1a65c5afa57bbb901b4b537dbd64be78d3e4b56c60f38d54ee354039634f4fe978ce896cc8d93a3383a0865cb49ef82e61f5dc53948fafba887fe0e731d69c5f1deee8b91bd9ec290a18a19a5f0a43dcffff6fc3bfa55ce259cb06a27dc3e080039a1b6e570fe3a5acdc3b99e6545f3188ce56ebbcf790e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118d1e02dfe7f5d4ae455b8da6d66e07df992da567f2267dd82701f64f25bf062b38e66cbebdef160763dc553d3a4c40e3e28e6da1a12a60c6aef661095d22d12527a38e9d2c197a6d484153a0e6873acfb5607193863e409e55a847ca8863971a5cf30a479307faf475b0e184860e048c0dd1b501d4a9321;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h133608a3ab93ff1895c6ef681df8f139cdcf692e1fea56c5cfe981f50d420f9357af08b55963831077847554d58d390afe08b3d7bac5386262e1ce6e1aec96a156970a60d0d67171154502ce67a783b0b6a54a8351a53f995f2d06a11a5afbec2000258e6d6758121055adb69903d570ab8d7682be42ef2ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5dc8a6f7647cdf6c4e52e95656c7ae79c64ec6de0196c80a31810242571c485af0430f04c6131ce778872a8f94ff1b304edf8c30c457753c14b04a798ef7661e8b541064e446dcb4704569bb1abf9629211af58b30ea06303074d1cbd683913e5827e8e1639b6d9504b5f472ba784820dd5c6959f964109d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb7b3e140c7bdfcfc3fe6812c564f985c316497b1dcf83e04d3585cdc89057cbcd8f56deda29f4fae1d2d8007dad24ec52301d2af0b8f77aea09bb784d880cb1b937ab027aad187001f93124d3563dda4e0305e3816f41e768c15cf341a7c2e2e137bd73d5a00c2840d4c634f63ced20300d0ef0c13d575a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2a4a9f7f08ec793ef12e8dc79fb98f3501a33eb6f4f27f24b062ed47dde201865d52970a33ecfe9ee0096cc76601f944858df149af8117ad2ed33b7f6da3be8d61d8216ff5bea8c5255670f01e920620f898e8a8f08ee072b109fc310afe3faf297bedb5c0d9da485dac8894c2e5b19b4fad23d85072aa1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h194d88f2b269a442c4072a2d86177805b921acc7243d884fa3c0837e286a9cd0090e333869c70005274f0454fda21879b4bad0060baa7c0d3a78f32dca750dc680b67797844d640dd3cea90639bca419abe29312c9c785a65390dc9b4601f29f098725b86586ceeb43efa8ce9cbbe6acd0c0df2f3d93abf90;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4ca2e1e51208e843640b25cb7661ea9570d625795e293fe4436a06f54c2311328ac36ec6ee8427afd27bf4190214e67ab4490ff3b40f27d497ed1b971271dea605bcaf52e4acbe7c05261a67e9410811d0aa1d7a9ed87dad4eb22eae7f82218bb32e86ab70f4649fd461e1801465990e33b4247d31ae558;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6945f71a7d78e6c4393b22bce93349e445b7de20535279362275c544fd36faebba10417c94ea7a66b6f58b1aad646f33c4bc5e3ceec1fe8768053cf11fd0bd642d4061893d08d15d7e2f99c399e50ef4f7ae379553157b3f04deefa40fb642b2887d58be4f0760555c46fc97f11de99208c98706761dd2d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cacb62e3c3ca472d77722fe8f6178ba5c1f5980e6ee2da09646eeb53d72a5e5253520b9f75e4407c8040872fcc5377cfd575e1a840733288855e7f5d18433ec8dd5bb03cf31e16cb6bda8fb338835ea5f7c804ce4fdb5fca3b1271b7279a7826125653443424c0a91b4d8f970da8e6f4977319b454677704;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h197ea89b2dbc1d3071e3cab8830f418907fc3bf1f7849aaa0b5c198fb61181659cdfa0e43b9f3af9b796e8287c89cf491e91efc517fd68b1ba0b149420121b8423866c1d5fa39b6d68715a1b1e54b84cea6173fb66543a02e6b7a917c29048c882cc3b430d559e2f2284fdd983870e29e73dd3d718325334f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae5a13f531cf70794d14ddd6a2fe3eb87c699045a0143c56c11d03e33882497dd97040909949da7b36595a6c6b044ea0f49315cc2491294f41c5ce842596bd0400999937ff067cdd1ceff6f0989cdf14ce4fa7aca00436d01aeacf5189d033d5b30c747666a01bbdff8218fa13c4c2b494429c758f8b8754;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a31ef2d02f14796f13d720d23ecf8d04223466f6fbe8d2c98b6aa73784a9c152575024dcce20bfb22fe61845a89a2947a8f4615d0d5c0329e93df14066331b68550c5b32030cce8c25950c840282ac9d8a57b88de94885afd37f0e5b65aa4771000bb5b6ef94e70536c44fc3b0655c81053b1de4ab4668d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec12653dd86161b76553889d4f9677e223a4edd683f44ccf2d27626eaba69ba19febaa2edb8d1eecec67f747efd8f6cc01a3517cd91430b13f6684fe489f8dcc9b07cb4101b62a256375c2b8709de7d79de79607b838fa6124b9133c1fddaba0926d71516ba58d3b95ce1634b4ab656c5157ad59bd636be8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1572d0c6da06c96511a4c5c160024c7adc3bb4aade3c5ba5ba986249d026988704300e596fedaf46a8d0dd6d9b14db9f68d205da5e4007e7c01ad75a8def99653462419ae3078d5fca87ea8ef03c431791b7431d335e9a5cc8e27f153be0bb22a44b4238458dcfca6080f7f7db1dc9c9a0eca1d8eed9028e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb08d6b38f1aef96b636b66c5acbd8849297fb0cff1a8e0fbcb50e90a414c7c3ae2ec071e6ef0a24c6b4adca1014ef912566bda31d1541dd1fee5620511311b54a56f99472f90ad3bd620b5b59c7cbd58d0a7ef9e352aff1fc545bfabfda47e4704eb4ecee08bd76e8f408a7bd626f09a169d2977568fec2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c30550da2946456c889d24f0ce6c5283d2d080f1c5b84642b276b98dcc8691bfe69ea6e08dc4a1a74eb85f61c665d91ea03588bbb489e5f0ffd39937aa35b7d34476f3159cfaae261bfa74959992388cfefb81e576ed510b75a289a2afccbb4e03c47f6de257b3ac62fe08bf278f234fe54c737818b2ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h403143761f09b265cf1ef49b26b3f81ab8d9d540e233608b3de3268ab10156d1e8d23994d874128140bdba34025989441580ae1be406864cdeac93e48e42da56b59910b8fe99db2d028c46d1adc9ec971f2c541ca6ad94d92dbcaf0d60f36427ac948674577199d61b9f2bbff207cf10223f3eed730e5009;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ce5ebf4e833c5f636eed0adc0aa50a1ed5e282e17f5f89e401cdb0a2ad59a825050b0b4a129b15bce5bb934d168f0e0fafc81f4ce0f0d38860db77cbe32ff6141c2dd6b4661c0773fc4dfcb86e1cdd6c27affb0b8f3f44fe9c76926c41abb7fe702cb420a44661e53c1e3952c6f25a9c90ddf043a578ff4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f6302734b26992dd6af74179b2b287cadec9af7a5ca563ba5f1084b1178ea8b53aa019e220553b32edbba3ed3cf75572c43e12e2fe126b6f920cdfe4584051a3fdcc8b9c321791009852133bc74852a67126094105f45b919965e27420a94c7841a7700fa919a41eadd432f40d3f7b51b57e1bf467e3368d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1030919524a5c22e061cec8beb2d92321bc7638ae6678636e1ab224c65f91c693afd4e68665342b04881df9d1f19f95dee6012faa7da56b74f2ae46e00d5f2abb89ead1d4900645724634c0b7646cd3fc23a16ffb719ce896a51dde38aafdad02aa5d11764b23cdfcdf82f39942194ee47240396aabb0dc1b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h418a57b12371698aaed8ef4ff48bd566c42cfc6217579b1f1feb09a21c2b56e4bb87468170e3cdedffc494b8067f3ca4fb10975cfd8018df45aec3f1674588208ec79826956ff7214fa3cd5d92e8705b4b14070d0637c63b3c1a21c7bfea31b11656189a8cb189fd171b9a9f084a33f333d73798e4db6b37;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1212664e045a7d0d3a26c26bccca005cf17a062b17fd2b7887ab07ad49bd8cbadedd7d2c31e582cf7e88723f29ce0b9133d64f854e0aa097e0be27abe2748401d2456beb844732a4a6d3749874efd996aca44b01eeca722f5cd7d97f57c176c9e44ac4d05e6e4e0707b14cb7c1a0a1a18b62a3e5537e187fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70375b1548e8c5947784d7d93766634ca5f5fba6c9bd5af7c0b941662442df91196265ac7f7c8fd47a3b7538a05298d96d8783b301e069f9dc46964f72b2ef8c460e70c6045bf6469a4a3cab92ab037bc649ae3eb02cb1c6f74c337721a22f792ad5967d86009407c5701b67c2e79abd89dea258e6d504e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1999e0bca956b00f3f4393057b63e3fac1a62ebcecc1cad09f455cf46cc42b97e475226bd6f94fa0856384b57ba319340b503056b76d65f5c88e2a2db9e32014532502abaa174a7359c20f45a4bb79e451d726840d99538b66f2044e1fea2f1c6842a1be018cde0fa1e7bce4957c9602e91010c8020240ba3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he2341687590c55f44da3f59cf1a59fc5768dc079dda83d2314a277cdd96e6ef674cd2985d1f50705180dfa407a795f7a47a9341d06e398c470e371ea18c8d80365aa0335a6ea40ef868acb2141dea6254c10ba34185ed894f3786dc18885967b5efa32e9d49aefdc5bfe9bf4d92581e30716d6df17378340;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he3dab8d8082ff706cccdabe2ca553d4ad8e082496815d88bc5f3daf3bfb1401b2e622b09624f81c8fd56af05f1cc763668a3045106d58d29256b9cd98d17c97ded6b1d048b20fff3ad1ae70fb209b116938081c8ee81dae92675e3ee9e7af6cfdd06e185ce458929cffcf767713860b290ff29ec98b4f062;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha7740f0b13dc7b196b7314cdd7f98d8b9366dc9f643855b7a5f6a45beea6f41dd202d2e385b4f7c0f5586d351998a4f8b08da3b15676ab67cfbe938ac51bec2ed1eed786dc4d5d18ad98c736f62635416c2a5969ae3ade4dd5dbe304e774357960c6f9855d19e1fed6a69c72791faad02d6608348357c488;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h327ef1338078e35e3ab7e2e0ff3524c72efb57d94905ea766adf31a6ad4ac8b774b1aec27876fe5e69d6e4672cd48da4da6f3b2e5c4716199259c7cacb1ea112ed60ce4b05d761c140876430bc3f44869f380810c3d6df0725e57bf84ea9f5757c827cb8c6a3bf3e44393b4569324dc06176705b50f36b44;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb6cfef3e14567417947110a95982f36eb88530ee90e9d0b9bd9544ad2adad5386fcec28c648b70c0bb5f5c242d256b3954135be2729259b262e0c280a4bef3bf22d56f93c0017079f5fabdfe4076de53254e70c1bf9915d3aa23f60510aa2f7aa24ad530c8ddfca7af909f0103e43767af87c1837211f5a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h81dd6535c81a3f73d3c2e64e1c42db979ce12a39fd609e58a6168d836b23887231c1c900a1db52624fa01842d570237f0e1d6294b607ec92cc195c4eb175824f43d0026ac70d378f841419f4e9712c6e9c9a2a3203fd5a7d2c150c5c6f01a3265fb1c3a9a696a155ae76f84b87fbb3b2915f0bd3b9bf2abb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hefba7c7c1919dd336c081ea0567237d9d99cd26901d8367876294246693b8119e754da6f33f95410819f87ffc2e71ab6aaa364bdf2709c9dc42602843e5badd442033ae642270000e571256ab4cb773e60832b5c8302b0ef15ff5296520d2cbb34d12ce4140bbea744de826c9c5101b69c88717f9f63913d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb67a03a738fc403c7ed66bc2e91a904b2766e3a79a4b843e9caa495bd1aff1d8d875db4c692b6f6c158d8d46ca3d7c24baa8dbeda47201f8ef03d5388a1d43ce0852c93aec4c2839b13d2f93252200e274aa0ce38ff881ba316302f07a3b30801295fee1187638cd59edda644ffb019fdddb90db219f2c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h811797803d116c43d4e5a604d629d06e7a3298bedc5e1b737af5a654fee5cbd84935d4572f1d360c356406944204a8a19df403b9d1527d7aa20411f996ba1718699c62d2a03b2d946f4d54eab635246b97385e04dd4039eaaa058e8150162e70a8899f091ec215f8425697fa0c30cb81cfa8c95165e075cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd27bc3a89199941d8f9c5e4f0bdbb6c62d12c92ae17f8f091deff1072eabe10bde6c387abc2b6adb56f3748d2152340becec42fb29257fd473fed53fb2093174aaaa2312a4e0436f81cdc30244631f281caf7c29b022e0e5b80eb915d37db25be6e05e1fa6fdf2bc728f23be0c9950efb8e8d82f4328cbf2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb175a75d49650d96156e40e82de7a53fec802f6bc775f8274150897c2a4b0512ca490cbe6ffe56cf0f1fba0f95cb2cab1428b000647ca150385186b0b2ed5b89c2cb9b66a351068c1629ed4979b4db6e61d92cbccc14770b38397d5fc734166fcf8aadedd2cef8b913312444c3b5568e23e2c569c78b2206;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137eee51315997b12b9b766054127e29de849d17f1df529f31e702bf18283b61ec23e1614a685d96070f5dcd743831102e5fdb7378b4469a8517f751c80afcc6d2eb93bfecf6bbe1091cb3e928136cfa7125061bafbe3a14f97d7affb2f31fa0e0bc8fa74bb31a1e8c19f409812f29e663f59e3eb15ed1662;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4fba26d0d7da6c414e0c9aa4c06cf05a84824fe2c9cf87c7e89ae9849bf88c53f77972421a68d64cd65794a3e2902092e7a09a8511e275622203211aa08d1c215ce99436bfd9df72f231a5895ccea3157a31aa40aaa9b9ef0300f4233f3326e96127fec2b2b7729d23546fdd9b67e6b92422752e194aa823;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h203d4b167144532897630415fa6defae62c7dfa92a9a96d3a82a201bd86825ad24e8e2aa7b5ee0fd2323b4509fa8b2b899a3ba08fe4ffafe48159b2b92fbb2fd0f4a36794f4690ea81a44dec2a593494eead2bc64b35eb08d489f456f9fb5129ffbbe4e2822b04421fa25f08c734746a0847c73e1c38dcd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d38751c520436ccf9322fecdbb25ff099003a2ee1a1bd058df54b3d785fd56c6a588c5d238cce3e6ee6f1cd2c40128ad9d804672c1c099da4e408b1a8ca98b28bca3f7df9813b3c975db0ed7b113f38417208f6419448e044c7ceeffe1680ca7947404fe3e10fa940586ae78a78c001c469accb60e86d86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h230564897b6b0f193c732b7520c074a259a1b8149078d72eca394c3e49917bee52eed183d161c25fffcffe067b2cfa1b1641acd9f349abf5dc6f3fdb7e9f28ceecdf2e9f7a7a825f533b2ab954193ccaa3a6a02fb4ebb6e5457c4ab89c2f07e63e86dc32a110053b57da4a31af743f387c2a29a782c68ab0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he3f6c3c1951514b4269075820615c870ab4b2fe80b5dbd71f67b7e347cd312fb92d8ad1a64afeea38a460e6ef5149f4bfa3706250d260568e2584f6cd15b575c9a976785c9cf4ffa524b859aace1b0be4487720cdf815b75e812b35aebee0cd74123cc7a85a1331561d9589678d693d96b59a65890bd81b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5603808569d86fe3ad1d777fb5fa537775df3e37e5fb93c45a22f792cf3dd3bad9370eceb0d63b5a28430868f65812e8e5a0ae769fcef721fed499b2cbd2dba501f55311cf253f11d7ef63fcc1c4bcf000208bef7e08eab00c867f405fbd8ae3a66504c68463b2831ef3ee5c2b63718e9c102d64c41f5913;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e38ac78578993612f88f5a104d33d7921cd859ac4913c9a3a50f818e652af67d72d73e764b82b20279879c3b64d67bc47b83a3d4f435904aeb3fed91b872da65acf30bfce2a5cbbaccae5aea968bbab4f56e30e946a0aa37bfddd565b580751f2afce91592f5afe3bd333838e7e9a7cb24878d420a9a0224;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1623db6f97ad9c9efaa464611eda3ffcc40bd287b74dc41afb7ad8049afd0da60add336d214cc2dff75d6c4b39a628faac3a0b886fcb2330e970164754fabebe40fb90ef9be29adac57297befc447b9b5510dd748425e78ee5dd94d4357cc1838ff795badc18b0f879a5cc1d91ac703b758dbb359baec53f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h171e610e483a3f1615d05e0279e11ff43fd32f0dd1ebd79f8639f19790f0b1cce1474f59baa373341e18f2b0e833314df5f488a64f3b3533a32905892a456b8f33f27e32f2f1a429411be0c7f5e6d94fa403b179e5f599f76f0726c04e0e0213ca090ef67b67f48c425d7ed3e6668d9d01cb849cc9974989f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5f7568ed475c2cf240cfedfdcdf8c7e903c0738f8bfd84dca221e494f16b3d9c7f3578a888c3e27a67e95c7825f31be007abc43a7f3d6fa0ae40beb120aacc5f4299b1769b1ff56054d083121dd5db42a41b8731c0490dfc3b6fd59c3052c15ba31cad68b556229bcb325389fefb083a157d9a906373018a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h760721561208f8a3b06cc205ba6b229dda235da76dd7b2b20fd35581fb22e4e8a1e470a5378e5f5a4f7ea0b6a2c0302145bde5183443ceac358a83b9f7cc7f60e59e0ea42802a22415f4ba5c355313c7072df70932fa739cb5e098f8570516dc5a955225300b6dafb36f7c5ef111c010441f1154aef42406;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1249208d60153f420e5ddb7edcf48b90bfd627ab4153f5860a67c9defde2f70cd72a6f6e63e0050c0d25f4a7856ef8c03a707cf0df9ba7e2340d43a394d37c1e2cd2e34efbb177556044585d6a1ed68323094aa2a07de98ef030b8c207644b614a3af8b5abe85e94cb0488aeb27ac43afff736905a5272f37;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e779f36cb5aa4f632f2ae73d1c734a132369d31bcbcda1d2e8a968049de54e76cbead959e3633bd5ff7760cf4fccae09163f2505502ab52179fb660c7fd5c867408341b24eb405f987cdc99ba56b460945b022ca6f360faba254bc7b4fd612f41196fa51335514b4824f9195579416b60229fa0ee41aeaf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1832152a8b850c6df6e3377acbc05c9f7f4a07f6991a70ee6f2b498315e36e89fb95540d9a035ca9557693ded8a061395165a4317ba88528b92f847e466c3bb9bfa11f4507932ae1ca69ad41cf2446f6b8973af56369afc4ea9fc6c68d731f9e92c41a41834d10a0cedda888bc9d726a5e3fcb8e3489d0f90;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1995d31013f0c44f582063bfe677ca8e22a553aed20b2febe09317c87ef979fb9986bf0754ec2c206878f911bb0cd2b9ceed02d11db1b8aeead8d1d9b74d1f30533b4c1d7271bb2991f9a40b5a5ab4b4145c510f1bddea134dd493c46ec719944f27326eb032c71c1f22cf0e973afe6ab91b658cb8069185d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h109a133e3e6e631ef37fecf6049cb7c16b53a4103d9cbaebf70e94df29b2a8138cea952ca370724afd9ad5ab38d3846535965bbf5d0f7c8d551c868123f3ccae109c6f77f187030979cccb2bec7aa372aa5f637cc786600d54d3c8e9b98597f18ac9ceac37a50d5496742d9ba685a75cf0061e5662806e236;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h834615ad6611cc366aeaed9ee9195d9deed9e6745e128e9b986bac0d2cca87bc13c32b852a7c88fca32b2d5e999cd0fe5b81a5c223ce4ff73b82b0d2d47ef3e9e1193d6b3a7c7cc85aa6b84917ebde09a2d529689ac3acc734e788815c15d50571da90f1a4e6cc7bc1587a2570ccd7a80a2152a1b1be173;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4342aade284bcf6a394107c5012e2f3db04867082707167b71b0eda0808bb594b00353f41d79b14879149bcca0ab5d12ba17e82f26be005ce00687d1d6dbda8491aeeb58308005e020478634c55d06095b7c1ab45fd406448ba8321b21f6a1d14fa184ac64f857ebc17ac67376cfe84b4bf8521d2562f3b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1394b9640175df4b937c991bca0bea401741c3030e1aa8f98dd1c079b87dabf16284826c1d1cfa04a5bfbd51572c3b568e6bb03c9b52940e122bfb7b875e2b93364226c9ad999fea7859f64d8c753f0d6c68787ef9196902d03a32e4e3838a0cbbede6cad379e5057a1d0b853450e58b353d8f416ef1dcaa7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9e65eff0e3f2e69b9fd1b94e9221db2a1133cc8866e8088aea1a34e31ac3df279624d70641462c552d7790400156277c53fe23e3896af5c2b6d7990d206055004c0e2f68d6a3647beab816cc870712da5deaa52f7c92036576cbf5aaad89a4b634b046d349a8bc35e8cc158a8faa882050cbb360fa2a4061;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1c9826386c5f975c09e0588130c262c895c5ae95134eeb44a2b25208f57b9a68d7a2156ad58982882784a9dc688d96e0c4fd19631df467c15cc5ce6d59561682ed491ab564bb03d8fec8ab20f3c0990c76dabc2fb5f5fe5124f30f775df42da37c702af426a71a21b62e7e7b3b2001446c180a77718e01;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12432ccf2c397ad3e2a6a176db90af0ccd9a7c636fba67e1753cf473724989415283a8002dc959dbe9b2668b517f643c80b5344975eeae3b9d648ab0828694c8ba384a8e2dca9415e0db308fd69443c3ba7b0d88ada9ce81267f907b73b9ba1646a6d540829f8da60d5542c23a041919c082c1d3709caec79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h152c589d84bf9f3c9015082d5e04ba0b4262b20f388c51612c79ec68fe110ea73f8ee2e298f81f7df9e7104970c338f359c708c2bec90e28e6eaf1bc974d657da8b9e16c87176a4906567a89192a544d93eada559f0fffe7ef7e3966355fd3ff6a2afdd47dca393dff3d1c25e1e80133402e89a842c928559;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h891c5d4e2dbee383d78ebd7f59389e6ec154702fd071f27276ec574d5576a1139a709e4deccfa3ac752333fd71bbd09a6c3b176e7e3ec1b4e158b921d387ad31bc4b656c0f954cc056285d0e607c6deeb54dc416b315eff5e2bf5929ab6d755600154413d6aeff70f05f41cb11f3831ffacd66459ec8c597;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h97053030bbda5aedc8223fb69e2c430d6668b9dc4eacfe57b682563d7aed1f8bfa18b3e9b176a3ebd729a842b53d56badb0dffb1a1745160795a5bc25d8fbb37afa57b2528556a99d7cbc884aaad0426bede77c95ea721f3bd31d2b64338d22ac536af6ea33ae5f3ed7be044fd9d08a3a66d55888d24158;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1db82974f826e8ee9687eed339163745443f7b4ffb4696c78f2f4255b3db8748de726eef3ae52c9ec8734ffd870d9b741a5cfc42442492949a2ecaf51b15a623bc2f12e7f10fe709d11b4cdfac24ae995fd592cc67cdbc532b82bec48302869f7f28a45111fd8c599833f89879447749c8f897cec9236d788;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h238dff6f5d78f6245990141bdb984937d59a32dc85e128df1868c552cfb80303688891238d6efcd1d5bd28e1d2dcdea2736e1b0a5aec40da249e6d9205da9d8f7f48a9a5959fbc26302d0d96af2e46e77024cf0df43668fc32a128f9ba662a56257317950da1a1c9fcb6b0a2706700b037442637581d9376;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3deaf43e79942dd8c43f7e6b0a663d6785a9a53f6109ed94f16fda58967b24652d2e372b757b164bcaae031fb20e9f5f93ca05470d9305291ea87400a470dcfdc61e9210b75987a42cdff84285c69aace40a4cf04d035efb1d37070404ac72e819d8fd835b52d235e841b0c741fd7812c46162be21a8143f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ea814c148028f81ce31b56c064ba545d43e7356145b4e312def445ea659578690b073f629aaa8c0a8fdc0278f7892dbaf66444e3956ae8cb167c020df307f37c5dd00375221732b444feb4d016b22f57331fae27078610837f7994b5e9f34c742d85c9d971b8fa979b4afebcacee0f3284e841328b3233b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hca893bb1bdd613ed318565d43182520696a6772cf54dce9a0041896e179ecd50653217bfccc1ba0224f9e0cd8334f8e9c41340821d366d4aa9229e5b4eb801d52c55f696bdda230d28fd53056d6a0aab41c7e4d456bd5fd8d22b452e4fef7e3433262a78c6410a1660d1f3d0c82c7421956cd14556db8a08;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d37b695dc6c050ad640ece424ca946c71e7f17cbce16a17c1c74be7fb0d2c3ecff58f5ff8116e3147880bfc7ac9f4dabc4aab63b3d6f1c748f1eb9a7fb50a0c7c36d2e21804704434fd0d72e93fb6f16c001aa31d111eac90c0e560274603748f97e961bb0b7379a6f19e81637d68e5f408d5eac534abe7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1adf329515dac407f8924a7c2b19206f54b2ad70134f6de491d130a2cf714f96603492b32fa84615db12eb1f2e1c733b1a9b628a584e853268317c148deeab616f34616aacf2844e2add9aa3a7eedea3429c0507a3218ba9b68a1e5465579c822774c9c61322018b1552bac91ab469d76291abcdf43f03358;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hff10aea0492e716a5ef64f659a8b419851235548e271fef76a4243485cce35513045fc2401a7ee453c4325e53298ad140f9584e1f6abacf54b6fbe8eca2e860e673b1f383a856c1b9ad809614b38af539211e69af3b8aec718d5815ac1b18435e6b5c347b5d041a86f81bca82523319a474c363aaefcfade;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f04953fd9615d3fd6eff24b7ea52dcaab8ed8bf7578f07f70d77157caa9c26c7425d39a89fd0f053c0be80c49bfc1ffbfc6c36cc49dde7fefb9ae74d3c5fe44e0f8fe7b783618f6c9a945e5f382bdd2de7d808fafc9816890c0a06ee56801d431263aa00d28c61801dd7132a9b7596077a2f08fcd2d747e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcee9193e0f42014465702ffc26a1f72e108b6c162e91c785160cdafaea6cbd9b325ae687e4ef58977a021b76238e89bab150d1b396cfc988f4a7ba8b6f28ee957abf05aaaa75b35e43df297fd40b3ea5d907cd09b982cb63e45e1bdf8835fa667a5a6a10305bd20c48601c2f65ed2ebc792ccf5097b1e992;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14b65c0fa5890c3a9f3b9aa286ab9eb4a5ecbc33f3ac0ee5a0607e5e7f41706aed1fa9710292daee59c3d8b601d611739d05ea9b7f901a75affcaf59d8fb922bee7b882e45634f709b826add20478293920d9433902a5190aeef173060bab0bc47be70c15fb40404d0aecded8169b206b11ca7532806c01e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h130cac5e27f408bc49911e66dba17d97b2930724b74ad7fa0349bbec311eb6b5ae2b86adf9aed7da4f27e5c037bf29b29f5d321de316e4f0edafa003c1fce9e3f8b141a89971d00a3c18fc0878c09709d6e793f8785362800526262ad42a8cce55ad477268f3166c61c9b686fd57e03a6bae0231cd3cb1ecb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc82ea61fd1362febae0e61946f386e7c3b9aa385d950a711aed9f74c252084b5050eab9765bc2613b46ffc756e4ab6a152b6c1fe6e60c93a04c847385de3be2abb1a2351ae003bd016eb54eb4b27b089b3a1d40fb1e0b171017c8e5bf82b68cf880b8e87c8644ee80d53bb91ffc7aafd2114d5f1d490557d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h25ba890d45e47a80ced90c698a7fff43c0b64335499b3d6801dd36a860e69dd8819e8c7a1d6b2edf2a55d6ebee5fba1952eed92fe80f772baab664e1cb88a77faf05405b2cc60602c2b5a86f9e4626e79a0c4d913ecd716decbb4c4df24ceb7a9d929bb6900a5dc02ab2686729e098f01f9e6a0a87122885;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f0171beb3f66b0d20a20d987d8d47ad86c0ac3a046d12f3bc8ebbf38a5df6ffbe0ae6a4a54d08c70ec9b6ce26bc1fd74b138905ebd1fb521dbc9dedaae1871dab5808417797d18bad8b5dcdcbedff191366dd2d90dc2d8897e61c83cea54965bcf172b11c46949c054610f0fe31efd1468b26639ef32f9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9507549cc3d4959ff6317530c72cea29575c3a66f7d2137f387ce7d7d2fcc6e9b9f2c4bc776ac3d5c35436a58f085dd48d3b515321227a0303db8b73bba7bbfa62d91e9ed56fdece647fd754007dfdd6d6444a47c53c9c01c8848274d5a0f02fdb29e4a329614e5cb1162c81bf4583fedfb261e7fb08062a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82d7e7e48498e2232fd70d360a9c428d8b15f8b71ebfb1aafb9f056ef7daed033beb7b0cdadf49b92119414d1969389eae418e439d131ad37c0e7cfa146dcdbfcdf2ba682980d0f9292c93525fd9ff568bad29630f66538fd6d21946424bec5b28451e774594f072ae98df367627675514d03c17111671a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e779342c15168de6fd6b1896f7f639cb039ad8319be063bc76ac0ea3843f6260c5c3ff85d4662e3dbc493952f1d87494cb881049d96b4a639807194803d9bb2741f23730fff9f125794d5bbe0dbb2798726301830671569a8b47341e24e2b9487bbcc1741ae50a9c4affd45f2a6c079e07ed65bb4b4bc78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18055e6844c9e1837bf9784f3ea12856b4f0096986d8f3a065045d0e4a2214833b3b0076a1c1381a723fc61d7f9fcdd28132edf984805f925a4f34ee5e111db12a5c90ee1f6f7cffdf168622fc312ccead77c7afd78e59198f2c4a5452bd6f0e70fead727bcf9871f938f6c4f9f2769c0fefc3545766f75d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9d3472b317a6172428ef2893bc43e1fcea11556569d7afb9b74dae19ea0dacd7e6ae92524c435416900cdee9c4ecc315008d76388e70abe0a65f9afbc3d519323a9e7443568e1fdb9aad7c5dc05a69c384869e2d93c44a63d349c0e13de85a913e1d2951b66261b5cde222fc362ba968155c3b19e7a41c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb902b988f0246e9eae2b4009af3b05a5848f9413fa79723b832c7009d6e34513aac0520c322ac319b5bb2972bc720152acbcddfb9f8737ea9335ac8ab356e44f4fe9fe30178907d38e6eddb0a5897de2a480675bf5ef649d07320970da12c368d0150e89239aa67789a220c120b340e65cd831c500c8f4b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1320efd5cab76981c8298fa79cd644b2944fe6e9723be6e2c8247307b4092633e0534716354f96ce8655755c03df69fb3076c8c1f8367fb921f376f3fa7797c31e55f1da3be1ec259efd1c4e8a93de68e42f510dc779d6ac02107f14a9e5ca2ec76709e1099f741e6c23a1f7ee63d7d386502a8bebeff7e03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha29569d63b09f3f42e04d6633ce4ea465458e6ed9504c203bfe9141767ea5b634526d65a6ea3e0b78bef7dfb77437e321e367187bb74814ce107d10775a06eb6a1a81a7f97decba9ca443d081eb7ff2cb4a535f8c64eb703904a3c4739dbd67f61cfeda8bcbb0ed038396ae74b367029f95d9b4da6aa986f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h191c92a7f69488b9268bdb17f7ea94bb60984c2cd77a539b3d5c56a36f693704e9853767e73b70716b33375ba45a7bf02c4c831ce930645db98bb008679a8121b00afa90d38379d8eddd9322a8970ee36681b049c55eb207e11210beff6f1b95406040b90a8a2a301cae9afcc8484c4ccf245ae73e0c3a3e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18cd4302afc44b50c4ce33a0b561884437bc5db579e75b8f86cf9fa1b9a9c2125c7096d951d22fedb0003b2ed8d272ee03806592a78f2d0825d65b2e7349494cc55485daf7a29a697caaff00909325af5a6ba0955e8061510ceaefc91aed589c2f57ce80031c0841121f34f17b586b80145d388bfcccb93fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb37d6e4acba7ddab895e5235379c6d189da30720d80bd27b5c2edc7985dd3904870aabe84bc93eb5365dd34f448bb65756b4071d19730e2d56c5834ee8f64302ed4b5ac2c3bda000883c05dd1410af5e74d402cd2c9ef196bbbd79975b114cd7f863fa4d9162d132601e13bc09989ea947b8525ffcdcfc59;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88b690a31ce2b3f65a042c554c5f2b8f2157ef9d40317b2e855dcce8cf48b72cd8270b0bae2fcf58fb63b256a65542853c54fb03ec378ddd700554c439d09464305e694b9ee0c952fe43d702c562051cc9fad068eabe7fe19537ae30d1a90da302aacf4b16d628c27ab2dd9a16a6b87c7afc6c40b5012513;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1125c702f4a00a7f65384a72715c05dae9224ed8789763905541b566bae6bc1d104dbc65fef8b18e30b78f94bf661c3a09e44ed7db29ca5602b9b2009e1a8fd240ac23f00307ff6a81daac32d7598a1ded4e1a49caee8f9a0d5ac4075c15469e10d56227aed35ce5f80c7d0cf396cee218d6e529ead51bb8a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb5e4f44858b3a6795cf4ee3f352d81981093961503ff9a54d81900cc2c5f4381334c2047a435f40861c68a7335c112308536905aaca8a857328f5fcfae471eba61ecc32be62d5e99fa331b361215c33b6399936b7f2e0fa051b21b3cec452a01be4a7756633e09e87320526e38d2b3ef4f546199275833c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h78762d3d03a1e64492eda40e92623173779953c5e9f4b39c57bc5353352d0f417997e636cfcf77c62a4ef5f13611ef0bf900e8c1e1819daa191862bcb1f1a170f96aefc95d87c5a0cc91c123acc9c872ce9db52acdb293f1a93b60c53e68d820087aaa03ba387dc114cb724cbbe8fd53b33d190cbf57e743;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e578ab32591befc9bff7bff0a844e570199cb171fe3eb5bed6a04e508bdb0e1299a43763b3c0b28174d187ebf559c48dce427539718bcfeacacc276bf3083c6bdd5682d716847d9b1193c6dcafce7aa9eebdfba33d37558b664a236e23e147489819e7e091d945096e5f2d0de64a13aecac0cb51099724e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6b5b754eaa187468b9b13dded77e6f6f69b583dd278c9e3b4d7070ccc6d2a0915a5590dee800f8fe8561239d062f4214053b1beec4a451a5118d7f78bd02e410dfe04c697543fa394ff581cde67b25941c6c3bcabdeb9c3cd5357c1eba5789b2fb9a57070d8b4dbdd38061cef582981250eb57df47382d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70fb6e8f1e6da21e04cf82a9d29458b5afef0399025604072c523b8d95952c40f02f7cee6b88dfd2d6d10b114d16e2d1bf2999376d4463edcc411b9ca1c68449f9898f5074bd1eba0f1928d69e856e5a58355ed24c6773e154a18107f0708d0db50d417c96f44a878e804fee7f89b348ea1eeec600f4d7f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h983f726fd98a5ec27243796e80f56452a78d66d014700445089ec9d7ef2f4672d750f7349a54010e6765f5f1ab090d3b255ee9cd2e7501057e1146badb7f4151a8bc85d8f362c75f77ed6c047a7fa71f471a96794d66bcb23e5ff0f30ba3a01c9251eea79f9619304c66cbc34e7aa3b9c77a3ff386b3b66e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h958c69411aa06738e0ed3b59dede0f8a2a7c84e76776bd447107d2ad7e6c4d47bfa4aecbde616ac7cec8ab746684f7992176a76ce6e0d77175c0719e01da83ea06449f7160461f52926d04b00b6dacb4da337e266ab92bd64df420491bb65d225cb461dc7277084b6ec00785ed39e6db74edf0b10b7599a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11a86df243576e7e16d6fb893f45cc7ac5c4ca20465ce078c220b336d27b515d9dc3b5adee5a50c27a458f193476e8013d9cada0d0bfbda0c0c799255689e86e9a2156f7dd08d7f89049a7df910049337c431e613f0c85c4d3d22881995f0b61e6cff7d66a7c74adefcc8840f8b73050d03873e637e90bb62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc2cfc5eabfb50cdb36ebd067d0326a3644a2f5b74597013197e042b8f08f248d87db44c047097c1e1fba9217592612bbce7288e615efa3a248326d15effb62498b44a13d89c35a679eae2f97ec5698a5a562bd4b584c44deee39017556ab67503e82e280d99f9efb7acb1122045a8a1a56c977086c2625a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1ab7f2616bd944cc000e17c8dac42e6945dacac0e4c224bb7f9aa6c57b6068fa9b9628dc813612b27531a525d92fa9d1e448baa061ec213b92b7ed64d0849bfa3a6d7587ef402855e8989770dd273caa18f2fa3afe6ad10cb3f7a86d033408c067707195b570399107f2fccdc5cc96124bcacce7fa56892;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e6faf62c3725e89f4ae5047a0ae5dec0774f91bd3a997d2e41763b058e239574b04cb8241f9380de7c8dbf3e0a9ae9875b4f401c31b4ed6dd6803babf3e719595a1c3d54cb56ceaa6d786c70d38a21542fe4e44bc8e4793624c7c8a84972acd7f7966b3a2fa6d8fff585dc5c4f26d2e18c36400d7915741a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha49a919cb80c7ed0492fdad33440dfd9a245879301c4886ea3bd0472fdbcaf822fe922c2108bd0861bf1ce11584a0f13b79f8ac286ea34d69460cd59f4a1d56f411a60aaab832f6600092d1c0366ebe6f06af4e82710928ccd76a5b19993b9523cc6bde2eb9cd9070ff64a1a86a1dd95e36c80d04f44bd0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee222dfa694415211e9acf3cf85547a359652f1ff26d6a1f5991e95f86d56413627ec90282ba3199a074ba743098ab7b77ebaf4a35e08c69519ed689133cbd7de6c69338f7b1dfd1b63c698c693dfd2aa6011d30e440479ae6c5c512eaf6147dc2478db206347ca4d6e95abbd8c5b05999ae4c71efa53e1c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1efb436961e8dc96e20e6a33d627677b976fd6192de213a82cf27de0cf38330fb8a1751ad25930f1c9a3cc8de85450fa89cf463a9b8041fb119414818a07f9c22e56df284ea927c107349fc8b37ff31b6620aef9840e77bace9e752011fc222451e962f015fb951a149627552a5a71d5050ef038797125d31;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd2a045a670d86c576cc3e891b594de1a13eb55056285924f79cb98f3d7b228eec59f95960fcb5170ef17881ccb93df13e66c53b17079ca831646bd0e469cbd132b5ea24acc04ce83a0daf8446417ee9e1d81b29f666ffd04be33438322a119fdf809cc0218fe22cf41397d6d65465c1f554359cdf44c5f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f78186dd8276f26962c65803d2ca8133c151884cc22963e543a4748f5a4ee09880c5fdebbde827af4ce3ae90c1d8425d55466e89c648a7913947d3e7e0a6ec6464956bc6bdfefb44afeb79f78349c7c4b8f4dc2d70837907e11431990cb34ead872112f5d4093fe4faa24f4d01b8d55b5b0a457ad8b38ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ac135d7a3e88f3c374432ce5c6e86edd748dc3a3ef868a42db2e92646319525126d7e3e3bfa7261d856b72ce365ca9a383b5f8801f598b2fcbb4fcafd35af12abcbb7b91f33e367209feacd98ccda715c93ab5fc132780e6b00cd547ffe32dddc29873fd2282f222946c0992a937fa8f24a6080d3636021f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1874ed09e982032e96b96cc9dcaea84478ce1cdbe0e3e20d7a6b4b400e5e9d23c3f21e7d864bff003df05efc150f5ea8f4c7aa790446203c29d5604085bad8f46ec905fbe725da1446440d1609b17ac74ed774471eb35f74b8b7a28e722a1d4efdd20ee51ef2e7c586f516be88fd77d81286d5f43597beb9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b2917fa59c21e476d12ae2808eb502a27baf09987cb854bd9ffa05dd8412d575f0cb2f6fc788af50ac097845455e705e9f7587f8646af95149d2650b997f95732580db7352cb321f2c0f7f8b4108c1831e1f224a02f7c71de826f0e1b78bafd413a45dc25c9635cbeebc496f4d4a381e30020f2bf9068b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f056584ef041e7a91d6ec5cfaaa6eb02d3fb1ca952b226883174d2ba7c8f345d20f9a63474865f991d64f5c6b16c67df2c75b35ddb8c4adc0eeda9b04a095e6c1350d42f772d621ee3adb9802f66e829586e283368c69f830514cf86e7684a5f43053a6d44e4d7cef9deb347fe6944449b4da993c0cb655;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1440511ee6a5942039baf79db4f51ff18b987648d73590a49ac64e32a6333cd883611b574b3f5c1626e657438fc1a1a91ec529d59f734b97540a9a1afbe3a0c7eac0dae0f4138670dca1e2ab2f7e35ff2f6c4524fbec177c3099355e4ac128ff7fac80b60d83dbe13795fbbeb25971cf1f67de106194d5f31;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b6449912e9ecf6b94b513bd2186e29e99f29801ba0db4da5d934132b66a7a29e026e4bb376c47a0403dc24d5cab82055e256fbe048a761ca7f790190f6f71a61f7ec2e87b5194c7a558dcae8ddd19def580d321c64d90d318000e83471839b39759654e426f5641e5d85c01c34e2169dc988370264ebc3cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b18bb14081cf4077c39bf4b9aa2dcba2055a87a05e74a0cbc2328bceed7555bcffd5817b636aa7a487d6ad637030af650f0508e889f319943dae7d8e7cf240125f01579acc70d883e5e34febd1bf160564a253358923ccd610d924ee8d4b6f941f9f8bde66de6ebb0b2bf1475bb11d6eb2006047849fbc69;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18745cadc05a60f2179bd5dff5303c44846e9d988f64f591a8a1a668a829085e9201703784868cf0c5a4b4e7a4638a3b088a3d48be6a18ecbaedbc299a758f526d7fb70fbe1b0b2e9344d13bd18e46a9b6804516d5f508c0245b162d6c59e26aed89b4bb7545b16345f0f390fd15af22deeef546fabddde7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef553d732c8a5e35524f05b03a6af55d6d990c8bd952cf56f90ef9b8d297ed20dc13700de33ed835ca9972921ae1f34fd18c17cc430f031a6939bb29e199b6201872c03df70d5edfa1765429c880707e669724ab0709ad3adff252822bad1b5519830fafae22b3e6e4394bf4020cb99c3823cf4278ac766c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17100e26bbe3a5c375084fba859871be392f8205ad2996de1ead72095f4dbac4318be2f8c3f547c9f1422470850f3782fcb74ba31bf4a795637cd5c86b4249b773c32baab9617e7807a43233224b06a82782508caa9c86822e90eb28bc29d2ddbbd035d7184851e996e91154216a3f791d33b9a41e6dcc84d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haca0e3249e1c3d0af2504b5ce7a59389acc66236bf6090e721130bb9a22492c6de3cabc96e84612489e357fb374f8d06d46460aa2995456d8095ed03c95d5374e09fa9352979cda75821a9eec8b8cc303dbef1820860ddb77f6faced64e416accea5566e94355721e8e2286ba6ef8fc2f864e402ecca6eb8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc308dc96667180ad58ea4c3d33f5f6360e6bb74b8b36f769fc9d00d27c39176a63593ec41f6ce9b97d7123dd2a447bdbc727742f9c0b0a9690389b24e625de9dea02476b4d50026fb307d11e7688d778309afbbc8cee23796f16cf5f80305a98fc6fb8ad0260c60eedc4d8e674cd3aa88ee82b3419ebd85;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1837d141c1c220101c593c392b3ae71514e1b208cb8b0583edd25409b9660532a313df49630714364dd9736a5e932b4847e9eb95042f4732f9903ab6a7e32970c15b5cb2b9c89625c573e34d1beabc8cffac6638d13bb9948b63dc40fe18195d5fc8873f625c8cb4f38c781183fd801277492f42b7086c346;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h399d21bb7a823e3a56f975c1a198b0854601e5870d2ce0a482ba03c8b0a1df0b30f848f9ad2d8fc680df423ab6554b6f9bbbfc7fcc6fb52277efa8d7cf58425b0f724ee2119b819dcb35f4fec9a7b89777bb0042d30c8ae73d49163990c659c6984faccf5b03e069eb4e60af3dfd1f310622913c8a517d9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16adf4d8fade53af6d53ad93295463ff30d8c85e54c6e41aa7a340936f396b9fdee284f5dd30050ee1445aac25c1d13bc25b8b9c87bab7ed1c9a2f0e16e3a54aef6393d69303bad625940eebaa197ecc8e1b5cf9c9e7cb9e7e37cecdb64de0f04ba7059e59f9ae2e0d5646d59b7901e391ea68ffde476bbbc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1191e56680393f0818b22f1e25781def438ede4ec7c3a4908de97310d9b171b50f8ab548383202100a93c8799359dd6b57e382ff7b2b2b2569748c9cb651d07a5a22f42a162317583fd8ad45d7e22f0fba413dfbd8953ae6aa6d41f037f3a450d7dc9bfa247f43a1865e19ff86ce66ecea8347320a38630fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5dbddcdc0cdf044a0262766b264e0da85d396a33edf837c9dc5f0dd6cf403bf1e019925d103ee6ebf81d21dbab976bed22a15d709d80a9026f3c8396a53e212f8c44e0cf3c23cbf79a59574e876ac803ecd5bb3551e65b9bd732b864bafc8281625d51871a3c58db07b45d181fdfd5a508b80aec3aad8e02;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h120b67f0488afc3519e7581ddbeab499c4dacd69faced80b739719951bcd5fcfadad8250bf953ba8d69ba6fca5410ca73c74fe95971fc1c3dcfec3470cc9b491cf3f055efac8c122d215f5c2017e71c75fcf13c7ddf03c0ed4c9f23046fbd75c25313f1395c1d28bb3d66b082e2ce65c5e27bf34053dccadd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2754f6b12e27d8b089589274a0f2e9c9cb93256fe030e2eee88a4f21c6f5e1e02c2c0edbcd20eede8524a782773a4b9bbb1287f12a7959d7bfeeb529ad2efbad1a910b1d4281ff484f1576b63734d4f8c41c55b630c5ba38858059f3882b79923ca80675fbd571865fc25b7b00a4350d751b775bec89254e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h131339fab984d04938b08319d5a8ca69a66ee8904e1aa7c4ecb0f54fb34c36a1d070201f5dc6166815a630e3f4aab4cc0ba4d983b10cd802d7894a58a100e8cd41146c5af011c81181d4bd8a97aacbb33ad53b4c49300ef1d29ba8dedcb8514a6083f3f7bfcd0f26c47ed18af5483aef36bcbc6c29e959c8c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd29fbdbe062998979724837b46e16da1eaf1b3c5b1f1a510b4050c25b65d5c05cb34fcaafd8b60a6c09e2f6b2e8c4a3c1a2ac234a14790a68f95998a70b0e0469317cf56aa7044af922dcc2959ec93cbcd840235a53fbecc053a794ba10445975b5df45666c5c6bba25ddd32dedffd9220f90749a242b8a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156b9f6cef73dd76fa3ff6f01122eadf238236ece24043886f22169a358a20eadaa87f00e2bded407a74115bab924fce513b417dbba17b6a2d33a3bc5c85a51cc38bfe3235779f18ea74ec455d77f91339b668c930d0f5873289d4db3dc46a85382d1261ef8ba04fcd55314b668fcf95132608e32d6f75ba0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfd8ef0c78f0ea10e5cceeb919ccb3a5230da12b1f4fe846e57ab1609a0a30845592ab19cf027b31b187fb1161d897198b17fc892d66107e2444ed9bd61352f43f1764da0bff490809f6c8a55d32353df7cfe7ca4d5ce4fa383aed7a6b23a8bf0e2e57579457c7690f425c99a8fc6dd62fa095e90c89eeeb8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb92df80b4bb861665448db2ad6e268153bd59f273c3872cc60f59759f5259239f686954706ca0b491f9f8567856903efacc408e0ccebe014034ba2bfaf001290b703008c6ca959f85abb77bf3848543ee5fcc6c4258901b4d8c7dbd1a466f534c46b00020448de9250a5b1585264cbcba8a17270850b1e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9cbf769562443aae79421d280e3d2a53927bf38c8dd02258f94628e8214f05d112bb50a3a283335a7ebb81bc9ada68403eb8419884a7052238c0d6536afc8ad01c99e8d8379dab6d6b4793b402a8d6c837172a419960a77a49243d0328c6a40a431944b3882e66cc820d8070548ac523e8a2da0fa509d401;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h452958e3350d3f44b97017e9f973d8665c8116e8c6223a0f3a80460133b8cbd5d3ce401cd7e0602118e1df8fb41af133c069c07f6e1cec190f8ad20ffc981dab5fac3d707161082aa22e61be0ae05a7ee2784b18e86f576a43f8c55161cc5d8139f8c0150fe0cf575b6b4272ca2a0f579d396409c130e265;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5aa06e09e2f83713b9f58524f50567f063ba825dd2ec3c566c77656b204e74a62023a48612af5030a9b6ceb9a7a645cb2b0f52018f2546e4cce4d2bf70361a093b987601ef01a5a84cc687fa7550ceaa8f3102fa8389230a9ea3226bd08595aca8a2abb163054ce6ad52d2c7ad941843b873e2078170eec8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f8f43e180700f82baeb8f49ce47ff03ac0bd9ab37bf3473c1ff4641bde149b763cc1609c09e38ce66a43345c290b6893ffdc6b2bd970aaeee5ab990674d593ccc23a261afb8dfc23f0ce3c68bd89ea7d66f25f1f5925d7e9c3f571c23b3ff63c17b5e0503bf5b4e9e6af95e3931f38f188cfb6ddf2fcf2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1baa110cea4e5dc91757ff39fd57e3bc3d0558743dcf88f65cf22fb0d99526c4ec3cc1dad2c71049e93d54e7dfb4eba3550c5c98345099feda00ca0bac0ea9aa6813414c0051e56bfe9aee437ef65a3e98a0eed92aab222963c3d0817f924666e5014cd6b6cbd25a3639865e3aca74ed24cf557da901e2abd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbd073fccfaeca9c3027e4cef58cb6147748f0369be74a88d90676a1ab66d4f6936cf86a6b5004f3eb31fbda069b40a3a8ac44381555ab8896cebe9e457d2ad8a722935b18fb92841bef1ce5c4d880aa3327ffc0cc64fdd613569cc8f903b23e33c6d08c43a60c3084c63f006019d1ee89a94662a5a22000e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18a9a13e2663b0ebefd339ad8d80e4e9560dd14b4e925bb65187b27ceefbb7c397da19d7ebad64fa91e44adf303d9c127e0316919e23d62a87eb25e33a3b1ff7332de59c563101b015f63afdb341932ef1d852f1e465b8f2d6ebfe38ae82d286187628da076f831134309807cb2c5162f86349b285e212821;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17d6988829466fbc2fce8ecc5746c8aa03357686b35fbba37ef9237913f1cc496b55cc0498c1a757fc918a1fbf62b8c24b355fa0f0aa802029c48830f8e80cf29c9a4c8ad9c6a1a27e5264eb72af3b91fb87d49546f8b1955307aa2809b9a0c020e6332ebc3bae8843fa91bb025abf4a1c429d08348e63643;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h22fed6dd5e6d6a792817f683a4595d5b8ca90dbdec2bdd87a54fde8abceaaf7a8dcaa79dfdc7bc262413382c80f6283823d47adc09f161d1da8cffecbb343f8c8781ec26c65262b1b9cbe5fc01340b891dbd80c5b688378db0fd769225df816c8025378e45e18d1c61e231722385de4adcc3df705699d263;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1a90c33702cdec95d486a41dd46a38fa4aa75acc879930904380d4799b346ded02f8ba8b3f273f430510be362ef8a1cdfd52e19433302402a25511cb61227ac0c78f1bf598847a3a77a88dcada790dd721d2e50d550e72a9893eaa846ef470556954c0010bac4fa8a5a66a747ee3a2709ba79da20059573;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8ff7b326bada5c6c5031a3b5d9dcefe3517d567ec5f24bc29cea6f7a8edacc29019014c5e42925cbe9e1818a6f8b3976aa96e336b0b80d11c39c1ca9dc81d16926233c05dbf4ae0c6ff0c178307db14494bcc6c79552cb88c6383460e7d5882473312d3c18d8869f02a03e031877a08b7d35cb304d18084;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5cd74ec5081fd53f35574b5a23fc1c71952e16ef2771921dd82e5df8463f1ffa9224b3013cfa6aef4c560f49fba41bd1f8ff32924266a407ae25487281850383cdb7ffa681facd323846397801ca71f492ead557b28bae5efcc84f636d52309129b1ee310050d5e743859b0cc9ffa15de558fcd5685aa72e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf67a4e38bc6b296dfb803a3ab3d79cc2e2b550227ad0e35bc7db6dda7441def294e46fe3f4ca1a677511210c0e63c0a52501c7cea2cf8ef797a87e32828e6f9b0bbf52a12c3bfdc94fd144fd97b46abe6af0333039d24bae03f64ac08f3233158ee755e65262cd844de648062d77d02761655922c44a14e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da0bc19f5d2ae7fa6c649a470dcf44fed567725982b247a254cc08c7f683a7b03220acff9f103c65b9a930331767fc2ddc70d90e154ab844452c3e0a9eb32fe79e8161a99579ace7ff4c9568d8e8e2573dd3e35e111d925b3f2632b7dd7cc1f8df198b59ca09f2834250560d856da62212ad253f71970b51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde33bb83ccff34f475b7bd098ad859fd42409c9b35d8722f5bc09a7d98ea750632809d02abfecf800ce5035ae78f4315feb602a268e553f6616b908de1569a6539fc1791e41a3aa3b57a1e63487908c5a68bdab8fb131fda7ed9d27df2035990e4ccbce0063b61ea52714d1e2fb7795d94ecbe21ad3aceba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18fbd9f9a54f253c22992fa76a819e8d71102394f5c2c7be8dfa8b04c7caab7d11ddb8190554cd53f18e2e27945314c53b4bb2a8982efba944ddab3f4837103831bd6c025e91759be8b9ae50a74ef36d9ae337ede05ac4777e1a4e246dfd35290abeb0cff9e191286f73969f1f1bcd437773a7c180b2a5dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11521b4431ef686300d4361f14940cd3b753a193115355f28771ace7a240eeb07f4f22e3bc97213a4457095194f10ef4c70b9dab86f0779988023e94301929c16f0e7b9cec938112d650a6db451afdb58274da48c61d7121d8d3d2838c7a9ec9172676117f9e553db254f4cda8f58efacef8d4590f18117e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee84ae9ef2c3828661fc046b8feee4083f6ea5f3eb00bc75db97c4872ef05291153b5ffe450ad47b3885cfd4073882b5773b8d1937ff6c3b58b1ea611eb096a3baf91cc5c174c9380bb207affad28d96b5d25018c54f33e7e379b4c06270626106ffffe73914282412ebc631ca978c25fdeae19bfe191fc0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h198cdf13f1e183e3c01624669d22efc0d6f3d53826c5da15f05f53cee13c38d6bba3bd221b2d1db923d9d8e2bb90add33a5e7b38380dc44e14e1cdd7847fa4a527c90a75e3092b8911052c3eb891f1cbb33d28d910d47c4c08c37f8fb9119b59ac500197afa54150ab3b39b067cbc0a652d06e6e0d5eb8635;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113f0695747e52febe30231f11020efce7a7fed07e07d7872cede3c5ed0435d5de098b9825f08edc3d65c59cd2be8cb58dd06bebecb4eb8dc4e4ad9522a2b609243372d5471705a722c3910e54c7851a947ec99636fdda72332b08b44f61e93bbf607f36d2f3ad71f752b2563f4ecb87a0830a41b35254e31;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf34495855e2514c5e3f616984d08edf2a237f23093cfacfc8c700fddb0a36228ff944218905f18664e7836c4afefaf9365daf7a3452e36b3182f6b4e977b409fd4ca7ab9f6a8cbc72da46be44369587dfc20d99d6620f7497274193e287e4a6b9c55f505c830c4bf97b673fb5bbc82570295e30f9c1c1fc1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d521121a6c010a84a1af93af55a99fe83b3e40109e28b4076a63bd6066d90e07c82b6b70d6503ba62a4b83b90362dbec6c0bf6a9b623332a2092cd91e14b1d663bc8d46bd63da6699a67350ff6102c79a76a41cac96d71e0bcebd61aa1a0613b111e5224e6baee2fdd451dec7a99121634c294ceb6fbf1a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1007de5d7fae781628957333abe1f72305012638d800d621e063a45509c401fb76d5e398a4973fe409d528e410768a3282fbe89bc984a2c63613436551ed0e391d2ec5cd41b8210254960cfd58fecf7e3fcd1db0ce3c807e5714e00be5553c178e60e8f89af83150428e45f8e5b3a10f8119f3d7924703643;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c0d915bc32c71c616313cffaf7faee93a9e4c0512c812d4478f7fc1f8c1289ac78a5a4dc2de753fa7e2e02236afcd0ce204273a138d8cc903f89b7b2399d309a81947d39fae055a2c7f2f651a5f962c89d0da86642f8fbd239c6ab8bdc02b89c59f306c050cdba25fadbb7eb38af5cbd171e9db4b2aa272;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h957c8b88764de907ea21a8ea6e74a36c370e9ded0a32d05c33424b0723f918d7e630c00340769bebf4d5ce8fb9fd24123b85cb384aa473eb6001d92340107149b2529c6d34b6c9786349c82f0845c7229af569b6e4e4d49118c663e337d1c4b94ddc96c4882451c539fde53673eb6fee453e4ef372c1477;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he1c9923cb044dea010170b0186be208555d1ad24fbab91d9f61704fde62af1951b9e39d894f30f88c8bf5fbc35b9bb15874a13a89419f50d99f2d22951e39261294e87da04b2873e60bb7ce1253021c09df94c7ed1b1a8020f78e8123faff040aaf6a9dccfa42a22a9e568feb53283728f49cf3731f03c96;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc843d3eda2b48a368ef2b3764ff41862169be5724539656f38258330afc0d8b1c2ea3589cf1446ff250b53ecabd22f34a80a27ec2c7bb512c6596fe77a08392a1d4da999f91723bdfc07a80bf2aa23e8e94047243bba30abdcff3d2a4589aca1b6e951d7a413dad1ac58957a2821fd0031b932e84c628c9a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h92c15907ef850f31a51d71213f7779e091e886477116753b3018733cf5e39936bcd567af301b6a34bcbdf1e38dc5d420333391569763c8dd36c645d56ee87d5ba36a8c60792461b86311423dda9d2d00f2a44b6d898c847a2d603dcc4c3f04f76c2a2d292b0b047cc8b509a84ace9c928f434b6ffc36cf2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190bc419ce02dd94a8fc761dd788f53a97daab35607703ce681db70174e7f5e4da52bad8f8244bf607d4ef8669f929df18c93dd7e6b1eeb111724045780490f41cb8bac634c6a24a16e82c4a7e089fa9ef8c00e71d485db2938d4c82cc53bfc0f72ee6841b35df4d3093320741762404a55abac0a2798f01f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc1104b4c3b643eaa8435654e9dc357bbf9efa1aaf1182cab486a65e76fe37e367b444d5eb8ac0703bda544eb2469eac826a98a9e275b57fee3051af74343f008ae9531e25cdd2bac5291f2922056b1e166f4f4ae30c2923d162859228fe476baea218c27537275a4c128154c00edb210227a957546f2b46;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h139d2e6ea8e74af481da7cbf4630c3760b58d7094a67d9e194d6c44efb2a5b7dba2f11fbc7a21a58f9b88bd178887427da82947cc9e95e8e37b4a32d33da82e5233e08c38470db4b7bf67e8644f3af4de87463adef556ab69376ef6c287a31577b610f48128528d78c1aba838301a2c48787112807552ed80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he3606dda03f073c41d5c7fd18b94901f2faaaee8b57adc41d62c22a3591b83336bc3c406ba66427cca7fc5a0c1f0158a55952babd469bb36254770ce4de7ff9081a5b02e1445a19acdf5dd8a663a49642b4caf54d89c547568c477488c2e0a4698d1330be97f174d96a90e3265be51b503dd265d2460caaf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3b4b7374c42790c864288ebbb2b923c32ea1f5e87c5e97024ddf769cd98f631d310f6323c7605e338254f70ac96b5680c9caac3c2237611c486072675eccd7978a31e399649da9304d7cfb5158298e235f1720c816e9d8286feb8ba2d9dc78e06fc9169796780c3e80854a1fe893d2a39c24d5773b7ad420;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2d0f3857e5fea35216082ca14a59db9e1cefee90b262452681dc8575588e487d608462b608dc37384d82d857ec458cf93e73fb5c3dabf29e284ca6d70457a7558a94296903ad271bdf2c33a5d3e9f8d1416dabe52efa97db1c165ad00b72c516533b6e5a35c39e6b93867c0dffa6e810dff4657a83fb0932;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58f6ac78ae71fb3d227d6debe24fdbf94814e90c5e98d0c60beb16a2cce9b66450bd65b41c506a1dde4eeb7279cb82ad53aa36890b3343bb44c1c13e42ca37e2b5f63a05714c16ba811d2d58cab6a270801120ee70221b3fe1025465fad9ed1fa2441fcd2c43e367bf0dc4d9103ba4d2d0b3333850f77841;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5aeb7a3be72246ab53fb6c30833885e1ffafcf40b654a6cbcd121842710f3044849d67dc6ce7367589c9cdcaa8026d67b39d929fc23f3123dba76602ab8afda8f4bd506c787356f6494e1851fe90b55a0191cff864ad6c6c566d8512db8461da9a908d67d31c177b672be0fd8ed69a9ad21fec90b538dae8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha54a80bea6b2807272bdd03f573b45d7e7d3bf88ce9df7c05b176a114a1f0c41ba729c4109f852452b0719bdb3cf270e030ffb3cdfe6c2d9178136be389d83f0266986db32a634242f2a3b2678a15f23ac1c2709d7cb2201d77319e600e4278dfa6dfcd00f9fa4ae139507174fff6074436085def8b1dd1a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc5e32bdc77260f416a546aebc55ee0502187df4f8ed6d7c79ad22274a44e3d200363758d269ea79eeccce3fbf35a8be7aeef71bef401f4e01302b1c82ce9ed0ef2d3ceb97e43972c9d5c020ecab1199c93be0b9e185f2858b159587e16e1ab09ca102f8b2864b40d7bb31a8f0847c44e3080f00f8483d5c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0c9b0438e05aeaa8bbfcb977749baa127fdff998407d870ce87ad4c19ef3064564d8bed760f1326fa110567140bde9623a366b3cf0a0f94b5a789a10bf1c2b40306d6f3ab8903ae8a4e17f9b8c84a63634f531e0c353f3ded70599047a42e3774425f249d8053a6bea5ec92e22268e58590417c655c03b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2160ff852ff68b4879435b6f017d11c619aa5ac4b1be9f0128940aebf3cf10723f4bafc0b1daa25a24c1c3c46645695831f3596e52f60c239c54b7ee4dc61531fac02dcaee7262773aa4d071b293640a272f5723824c4b18155bfb8123c7ca113cd9bdb050d9b97ec0cb5f4d3795dbeac73f1b59ae6de881;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9e344760513d8eeb8243966db307bf8a8c49e1cf953f388a3704871446966f9be93f9b7462f69059c3c76fbb39b2b6764b6d34586c17d91d23f0fd0c69d5b9dc286ac369bcdc2d697dab6594738d34f4575b13d94705313df7089d011e6be9b1910ea620f7ce8e61fe143e35bad3c3ea7a41b9b03c9218f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a7b8725a815093c9ccadc6b769953ad122fe8954fe2af9d07a6f4813472e58cfea18d0b5dbbda23603a9c5f99881a925e1bd5f1f3463bef5ce4b8c7d725f058af69197ed7fce10dbbb4f3765c4be3f2bcd9281042c758387a130017b4d78a01c9febf3fef1dbca4fb985c874af3f07c514b88ee32d26e242;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1920169aa710a583363fbd7fa6e556d140ba835c7df4feb2a41a052ab069a1edc2f4cbd21e5d5abea066ae1ca600b826f8563dc6de3151e3dd327ba7ae4cdcf0fd977644f9ddb2689c6a141d736ed54bc15cfc8e1a2b6a78bbb1a3ff617dc2276a67cd36c9d00af45dc87a74dd72703bb87a290cd4ce1e146;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11eba0f5f674815246406ddd3ebe5edb2afc3ae4ce0b6cb70833eb88564c329ab259242751df7b08a3da148d1fefd859f45eee9158777f99621772c3431c71377a86e7b0cf47fc5049a3a168cf4be86cfba8fb33c3781d0cced690cb82d103c9237fa406d4f8e2cc401cee4e331472b68fdb52d2235e2af34;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44efdd6b78bb333c9fbdf36fb1baade3c9b8ab581363d22f2e68da8faa35ac887a5630fbe9d56d7a989008b4ca54a08b47ee139fffb854ea9ec2cfa30b61920d8b4cc817007e47ed71d3e417000d8e55484e449e8eb80ae74d0690e1b1b254bb51fe8fa4ecefd8c1ba820148f36dadf9c8c8bd6e5f15e0b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h188ea57025e81041f80b86b25fbca8f15c160f620fa4fbd61f50e67e82de95fce6dc7a61a56dde8b5fb48c2b731ef50fb1ecaba6597744e6fbde5a3e7c404048d4ef512984a5ac916f824e4e94480de440132f090b4dd7b99a4db9675812cde257a11267d86dc68e9647d4c138260f9ba3ee5d4914afcba38;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf374865c42641e6df782dbc9fa8bad36e56ae4ceb7b23d963d8749d6096777f0eb1ceed2e6beb9f3e3a8fd5bd0dcb9da125cf6d031e6e07a2893c6e4973f560292731cc1b21f6822bb3f9241128b2295f69396f70fd14353617df20b52c8da5f87cc8c86ede7b28e94005a82ef0fdfe01bec1dbaa6f4da4d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h120e689dcec72429eacbebcff6541daea8067af9a92c9ea372bb87486fb12fe122f020ccd36aa3786268e189783935b3a6212b138aa21bae6c8bd819e5aa6b38d0d8b94bd16bc077bd13a50469998c59d0de4b3bcefa4160d561fc78a9f4450dfb68a05ea36d4c0994c4afd953bdb62373c082e0dee4729fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115ac82e56f5c25d2106665b54b6117046015de241cf244c83950c9c219fb68901c89b0350a3a7f18e462212d566b9357f7a3e42f2b2ac7861643ab42ac4b9bca021d4f6f53c966d96c1e94a5ab62a8389c54f83aecbacc513ec02891f9a379559beb6f8c49f7566f3b266ad7c719f0671db478b724843490;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181b85b0c9c8fd9986ae5ae59c5f831220248fa2ae20d51ce7c87babbabbbeef8545a6a1841f59e370a6efad18511898c23fa8e7e99d3765b030b76e5bb54727c358c13e12002f15a1e950623576fb82dcfc075cecaf7a4c5605b79210d179ffe3ca42814af8cc07a2410242b0317d203a48cde8799f6de58;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d96a1b1569db5faadc024785607f9e58026460506bc488207b251d7c97ad61f0b33c7c6998a931b947725024188f864dd2cfdae8eebfbf4889b678f8ca7c4f154234590f8bb62d40cd1d3b889bb182a96fcf701adf2e8fae98e1a962a5f59415c48c1ce6d883c1e41c8281a25b0e5b4c626cc9c2fa9ae38;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa9837c155e4bd93c5c06f693f32c4b1a048227a878ef784d484853150a9183474cc7b7a1c3af7dd89ff562a2026564b1068a69e0f18bed99c2e863b19c26cb2ef155921438279964690f4860647e8ed1c7ed76a73fbce2b3703666da0131eb52f7b34c38ff19a070c3e13a8920b719f3f3a4acf7a2155c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132ef7ac7063920dc05922a9f038afc0f475f3971fab9e98f4e2545a7aadfe9fd56a06e7cbce3eb4b437db5c5eb70d373fa043af7aa5b156b4474501dc7752579fa8c42b747a78748909380a419857f482e18cae987ba2804f241543526884631525403260c7920f86fd008ccbbbe7beddef93910b3da9798;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he220aea96f7f14746b78fd3aafd28e2d712a53572d83abf3ab34b213c5813a8c4742561602e40ca04eb85691bcb72e67c00fe1c8a3c85cf3a39aa7c7e83637ceaa3529503d0e60789796436626dba56fcbd3e974068963ed183c75c9811efb53b5b9786a1a03ee967fb2d01f3f7093ec41df191052168539;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a35e1ccee8f5a8f4df08118919ce1ba18acd1f0083cacf77436cebd7100bc85af75cfd6d00c498939703d39b72db4bdb942ff4497f3c5fdbdc5e9c24d1ea8e75f5af51b8d096d51e279755adc31a6041aab83f701074129687343872c87f261ab9c241389f05b1cc744cd5f523ea25e14fa54e614e812948;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142c851923793a2993413976433d31e2fb963f12edac36ba887b81febddef4ada865eff1c87808ec0c3f55585f39546ef8ffc47d2d316596c86dc1eab5d5c1554c07af8549d7ed0afedf007d7184afc3865376250576d35b180a7acf4cabeb97674fb6162d3aea8da179a3ef791e22bde93591e0800b62aab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa4c7d77221c506918cfa805b9fe84414c237cc798e6eabbc906ede5ec83a47b1744d95252b7603df6bd8f30547190f2799120abed9555b81d6afe43b79c935d8bf504a9dda8eaf39983acb58dccf21471e71c1674e290055e9fa327fb20215a1766a0feb77f44f265756b695acbf9d21d679913053295ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8019c8239364d9d2558b974d2e479445cf078c7fd1d381f8af3b22db2bbcb8850cd6f7f1d1d4f7817d46b5fb0a37b77fc655a6da33b6191bdc0faa7ca0ab861f3802182cae86b86c16b85082058f36ea05a9f19e000ee57714acb87422f6587597999e148107b9fc6c30447e32e1ffb55303b2760e49a109;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h815eb67c063d3f3810f6aaa0eff77a4ecd0ede1da3d6484eb7b6f5c9267cbeb843512e75b88e5f841aa2ab1146e9bd19738820cc0ed7c2e8c7d0bafe9f453010959c8c736d9500a1668c8419cacbba7924adfdcb9241f1afc5b1463205a608a0e055caba05192b15412599758c5d35ea1c8ab678b1127bc7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ea5f638f53b52e12dcf4055023ea4a0ea1d20fa5df24c13a0a01b2c085e2bd868096b71515b1d298ddc77c16c59167df281538fb51c1891cfe1e98fc9f61dc7c8dbc732b0c5070c63238c6a726e665ed85fddbc17e628a7cf2b0279c89172374a9592a725fe80e123d21bc15f7a3314e39323856f05cf77;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc5f8b3fef9cc65ec5f62523dffb96f5e4fca48d88ec381966f47b4dee3cca03d676d8fcb90361c0991d729655405a54f03401715aa16041c71aa25eb6b978c2ed40f98ae4fd402f0dbd28e4ee7c769fb6669bb6f038426c53ccd1fed23c8f440e78a3c0c6576af3614446444f9809b7decdb46ba4c52da04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h462ff9f5dfaa1ac86bc32a0a705f4de51b5d155718604e7688c53a3f44cc1bf04b3429a4987410f199eb03955f65762662857233475fa3496c35de311e13d4e0bf0fe5c656b2b5b63a73b77a9faa37d9d20b91b0abbddf130bda072751a5ab7de74f7d8fe1d96658c8edd1f5ff1c88859d7e2f1e6cf886dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h94f102acbe29908046fac75a744b2ea4b42e2f1d84486412511da02cad70b23e04d31f709f8c4fe8cde4ec53d872c3191c04c5b1ee4fd6b6206a2e71268bbeae3d8994661d223d6f3ea4cc93095a7b3772b0f67dc7f6bebf00945278ffae0b4c6c46ff55317bb20af2882fd0c7c81daec9617b58f4dc56bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa61ae49d6b5b259f400e7999d34e32fba1af19914c20900ebe4df60f6680b985390e102599d88958e272eda65fb169e8ee4cc4373dc153ae32a11c5546e45e093f922e76ddaaca47133bab92d23a4e91a62fdfbe3ecc97edb2b95ff179929bd707b71de880df60743e7e15a3abdf80a473946110b0d4c80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1701dface39926b95076a386c425787d44ee9ada1878146b09e460c6c53887c9b6cc8b287862144f6add50260ea5ba20129a09889915f8a07f8ce7d218fb08d7b1612c265cb80da149cbc403b491e7be3a80eeb3e3187081ae070eed82a8534e947f03a4e9c9eb1e708d866ba856a9c46726bd6ced06eb306;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b18a481afcf49d0b85d7c040b526d92873a01f8aa432700c1e07ab0577b94fa2a2bb8f12fd55f5c5e41f0f0a56df2a8f5c4e6f08f8c9532fdf1c5469c0f2b82ac5cdddc595eb91eddad1f83b702de4b0c07aec9241b494fc40ef3edabf098b69a6e88e6b3d7186317fb526582ca910a4ef2b6172cb59878c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d711c3ce937f07eeee8885b90b92c995b4ce14f90553805317f438fd783c24038ce84af95375bccbcbe78d8b1fc2dddcf9b4b8d47a92751ec20e2f8263ea75555f06362317e0ea3337ec50147b101e0ce90f143aeb3d53cd91a55b3473fab76bf32f2e63ed614848efca6943576b44a0057fc1c655019012;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115627552f5721a40667aedace2cae9118e4e229d8b61d90983260a553dd02ff72c401adcfeb5feed1833c9d7e9b0593eca05c9527b105d83427e3dcf03bdd5d653f42e0cd37eb2a5fdaca8a73abef175c842a5d93e5c804dac8e390e3739b58e27e3ff0e5fadcaafeb1ad7dc99583a8f8f7b9f04dd61c324;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e7a63fd690e7f2ec855ab0f156871cfea5aae5bf47a246ae4d8d951906695187796c3641595aa8bf4933421d8be4b032312dd430372df34b2371c94498adb31d070f553359d7eec9d703a8467c64a879cc4c0d42c1387ba5348c98026a9a68665de91db416a6fea98e057fbb3868e9e6643bebec43e2326;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h191d999ecc09d973712fecd7e6d4e34db2e7600fb427f11afbabb1c8905e2307de6f470815ccb366797cc57dbdd5421f368f6810e85df20255e93dddbac73307976f57f631e339fb988497a85a06b4adb3cebc040b5ecd978c4bd859bef4c40fb78958eba17b639e2c51a6ab342b007a03c403d2a580afe39;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf495504ac4855ad1c74f6da10c2ef546b5dc4b70bda891e6bd0b80c6a032f84b7d51224c9055ad70ee70db32d97c643452480406e09747f1bf8f13ed5d6bf0e9c4eea91507de6b48bb0dea7dc9392cb23b26f5c70e7f18a329d27ac36d035992369cf15b74495930310eaa0eefaf99cfcb0bac752be0f62e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e30756536ea217fefa60d50b7cc174ffc5a3e9abdd0ad1d5dbad915cf4f855269fb85216a4118a514f10b82f5f305ed8067f5ca39361d310d4bd6d3bd0a8b824d23a1c484a8bb0db9f7a83f18711bb97150dfb010457dc8f35396020405248f18e801b515fb076521dd133976a8058a31298d39ac4389f64;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he2bd5998bbb4798c0006b36b7f4fadbd1c99cec5119cc8ed885f3131e779b372b2a0096d3e663d2dd4fb0fae84b858b7dc8db404aae64339801b4a606c8e6175742f6e9ee8c09c8fb407ac4b22ad91b80458365d76f16fcfc8a86f52b579eeeb98706cd350eb86b5b2ac7cbc91e725119dbe27d1b8de9c7c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h131563d580c27f63cdfa658f29b59ab342d7557567c986cb0a262bd23c1bc67f0a80ba1f1bd4a25154823366b0412e6abc6a6562944e75cc6eb6bd216dd543135c8fadd10f95696b67bb926c44fe334876a1012ad3d2e39ef7601d448dff694be015ffae219523431c0c4dceaf880517dad5eb06518dd7054;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1375f6cab468b165fbbccf38de35533456137969e62de1fbef089d03e52e2fe3dfd791f475d4ee9cf0d2395c2f236b1f65952a7019415ca6d2bbd37cbd7704ed88dcbb3e335ee20e99d9f0138a5fb4031ac443aad35f37067092a515cb582807b85032c2d322df21d482701aba3f4096d57b5473d87122f2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hab1f9b78984b116c3557101b105818cc39ad9acb836edd293ce15f5d7db3b75b176e08c2dc2fa61c4f1c2e8c71978e90c6d99aa44418190b666f8ca5ade1cacefaa2e5292401b25741c894d7bbfb6fc72d9feccce8d5ce86d9d90d95afb668d623205ab776a56973c8563712331f752eb25f382eaab119d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8223ee43db624bca86261567ba87709dabc154a7b564c92da4ab4e7a2b408b7a7297862dd33435cfa1435580731c4541b244eb6fb409b77cdf3249d0ffc58063ab14eb6bd13e814606a71636de064ced4beb1162ee02e379a1b8ee122b68b4708f2a4b2bc0010c43e2d85fae0c31ba3ebe877b4fa330d66c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h956c8fb19dc60d45bcfd5387788b76d7ade389cc0f44e0dafc76fb4c0645b4f10673d2d49b4c88ae17af68206c3b7c8de2fe564ff9db25eacc4f31dc313001062461939f321153fcb0cd4c502845c298bf9903c0571f37402b7b43dc6116908b63340e41868441509b41f1dbf99a7cc0473d6cab7b49715b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd19f0b01c009058cd74d18c34a585c6951ff4abdce31f990161f5c39660d59a63429af2761bcff1d54d1c65170beb81b70bd8e104d43e65e84a24724e991dec22c12bac8c436982da5806a1dac54654f2cd01027c05e12b3191018733d1a05054d166cb5a1948a412754eda21de3ea74d8e1ad1344e526a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8c2db4eef54007c3b9c37a81716c0f9a1c2a7da4088b4101554f601d80518231a279eff715361727fcef029c4cb56a14e8c4f86c4409155cd7d31f78ee88e4f7a581384c7a25e03bb489c99bd6b49cc06113f2a1aec567400fb7696b26aa562b5924b963faf87a3fa2dc60b97a8a66775d8cf00b9f82b25;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d3b0198671abbf95288e5cde7a91b972d47700450e1b61187f8e604d278c00f26b75f509e9230237b445ff8552dfd9ec6b2ace1e541383afe5cc7d64456e994700034e703fc1f6f7bd351629a9237ec473e835cc1f4de0bb59fb5897843340ad4c3ab989465e19911873aca7e1754188925b8d5cb246e2d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c4102a710372cbf4f0d140abfc86fd06e1bf9d5c6ccb6e979b92321c7e7440bed286d53c3b306c5ba388c3a7f0a55ce1bf349dbdb3944dc86962c0113be3fee1c03e8896011dd4abf585ad2ecb1dad3eebb80dfa3ea7ca0b387011a3ac99c639e8ae07851119a1a307826a3b5a100c0a32ea8ab10aee8670;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf75b4c3edd4ecf549c99acc820509880b8c231febbf4a3c532ea589cbb5763a88e5b4238d04e8e59296c102877f8e7a5cc2d0c87140d8bafc5b8afc472cf171c5f4687cf69684c6b0f77c237853134c1857dbddf3d6b683fddc622824958cb1dbeda0dc5121866e6fdaf84bd6ce31d2367b0ac7d7ce252cf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5f739c7afd2587f9f99a640dac7a18afdd3a8013c1016c29192e7d64cd7f43c51ec9aef8f5cde5c519c755d65e890ade1374006002b33488d151f189bc70cb86adfc8613eba6d27924da5a2d6b1db535f468b51694cb4b8441f526bd8ba4dd600890855873beac956e080ffcdc7616f43a2821abbd4b1af7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d8647ba24378cf466de5b1ebf5051d2815abcdd7c7c063600c8525ea53b8b43edfcb1f63c232494ae30cdb1fb3de8151b30d087ab5af095dd02aa61227021b5064d001f1b98abef924eb606e42cd3e25780246753683afa0ebbf7e9e5f3599aded6826742f1793bd7ea8253a99da1cb6e3813ac468aa7e9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149781755023150c908170ee6fb1bed742fed634a1bf107140d2b523a52632f02e791df96eccc64e81c5cef8ebc6ee0c5883fdf83be48d3dcdd14e8a740406448047fa49b89e75ec861864ec4155c7188340162bcb941d64b8d89088b58911721250e7a1d680e09c512f2fcdec8f2e7bf2a8dccc529112c68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ad4f73f50d4d5e840630cf3ccde5ff1c44dbd09690d85dfe7a8b435655111339fb0af31791d93712da9ee9492468dd7d1e9303c7f7ea6073ca323fa8a4c115e911611b75984ab0a1249a40b9b0bd3a71b0c57f59c28cc655f4afc8803ed1ec9f6c1bd7943f6b4d7a7eddfaf2f21be198ef0748d08c36514;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h134cc6a15ca43290cd4835259dc5f257421bbb9b1dfd86720e6431bfb4070c600f43f546937098fdab7cfdf029581490d41565a17b152ca9cc40e117f0733c210e4a13d7828694e2db2800c85cf036a6e626ef9045b4998cc4e173149b7e5920fde9ed3fbe4ab6ec5e68e8a6c9522694a47e32539c81d4680;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9fc12b88c287aa1efcebccb367deacb3a30c430063b4bdf893ad442cff5ec12903a5bd87d8cf89ac981d5b348bced2a5450ac868ff6149711a1fb3c2f5653b7a04d1f778e3cdb926f6201c7c232ca94e93bb56f4ef3171dc388ced372c6032306cd8197afa2eda834cd37eee1d205893ceda7bdb0621767c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h188bde3e5bfdecc0d036758f79ffad1c39de4b954cd2bebce3c788c8d72f472f7d6337b3d8d541e14cdab4382e762484a9c079f0ba4153f42e5d4244a91a93febd52e6770cb62b0515865f4fd1ac1e955c3922fccb1c8d000e16bc6feaaf8849868f28cdec6d01fbb036b5662ec8ed4ce72732906f5446b00;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hacccb2bec82a67167e230a8b0ee9ec0af43e4624185a5936b110a6810f3e8dc80eac5033c6451ac5ffc953434e79bd1f51077c77d696e7146f48bdee5ad03a6fe6d52be54739eec53e96c8173eac8c8eb28b3ae7e96d3befaf5a0e5e5e70686cf85697f88f40f27dd10c707c2d075328291d9046e3177f46;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h32485260c12844b3f39da0f93be9a2c0ebe01c06035428c0a6010ebabc804db058d43130d81f22b257a460d4d06b536625827a7c3e8585925fa40c8c1e47dae04a62f1acdf3e0ef702ca924b08dd10c9a08749816ef9b5cccf37aa02d6a466b96e9cc0e722d8f4b06302791342732cc9d42a85d189d4b2b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63b26bb83d8278f3d96f8221082bf363b32be7a3116a10ecff03d7dbb156c15fcb5233ff17990157fbd6f7321eda39f16d6d5168fdc882f3ef15e4b398d267242549dea36e5308b1aa8b7e41802f6597ba0735d75a3f82cbe8bdb2fd4fc4e3feec0eeb4553e3e9b7e7ff937086618f34f57d703ffb27db90;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h112ef78fdb05b6b19978c7694785aeadf0de881d2ec0d8ecf9f8471bd68e2c3f7a47f2bec35550f4c052a939b33adef92c2bc72c4c18048ec4c4d445954e2d64151fe47d98c3bdfe2badcbadc67ba636c27cfb8ed70711bdac51a7f318ac94ae8cf7145c0fdf35bab04eaa4d97791fb9e80457f568f942ef9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c3912893986eea490d5e7ad79bbe5a06d5172097a08b2c04f7a793782949d7da45cf1f2e13f8e8c6bf92a012de7ffe3857bb4036937def099a24fa915fab739956b3bff93e4808ce6e1661ac36441e26b28b2fade57d8d2b513668617623a0e02b4c42aefbe25b5b9bdc02ec921ca17a1c65ff935baf4885;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52857804bc15c0b07913b43fb3da2b6224697c0f1f7a8ceac2c9bc4fe7ac93285c93a8271c9add483e48717e3cf62cc9dc3eee347fc6d36acafe705b37a370f079f0948706e5c3f31a40afeaf5356f12ca01e66d63dbf558fe93a87687d45e8087031555332e5c975645ab99bdba70fa6a4c618602e6fbd2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7dd2bb058c7b2e157d14227d058212e620058ae422d0076e805a2df729a54ab42f779950de69194b553d287b64128058a589f901b0cfba957f8daea38550f17dde5e3d60b8ce7c3e4e56a3392421ba0d6fa148cd04621f3a324119a650a6b49ca27d60cf7c3943d4a6cc66d418de5e5a6b46e8e5b4e903b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13875fbded7e975d2a47e7a4a2cad58fc4f1b01edd17407e1cbfef1e0c60bfa1230b47d6cccdefdbf0a86a11beb5ed36c648dc1ccce42c4d78e29972e61377ae8440787bdecf14de5e5b5548020ca91274210553294963686834d4dabe32f5e820b9a0d25a2c1c05a0c5dfde71eb6628b5c24621a29e4dd17;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bed906ab1c66c2339571ef6d93ab778a5f5aff50f4aea02e0ecf4613dedb5419f6e015c322d060b9301b5a00e73e3afe8acb577dd83616c30aa8343b2c87126f14ec8460982d357865a38f5562a04aff8a9e245aaedcace186cab7ee595ac7870bdc67d8f63ac7cd4b93270ffb7ce03df09d912b9180664c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5edb50c98d3d38d8fde8212c6a31111d1cfc1557e92667539576ea0c96375d2fd7bb06846a2570a668bd94d7a68ba3b065e8bc2d279e42e21d200dadb5e95657b084d114facde6650814bbc775514aa5601031d93728bc4ee54e00f92f9b9ce0a63558b0652d588de244ded8fbdb35856dfc6c517873507;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd5d2018d412bd6754e06fe55e1a756d6575a4a5c4cb14e3067ea3a962160eb34e09e588438866393fd7d73cfb4473f58ff19d42bb1be8a2e469ec5eae1066be437fa881cb7b7bb06db04189974824508adb9895a09b78b17aa222d14e691c71aa87f384aaab71947acab07bdb4e8341daa82f49fef7bdffb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10b6e494854f7667c7efa3565769a0b4fd991d921c2e7e41c4258bd29802ec0097c6925fdf2da1afa9a8585b38cbfd59f09ad0ed95c9c83cbe8b0acf36c122d7cb428da7a03e7170d861d0775fb31ec789714720967a29e006bf9735c5cac7b0ad6e4906566a262b3de3eb9f18b9fae779c1daecc1ee819f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e0364e92cee2c895f6b09f8675517e7634d5fc72c306c62ffae4096671fe0a66eae11a4b30db1f712476debd17101dc636547170b415ce069f63dd936a5bd73b7e82f068ccced0e845ac60c332271bd387c0a5674e5e07e7d2fbd728e592d95be19e3a1c3b4137a1ea39f5663c600fa1bce53a066561acb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8051ecb720b03f3b006b6f5e19b8eb4700f97a22a4212dc7d53cd73dd3c0056376cfffe1283748c4e39417b7aa429f56be99075324c26c087da069af5aa8a41c49838e219137cbcc712de47605b0b093f710cde35df39a71ee81c5b79fc531d38aedc28a63b3378187534c7939b33ba6e24339093dc5ee9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10fa1d50717e0847c54312cabec935319aadb8b1f7a9dcbd2b9c2ea3116182af2a9d6a32d50133ceeb8bac24508c1a1b981567477d0fe25b07b0f92e188796b968d5edf777ae046f55eff5803ea1bbb1536fa876014a87d1c082be84f1838cadc512590725475e1a723584051aa059b1b6ecb9adeaa3b521e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1655922a2f547c8db3546dda374f7c090041f11cad061ab29d6bbef653fa2154321a385919e158b479a29ba6d43a097daa09ac0fcdd09d3e35edfcdb09a23f31247b5bcecb4a11648c2bfb6b886e0cccd27f5f75e7669eba352e40ca78401d632ea539869c38b52fa1828f8c32c8f6fc058f0c8ee8efc5daa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc4d87e3e02e27f2ac1dffae954d4f61702b84bf7eb1422afa2bb539950842ec32d76e5090a55eea6aee1cdc1083e75d3177e4c2775fc8697c5531bf13ac479fa392e2ab1781bb9eb15cc29a23bb5ee742c50d034ad2e3c9e3c9b586ec4cf2aa67a400817588ff51b2358509aade6bae87d4a39397edb7c65;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b712831ae46e7adba966d408b35e02cbc55997f26467339b0bea99339a13b468c96be5c463d92b177eb116cd5245065a65c2ba8337f573882575a13b0d4d235a8138ee17a861a756918f4d6bb564bdfb9c9a507e58fd896f80785c93d0cebc5c344249eee1662bb60593d694cef1cdeb003a6f3be9c63c23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a13a9f81bea99ff6d4341130b9c37ea15e9c0ca72849453f6d823ffe3526e2f95c0eb5a335fa6d2208fdc65c673859305d6fcbc493d498630d85f1698632c4015990bd14eb9f1a55ee63da5ee91070378088f9a15aa7ef718fc54af202750c87cf02b56d9f5ff13b5931d3ea3bfb9d38cc96b43231787bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1864751e67148d981653ef08c237761212a5645f24123d3db92700624807c81e5d55cf5b28b1c06778fca6d74f82dbea30a58d58a8fc892096f7f6d2b5c122970db32527d54282a9edddca597d2c09024c0679f7c9f7e3531813b2ff1f7119578d61ffa92c292027bec7843bf9b26d401874333563189e4f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eff3f8ced9de736b8ce23b73e38a7077ed217cf1b6652013ea003eea70d2933d39a57a7e8618ad99427cbd69acf34d4e8376b69daa0e427419742f8fff50ae139be4f6b98f0b8dfc957e72162efc445e1820a5e899c9b5fd1ba01b85839e14b79c5d162f904368052ab78ba59e413fbc33e2074b1df5436;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc06af7689f98150bcbabf978c2567043ef3f186e653497a685e2f8a0ac9f5c25eba212e578398870f6c00a173cbf2a1d29795ff2ca074df852b6d63d3310bf1a34912c6db88b30b1fa17984915168325dd6d05cd3e7d86afeff1217177096c656607d5d50a8ae56a899ee2c8e9a2e6a30bbea3328d4fd349;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2bd5119e89e4983f00ea8958262dea994fc946db0372d99d4ff685d4ca6e73174b990a76f0dbbcc6770d30a3e84dffc394f766cffc17ebf5765f7c73cfdaef2e016b6b6f2ce97adc4cfd2b379f201b0ac49b7ca1dc894f16f8e6104b8c6fa7056ae5997f6fdc3bee5e4f852508e9967f7db99fec19283d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdd00be0eb956c8ba78de3fcc2f86eadcfa223fba93b2ed99b6d45576375ec8af88b7b535cfd2501658667b41662d90ce5d895ac3e5ecab6d08d0bd16420de33706ae553d307eb715447bcb6f929a45b574fdb543966de020860a90b413f95af905adaff1df1416817895611da575256771e8692603019079;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d80e98fabec5475e538d03fcda4e1b8a442a4c6998558567ca62bf24b03c7c692de0e979aefa5a066b64b4013d879d89237003dc3f1c0870abeb2e81e8cdc26c8c5767b3c49f484a662a5c85daf102c458f6fbe819e34c022798c3200d7bda9857db7f3f29d8d229532d815fe573d216e47c66f4122003f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h391c86231eecff50465b07432b1bc514af836e9d2beb83a337a9176644bf085879026e87379daea28f1b8c73cb2ad458e37848cb1e7472cc2532eb56400b253b093e27a40e219edda31e14b216b26ee91d444f8ffb5dbb822bb303daa12815c9186a7d14906fc6db02af044805df7d241cf5307dcbd2d592;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h170a1977abce72a8c6d62be2c216df7f630083009fc19f9a28ef55adebee2bb723a4702fd26ddcffdf3403600637a7b36f7a3083e67acdf974a50b8cf65ee942937ec1b13d3b0119bb73bc9302a35359e1558d580527c7fb5979d347a161ebc4b6709978fc9d21a74b98f2c5ee0b3ebd830dad9ab578f1482;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d1477e42e68568bec51bbb978e05da89d5d7dafe9267bf3caf0a2f90954526cdc282e1f87e42599024d9af8096a3f26e1639e323ef55587b5d196c204a48058fe4d0be6b9d120157f55aa6c4cc4d627b6bb3d6aa22092bd7787d0113fd3efbba173a5df5e8ea3c5ea5e970739ed2f725d6f6a2e28339288f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f163cec9660af1520b377fc5a8430ebebb8f6269bde9629c6f7e646f688a455789d9463fd1d6264ed0455190b6ff5bb8b54ffac3ccfbf1140ac42c69860d64b39262bc26d20a7cfbc33c552e0b6cb23fc5cde0a1d07d925c4db08b40c0f7297e69994359ef0665c0d19d336052cb7964f716a174a9bf336;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8af922f0af48dee6e8e6be7b315d4201f223daf802d0e0d51b360b32d21805bfe0ca612721b8f47369fe0fe44985439a4f40ce5494f5ba161ad82b9dfe289235f710affc22361c756dd9f8392ce8b6b7e4e86dbd6ab4a9b39618201ada3e71f5b795887c8467c2439a18a769561880c1e1b680142e7f4f94;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1570a88142cd2b50585484ad1b8c3bf858a7cf6a56d28f35349b774ddc5d0211dd87eec3654379feceeb0bd897f03e5e7741025986a472f24d4a18b8a7f281d3edf2cd15b579da20ad13d5b2f892858ed487656b0b2dcb5dda5891570eb23535a98019013a99f83e6d70e5bf21975473acc76229e0471a893;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h114d12593552e1bedc708e7ecebf8af6123f60d973c814bf027b8aa3f0b7aa16f08a2119d63b20d123d121265bd512dc73e954446236c52fe97b26dd831059be5cd34c1ebbc77d0a906c54aa6cc92ca9fa4d29eb4d54cb7fb63e1323a3ad61c5b25a169dbd79ed6b1748b7b65523d48a1d1446bf652382c3e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbcea8805d0876e0407a76afe591f0fa5fd62ec99c832fb32f507fdffd25b4edee1fe85cbe861053a65a965adb4a238f2de297b0c7f579baea1b3a8d3f580b7292c64c498e7fd302b4b3165ffa528c879b635817ed6eb09915525fafd02d4386ea6605919c53042519de99c666dc0da0c0fe9107463fb4c3d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17260d133d091f1d73ecf596cc6663a4c63e9e04b01aad32c822204df667544822b5bee4508fe018346cc28e38b4f6edd3e1e1919eb826be67961ef41d6fccd4fa89734521b8a76396655d92cdf8d6ebb6d23e9817f3d29feec60cb7612769f73034a1cebf935d0b759d0b6e7fa6a0a3122ca9dbc640a5f9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab78d8474d99d9c109daea16a4078d58b468590f6bc3e1231a05afb1404ebce486106d3a0f65911294532c84f8a1ff6652dc93b122f82e5c06176aaa1f78ef9aadd4bb18dd2e9f52204765837fce6595062e540fd40f528183e596e274a4bc6e6682d6ad2bcb79007a8d12cb088ed00abeab2e84052ae88;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h194cbf6b49e46d3e3ed8ba14e8d9d118661a922c851aa1fb51a6173999655d411984bf5c04569b9e8471802145793fda43956cba506c57a011055f682a67e3689ee34ab625258e91b5dcc46d0b116b76bdf0c8992b9e7ef9ec580ff4bae724108f0d2f053434ad360e270da683765b5467db66f781d85c8c4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f91ceb616db89717f032cf693d864041498ef0f55347dc04420c62d23895c6f471f5b3870ff13b024a1cbb54fcb29c584f4a1dd967f60ab81e33b09eb648abc799f86f44d6c3983a773137c881de31b0ee2fcd0df2f0ed09ab336aa1b596e91ebe3c88adb37f9a1dcf585b6606f89c5ae8150f05795d724e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d93bcfc9ff675bec146e40ae0e415081579baf46adacc8eb420f300696a63d293af94fa3ddca365cc72f254e56abcaefc346cb2e33544a0b30d58bf9f88df3013c0ef2d09d68d0a1812c90a0dd22dc5a0a8de2d6f0658d4df66df05be3ead566a67eb0b90f6963785e8a9cebce0a4367d5c4bbd5c43d8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a67db99436f007b65f84739f016655165c39e16a3423e98d3f675bed93d24ded55bcb8163e930730a36f6d845fa371a3405a45f69935c1e63fb3d6a916ca860ba20a7e20eed60000e1922b35a48354b862c2b20de8ceb9f59ffebd1a7b3063a9ff7b9779c28871410f46d744f231829778cf77d341517f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111fecef198fbe47188353bb69a940b91e4870286a0d66836b94db68332ff60670a0671f0d2a9675c8fb32f201be0a3047b2783bb7eeeaba48b97537a49248dd717962d8b16a36c760f5be7d7f5c60721f44351e9e3b85151f38294b2e6299d453d5c32a9555f91d2e765c1547794ad942ccff889c2bd3944;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b90f2eb229911cc3be13c05a87e8297d189b3538423a40c484701eccebb394ea5e7707d09925361ef7420a2ca372b74f6c72c6185f549954906dd765aea08a442461aade9b6b17ea8acaed907df67041730977e317788b1f0d8ad1074be411626157c5acb8342f7db7e8f44597bb27b5548022e0698eddf3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd5535deaa2bc60e893ef61e3d76098bc63d2d1b58a1eb2ca27fe6b9c05fd1520a7f58a8a57b8e483dd1ac525c764fd244c11f8b885776f8b2c974091e0a6465c5611acea5acfcf27efc884addc128b058786619b1084ac217c38a194083745228620997c3c89514b65c47151ec8e6f3fadff37796cb71d8b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hba9a2208ebf3bce07254cd79e64aa2043a51cce518e3d64ad1ebb8cb0f27f21bd38606a39a64e8f1f5bd8b2113e4e29f6ee841aa62819825ee2f6375fbf4441d7e472e06408e59b71a518c12f02062131b88ba5ef567f221b6dbc400d4f2e7d19c22564d23d0c71bf16b8515eabdaee4735a00a858bfb4b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he2ac8e67c8d41877c6df69d5786c4a5ae44653ad58412a95b71ca391b80cb7130a26fcc25cd966f234da62863c90a8272c72937224b75b01b060ce671f35b3e5341705e4fa0357b3893579f7d924be0c4a09fadd18e3460ccf9afcf0ed006e818869d6a1394efdf73690367c632ab81e1816c709353a96ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15af3e34af2cc036de92cf4e8c21c564bf479dbdc21c25e7efbd086f401365ea5c4969e5dcce9acf368f50a922918a9f35af002a3507a338596282e16c2118eef77447106a53f91b44b946103a0156e7c5e96d1d556176f104f72cab39d59b8130943b3d161499c2b9a6e7b6fa17dc32d520cedecab6ac19b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h123b5878d49dffb5a221b7394f13a23feb2e9aa5bee6b5fbb51e69cc98be216c29ff7195df62abca3dd2aa79446b270eb1a48535256c028eafa71845fd58f2c303701ea73713dabcdcfa4df02fe42075615769e38e51e0e62e66bdbfd0d169a1c47520b14d803cc86bcfc4b9f3854d5fe07332d23709434a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b3c26c3322821fa66e27cbae2f63f87ff8e314fd9e2f84326bfd4ce8abb339383aa2bdc059a521b62493cc99b600742cba22dd5beb7259581a7d71e509dbbd240f5f9452b6993d2d1e6be6ab2e423076738d4276283b85855a2fbaf4a2893435172b418d1b22291c9270706d8b6d4488369a5ef2132f4a75;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hff7527f917bf1e76841797fc195965c6bea1826ec0ea4dd06e7342d0c795e1a37d001e6520e1618099f57feb69521e7c004e59fbb284e93c6fc064d5454cbd98bc79b202e7f873c0955e2b09d9b12b1111b636e2733972a70ff47832d87532b9e99fc644a42542353c6c33060e78634d34832c6ce1b23b16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda7837c2dec59c126b7fdc7580d6cf4fa5595d59116a8ad31370a4352f9d11e8fbf214e33a6f388cc7d38a4ae5e7150f032ebda3e92addff6c4b1583e97f6d39c0286e63252457453c6b2d07957fb8e488192111d1ec0032e1c3f9a244a7d687003760147cdfcaacfbcc1bc9d152eee9749bcefc4f9daedf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d6fe89f31f87eb2e6a4ec0e1544962e8e992bcf03b635a188c9adbf54f1e311f0377ac40a7ef3be4378b742f0f578e8a6a2d7c70d4b463140ede9a62b2c7805becf9f62fc99e01c916ea4a8286c988edeb65c2b5a64142b54363a6549bb681f1673aae8f60281ddda2c713b81016cd16e61bef6aa8669d6b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12608225cf05c0b596407b09c894304a499e142f131405174fcde207e6c717b02301f5937060e6d7f00d50e4c236736a47ba38281e246bdfa6dcbcbb1848ddccb85aaf608dd1aecc44147b6c9b3b1f784b9cc605c9fb5642de57510c8c58d02c6c07de7e21ada752947614eaa31a39a1e2ebfe9c7e291378c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1200cc83d9588a0c186e7eacfb6e3f09ddcd04384f879382a7007e326ae8d5dd6ae14c1bdbbc83a965c250e9c3ae7f044c0f960fe54e8a9cedc8d72b5bfbd2f2a451c3f284beba979362409fdf5dcf6f21d5a074b1d06e90ba583bf4acd828dceb38dfdbccdc12db715324d8f538ec68f391d988a6a6bb197;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15f40a3dc4733fc1330071d46bf1dc18374e0ac468bf0d9e1224a824427dec343c2ce69905b7013b9aed26f01a300d453471fd26fb15bbb86254835c807d32b499a777de7ca4dd493ce6c6108efd7fd0036c319ddeb7a438093f1a811f8efb4d2fd8b73fc7c953d60dfd73585d91b748782970a67eac875d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdce6e7f5e48aa88e55bbcf4d81dd01ad714cb950055c60011af94e88c332467aed4d01fb730d31ec23285a34c09862934969d7da0cc10abc0399e5a39032b952a94c1832d166234be6b23edf176fe0c6d048134a7b2d5bdbc01e19198360fda73586ccca44a860a3acf81a6214f85dcda3447e48f0ef03c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6eb0e8d7f26bdf9f47b1ac75c93d7d3cf10bb5a1ae86dfe8c3a298bee7ad28ce715b053403dbf296d88db90e214dda6cf232c520e9dc01908495b712ac3e691aef376f72e470dc347db246b8f8a47d13c4b6c03154f135dbf03ceef7d89f947b93f87ca8c8f0a7170bf982b1bd69184e00890661e167c18d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18a1f8227f6bb3ed8b0916778c529e426f6b2e09cec68eb3db41aed1bb4564048a1c21df8260cb09deb47b70e3b7d354a7a2d2285aae9182198ad39d68505bd896e68c44f276c09e75970522dbcd9c9cead6983ab04eb56acc95337bf802f0bed2316b4e74b14b13be121c6b8b66c0be53689dd31960f2704;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15a7577bff8dc820ec00d563e0c1dfc4ea8c8d39d8d7d950bf0723440bd920d3d90949682ed62e39e6b5f837b5d7025bf1ffec81d4945c1d8c0415832aaa7c43c3985ac50e29b87f44807953aa8c2d7fbcf34ec0c51b20c8f584a4efaf3ed11df13ac5d600dee63c816271e730b194b135fb542e2184ff1bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13664db376fcf37f4eb1facdf448e71a42ed3b9c7bdd5612adf4b439955e75ae09f110ff5313539391ca5847a9738a45210e980f9f7441791f1656f961c7ad60a1a0f991102cf24ce3d5f50eadf360f69ff40ffa099fa90fdb33d633a5beaac14cab90ff6a3c83f3ab6746b252a4f6440f6ea1162d3823ff1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d72c92b589f403a83a944da1f67b2f5976e9a4f94c76690f780a77017a44f5f06991da485694f494daeb2b5c3042252c337691c442eec9c59d4c6a6ed6132ab43bc219afc077756d8c1623fcb8f20c8e9e8e5992aaded9fe85a458284eb7ab8c443242e73301cfbef41148bc13599b940cf7a974701e695;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf533cbdcdb3556f3c11bcdfdc36e2797e3c12308bdd727c36b6b2272f3a354d2dd1ab8d536512058a138d5f342017863ba887d826fd141aa1e38961acf99cebb99a36d16fb440054db3f05214197ef6e878c5d5cd1371b459d05eda1ec7432703a05be03324dcba9d332fb9a8c8b4c6bf0e9fc3fc65c1a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdaca430cb38a667891e48ded0f33f3bf27d91082320c41fa43a1bc99ffd7aafae58a078fe231ea7941a12169ce400f3adf75a8bf7660655b439f53dfe8a9c1d566063db4b25d7a3d846ccf6f223b85e39876b1eca439c3b5c78c23060c8f06243e9824d7e9ec4ba7ce2711aea0b2ca13ced2e323e88ebee6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h189e3d13d774819195799176480c64bf565089aa2ddca92d43ac6f9bfdca563bd922d92baf7dbb7bd781477d59f11d2f2e8add49da7365cb8cc74bb22e12f274623b403349e0dab39e121e000502020c8dbcfc6ceef58a55e0644b33596e35248f3f82c4f6a5c72c28ccc0ce363fb2cdf3294235329e1bd27;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137e97dc02b44b9e39de1ff9220e8583afa2c48b53055c350d5927751a075951ee8d58ca86e3a1de2f9961b0d03e9dda7c567f02980237170e994167a928dda57570603e8987c66ce9138bc14f1fb85c62c74a5f63403bacc6df2f3067f732c18f34c600c13dc7b5e8825d1c8214bc2f6524a985d608e31d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h148b13943a9d3b46d111586d93a43b7989df27955e0c5615cc46d2b8eb5aa10c002eba57dadcc409ca153b6c71f47cb3e1451ee921a8303c4c0332b1a4118dbbd427e1a05383ec717768a68db11a994ce67bc545372e9abd0e9c8230a627a69ace4c28d93de78654b944d3bd5611acbe28dd061cf9714f52a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h160a7b54bb2fb931ffd260dae8a92b23080c984a011eca4945e9a96a2d5f94c7d9e3566ec6f51e3e7b25721ad97f2049a76dfb41d909f45769e605377f194afcc0d5106307f59279ca0fc86ccf993723fbcb9b12e160a3ec581da1778de48f101f3827d8065b24abe7756d293075044d87c2654eca9f9a4c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd8bdd39d3e09934097525ea0beb42f942953b8b03823a974a695dc6da52cbdd9795c7b2a42b5710eceea1d9948328de127843025cc963008e708826f7b55933b8a316b9575036b036a806b949e1030261fd5f291ab0a0f3e60363b25980593c996bcb94bb9100c406764acc099bd3e4e70f7909f7a6a8e5f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f07354538154f8c2e56d3838e17b490d707053ba3f675cbd9e6855bd85f21928bb28441e33a34a93a678e0b018fff41d5f57a117518fb8a4ef6f5316df494af0e7781066804d249c033f01305b70eb7fbf9f1569bde7aa8a29e25caf3bcf1ba48f0a7b5ddc43947eef33b93dd469216d1da776188478461;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1210837d122d146e301846359ec70d249ea122a6e25a457f8f53c806c85547a9fbb45bc79cdc8b3e1b79ff422fc51f7744eaa45f41c0458da99f2394dfd1977785aca1c5d0495dbf5d62a95fc02858056ae401f107fb685805ffd00b47496e1dc3a36a2b79939756aa9662b0c3138dfa580f7cd51c473783a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10e2068c431893f13fea30ed768bff9f3605d2903695b2759c77f358706531e7a27cdfa54fab89e9f60f9c4934e4f179ff47173a8244d2b0e203f3a14c5014b67a9fddb61781b10e2fadbc33b4bf9b2c2a373bdbc8cf7f90f287198dfc051f0720cfd2d3422f098c18c842b0b47159a30b1acefa624776dad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc83f13683121a60000c3508c8c479d4336b02a95fbd472f77c9e1c74dbd235046c134a1944ad5d5d09f14264b131a02a87d1ea0f401c7ebe91d8b00af7b2aaa705c18767d52c908e38d69729c9cd28a05137f77ac1dd209b60358f5cf94404d10d354683f067ac4f539830bdf3d1c80dcb3e0ca861fedbf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h164f7f764e192977330d1bf9b4a3d0843cd90ef75437c4714001c77789316b095fa950cd8b4fe3469ad117e8d060e0221a0a581dc122484af424fc32092afe04f78691a7f0566aef697aba43347ad425261afe8acd8a6dbc359d906cac52a69e7959f7c832e18f69e168f803d5821a0cf42a2b616d3d658e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190980f3295df4b7e78eedaa36c4b2d8ded6856060b6285d673a039378dc8cc4516e6914196626a26a8df08cbf83d16a11ea13291bb8ffdf8b769289c830d15939fa544308a61ed64945ba7076110e5e3b29b1dab56899f7dd26712610cb1d331a998973c54e3f31430d7f56cd9f79d409b3f8d97f98730c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d354c9849b5c1239c626298a0a13f1e3d3de9b2fdc717678a535946983646040c333fb69b3e3b2339a20fb35e74cab6cd308a136b9a4937f0492c2ecd006ea294ddd425f5e87293246f628acddb8b42061804e0ebf7a6158dde2664304c1ab004a1c24465f1ba688c41f8fb8e476c1fa0255d7eb036fa608;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heac050adaa86f32a9e8fdb4b9d2bcaa147133580b982bd8bd1076dde7c69a6d616876e53369f378c75b56c447b9cd21a2a36730e149c63634c91bc4cc246c9deca40b73193c5c9d3af7e64b53c7ea95a5b6d9f4246199ba54bd536198da805a544d7460253e080b89752e8dbdee52b580314a99f318c369d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h163c47cc41632a788f0e41b87d530d5d5f38883b7b7dad67242e002a44c41f1699e928808bf3d5898ece7218519bcd1871745c6392fb3c734ad629a342ea14d8591ec388b0a381b7e3f440047f7f1c826ba9b3057ba40fe25ae3f1cec198da951e0addeebedd98a4ce6e0d14eb654b9a0356d939825561196;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd90fc72444c27f1ab1257f08c303c7f5ba7f8ccc25511b25ad28af5e0eda71e70e06dee480e34321c1dec74af08a0603a2143bca09383fd13995665f67a5105d0e082d5b21ba39588b4b2a20d8b99bea1b4444af7b5b3c631f39e6520687a1e6a9d4b0c48e38e5d9958d3d1d019a5f0b53e5740a981b15df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h39be2dc4c3fa3402c972329fbbec1a4f6be52a07c72c1cd902654db91c5d60bf836d6bf04e57a4b8850cb5eb387617d9ad4016a56ec99f830dbdf52f87ddf0745e13ec7f1d79a1152e3847f09bb37ca70285ee5046b82045e37b5e77cfda5b5104e17bb82107c1507975fd00c1a7a92f24d564ddd5cbedc8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e35a207adf2023d46459653c47061098fc604b51bf41ee6567f01fe9a06a3489a6c95c140fe88d50686265c83e11c4a19915e5e282630714a939cfbfa10e77f8f5d3363c7f5175cf574e0712622c8137f308603306270ee360b73dc5ba03744c9f4b9beb477177525ac268b9b8168520e16379638b0a9f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17544b03a797ffa27029cdcd0ad0d430d98403975e4e5579e7fbc298384da0687f9d0d460f9f31ca88de98d83d58131e02b7215efffa07a76ec66f2e071b5db389e4dfca46f4670a3bab9763eb7d4db9a1ea7c8d0b822b2a8eff59ecc130679619f9c7736792a23c7f0dd13ca2522bc32267d2c7140f3a894;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11eb63b3d220a8db064d25088977c39e56d0e0663cc2d9919edb9b640dbd5193a9e56fe1e38f7f8dd24847a3a0a97d8e547c0bc13268605082a4359f357f5a9aa76e15008ed8b3cb65c4ee1a30d514a398275b4d199677156cff93f6f1aa9d17d7cce417c2ddc2bb1d65dffb0493a27a5a106db94a5574a9c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f594a5301d1cd6471e9c90fe622da59f9ff6d54e208bae796b67629ac2dcf84625f67e060f95d221aad05f4c7606c5014bb35df3797f74d4b6bc927f926f077b179ec24a536204b841bec2ef7076d809513b89594c73389a0a2e7564e40820f5fa3081cb4e762b1b2a02c6f0568878c4124a80c856411de2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fb1140747a41dfe860c830845c9d5edd53f03272bd7b999056fd598eae4d2a7fb7c3f5cc678e64ea77536ca2dbb013e3fb3f5b911705291f0f5286124c29ecf64c2bc38f1660b5673a70f2415bebe451656310a2ab6f1155e3d6a97c87b0b8e0557fbe925c77738ef8aa2c6e8a820b0bb59b2f0677291eee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h42ddb14dfbd7dd521ef674f9840425925f4bc03538590446ec1d8f676848dca08134c697c1c8aa2e63ef1c1ce96b53e6715845f2daaf3b7c45137e1ac96604e69312090759d1c170cd1a7932d9657c3e72f88c243f37382c3f97fa04635806687df0217fe7c2a06d44adcf7182ac32a9cfc1747de485320;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17061b10ebbe21f7596fc3937d0bfe8eda65fac8d9e1295049607d789bd9942fb7275c0e2d0e2197cafa6cedfddf3fdb36bf150c534dadc67bd37db2cfa9ec33edfac0069ce060cf39d95d11c03936cc5ea09a61eefd412037bb489326e34c90e1a1360694ac1e7745eb7fd63405c0a5048d7126af1107268;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfd0512573958ca4d535a7490689f4f484f93e1f78dc59d61842409b35e4916857ffafd65b80acdb076e2b63b5dcb552b08fc8e7c59dca2eb730cf8735390cc8454e1aff4e3e17c95131ecab60ab8501733ddeb01b05451e2aca25636c30b6562e6f56b2a8eec1e3af1bf9f335564f73e305c7995eeae7396;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b542321a8f5d857134a8246b79d9e2bd5b047c0e7b524db45dacdf9d839537959ff0242c5d46c95886c6d60d5f4ca0430e024c89e5fd9510612ce3b4d349cc964be5b3268f4312ae7e80df31c19394c19bac3e3537f3e669315e0a3bc7afa105f6b6cbabbf2ec7d106cb2a85e7b25f11e25ed4112582451;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h39d7aeba3dc710faee6b57bbfa82d1bc6a1706b11484d5698336dfad1c348c7475534716feababe01ec2a9cb96ee22ea485d51d9b21418f0aecd83a4240a22649322068c923106d45b58cf73639f8f53c1a07c6f01e93967d82328d787f022a10025bbb362d4b51be4b9eff5e6e872193a3bd925e6461ee8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f2246bb7dbe4d9ad44fa44034730a1fc4f3bd77ba4c48babec905f1c03cd8b99c288dfc1330c5a750f9048b6541abc86359bc40b9fcf9f7a45ad47595b11af31e9578938c1fcd12f22682997159b060987b664d8bc89b7c1b146748a96e40312122c1d367550d6999ea802506aecec028b87bebae573e9a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a611fdf5e72afecad06fc319c2c524e1959a1faa33554ffb3fb54043f836dfc1820af2bdd1529371230d042ce758b816d5d385ac9bfd180210208cb62ee7054ddd11b58198cfbff43295a274450126656d7384856c18eb7ba5be70e18f92dfc260e3b3c27edc575ac2462002442209f7f928704aad6022d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de00a62ae2a6f736fd1a8478bdf29971c8a99838b88ffe25720972cc9c7b7c0fa61d1ea67ea2ade508fe272e04b9d0fa3b33437772bc9567a48ee96344d0c0821073fd89543cd21641b2817bc9738c8c867fd7299698e22ef04eff3fb5e00333470adb4b7f6861550e68f696854defd8c568743646e0ed9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1507b04b2040f23d35262055ac2d64cc33a61d29d2e3c7ca7b58caa5a5674b35c42d454e419fb05ec2f4b70e5d4109f6430b16214c2b59db334076e87615cb1fb0f7bc2f15cb365b6d93e5c8fe7b2d211aebf44a1e160e433de0d5c101332a74acc984423badbaaf51b52249b69bed9589c1b424309f4eb13;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90190a35f097c7293b68d4376dc8b1c2f6dbc4bfde19846d90ad22840edd8f62cc7507e8d88378f47f75b53f90a6100f527c4692674a72c03e91fa55d7d8e2e21de624bb8d4f49578635b1c6816545ee3a2be5b6afd395ff7ed5282878373bf847c09c6c443fafe860777aac885e70218da60753fd912c0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h20eea10a95e25025de1f9d3c98a5877170861467a72ae16506e896ed4028a8a5687aa41eeeadcca0869f2ec2b728340fdd1787bc48615a083796188188a9c90480305cf4df69b443269b8029e18103c875479b3b4e49f2164693f54f51f8470647d761a884854c8d22e5633f797dd406d216416db3d8bd9b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfcdef07fcd74bad688e435862165de865a188e1636d2f82947f2f437045aa0b1b8bb1740c2403bff431e4e68dcf524e29a668e46dae8139aeb9f212824138c9ed90fc8b592f4aca30f2b7ac2325cb3459f3885e63c42bdaa3d1300688f9b87941a7ce6e9af5c9757bb9d76226c2956f75e05deb92ce063fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e63a8d270998481abddae28115af6590f1099b4b80266b28536bea63b584c3ee328f404eaf0366e3642c1718e18cc8edc16de6835b647e97e72f86f33f4e390d3e0326b4d66fd5adac87af9a4081da11d318cc7302b3388e037c1d4a1411949d2850783789875ec89e96d7ff8e28c4800998295c8df6323;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f65595130eaee5fbecbfa230c2c43ec977344d80495a5b3454e9356a9b34ec2737b2da2a87b1ee16d4fe62647b41eba8d3545e3d9c90aabf120a55a6b6819d9df65758f769ee25c0f7152089743afc49ee17fb23762ce4d7a78290f50ddc3f07ba73787a9e842ad15f747e2c60ff201d60da2daf2c5726b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfe178b9ffb55e80186725020aa31d7bff85336eb6fcac334ba3086d23f286022cca9d32acdcb25fe46e1dadaf97414396ba2acbb425e0bb524d38d9891aea75a78b7ac47e40695cab7faf06909e45e5b891ae0f326bb5fa0c5060eb832ddee87ebe7d783bf7ddc0dddf8948bdc7f609099ed707dda213543;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0511e9b05d743269e5510e15cd12a4d602bcfc4efacd7495979f81cc13920eea69f1d224e90744c9c2ec90685ce94448c40578d971b545af9a048ea6ad633d5b3ebbe928a5c43a43d20325819561bf1b372a8ba39bfb276708ce8fdcfa7ee32f80e657c556f3166ed109723ccc778f713639c4b40d0f3c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b878a78c82d1ab78f84900e43079d9a3738f7fb539104efa576bde5eccfeb460cb7e4369ed3974cb81fe1f2a8f49070ada9b4f0946e42736664f708b60917dd29da809d41ce22fcde019f7fc8f7bcce83c7a3f79781dac77d3ffc460f0810c5125a39e81b64d5afee42a8a72556b6a00472b082ea5952fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14dddc6559bc5df9f9f2d4a2e5673ff46257d1285a7db4d8602517306ebeb938fb35764addb419c50eefe15fe9ab09ec183239cf2fad8c5ed272dc07b0118c67ab91da25da4bb2c6388c99f1e53c5fc9ec29412babf9a449bf25d99444a394093c1982cab54968579caab26ff16ca1f529f91d62f0a03f2f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1badcfb1e2cf559b0b522ccde346eb6b797f840daf9af2240d4c29bccce06be8ac5778cfaab813c545bf644d4bac6f61cde94aff3dee7becaaf572419d72823e37235acbe15574b0d1f41f1017bf618a842c6b22ead36fecacbd8f7cce27cee4393b39f9945460e318fb1d09c681d1e88ac978c59154cdacf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13da6961d518dbc170826d6d0da01950cd8b54855963ff33b75b3fedcd70345617e3f9b48b804bffde9d36e343640a34f4506ddc248ed2a5fb9a4b9d17949230ae26cce0ca311fd0e43a344147ea4d2896f800aa47ae97c05ebcb88c8af31b76fa0f493816ef6928c6df8349d5905f36ceb34d1a3d54c673f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd6617ec166e3631fc478165a6967435a22a466e6df9652bad873f2fb6e12d7f90629219e74f857f1a4e10a36a5c385e53f8f85b48d3632366675742600758325a2b84e4dbf829ee9595f360b0ec8816fb99423fb473fba2e28be97aa49db2408d3d60da9571755b6cd79ee0a8de9afa1beb67846583e0607;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h107681fc4064b86ce60afa4b3b6dec32638031eb51c6fd8fa119c76cc45ff267962771ecd657b696bde81d1c3b16aeeb4b7df87bfdfb860b7fed5bf549696d0c6ca2965bbb76312c0afa2c7c82f0816adff348c35bd0142907ae64cde3447089fb4cfe91e05d6677aa0d168e5dde6b26823189da3d6823edf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b41f664dcd9e76d265f51cb3f902b10c3e957d140a42d5919cca94d68de1aef0e052a7f161d1cbc2915be27997e8500aceb38f0b17ac8244dec6640d2f25ec10c02aef4e045f2a16a2892f4a2701ee5eec129ce73fb2ef132c75bf386331c5f56b62f4ea87e69b64383d5d208c9b22047e8bc7b539cce68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f5aa9febd5d5215de6a60b8ad9d5868050003b76f6a8e53d908c9e830f85dec204a18445953d2c08c552e60804a96a62cc26d9659ffa3cca776ef59ff4135433a58f1de3404accfca136e455f80f96cc57c3d60553143f8c17c4d41066f24299baf66a0ecf7e4fae576c79a3bb2d50bee9f78ed040891f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a3e990448b76dab747421722df7fbad8d46c64e070110e0bbdd4cad9862e51f222e18b310117b4d35525d89af2248cc982d5c7f1710ddc099a6fd4d82fa74825fc0796d73afd6b1e8da593bb9f26197c571ec72bf1ea672b9e42a9a0569bcdcaa3d9e2a331224bd3943d36036e345a65c83ab304b629e67;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9c19edf60378cac71fd20dde5fccda843e9004d086a9ce578d9fcde75b0340d0118437b7ee3e4b97f55ec9555964d17adab0c3e081fd0ca56aa8803388c5652c9574f034e60ba4b71aefe45f7a143c992baf5503a9569ce665819abfc40adfcd4d2f3cd19a0562a55cd39db47135a78660fa0a8ce69980d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h98aeb0ee7991dcd863be795fec9d0322e51285c02a4259a09080f9f169a414a2feba5b04123d4323b9240bddb70441e509ec0e64c5650257a57eb04d14553938f7ccb2f060aa6595734602aeb5c7e42663a2d0e628916d14dc0a6cdcbcb4b38c43997b39fdd921e4e78a844a05bcf95febcb893dd0a13c51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10bfc8128be3dc3fed37f79c41ebc0474c1df3055dc1cc678f6fd0ef675f98188d5328a6907f2ddc2b07636e47bd4e272712607bb7ef12612bcd4498fa177e435110473e8b50e13ab508943ef930864ebcebbe331665200fed5e89ea662109310fa1fe7bf65f883ce8dc2f68dd0f1b732a603e6385bed4db5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b350b1c031d9a5707241c1ee4b351d69fa39ddfab7c9870647dc65e6b7e4938c370096b6e68f2c2a4e9f921e4a9e74696c536b121183a30d8fc50dbd6b87dff3568eb23ae3211ed43d51b41e6f5fa2669ed289c9afb007ca09d1efa4747a1f749f664ceae5fa380ed9d7df8522743a00d4de5a4ee13a8dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9365974351584626dfb7f6c891513334d1abc6c6d555a6b287139a4600a88adc9c8edad7ed996a1a1cbb614ff40b69b55ccb0b8d48481996c6867418363fc10b16043f51568e3ff09ba9a23dc9674a5f46e544682681ef9e636dd33c923f325bc477af54ddb6f85527c903184ac1a3460a979fde0e673e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa5d3269d0c620bbf4a01caa06c8adedf94b837beb65c0f1f02640ffd8cd74a1c5f603b23d0932f012fe6930d90be53537030e275f842a17850793b2f98f87ed64ff4feecf7c050aed34edad76e3b5d66ed673f1f70c07c9234cdb5258c2a7b8d33a769d568d694525eaa7c36304201238d2aea29558ec83;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h824aa9a3b3be068e58d86af95001c6f34ce8450a887742ee59d1370e3f7344dd1d538228958ae535656904d17ee20f4d3a2d6f243b615969e1a4d0dd888ff2e324e9da0309ee4f95c6956cb8c4a149f9096bcebb731393ff466433be7dc3d247593989d2f79a2090c2f11fb7f63b5bc8d971e44cdab62c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4531dfe7f78df454feda12efa23ea021414a4aa7ca6022b31bc81a4dbec1d31c4bbdfdf8bc579b6a89c66799c26bf4dcd1479acbe5920fabf5da1dc266308f67a3ed23d8891972dc79119c5f0d0c2ce6cc5ebf5a6c2af0e14a63b2943c26211103fbf5bb5352dee382dc4165bf6e160929fa26ea13d238f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcc56f6a448f1f4e0cef9a1e4dc66406bdb5e5613a678a8ac845385f76edd7580398de150620896b689ac48e7c83e7ccdef58754f517d7a1dab4ec73b067795631bedd82586ff1f6f17d323ec89ffef80f22d897c921825a6b2ef46195770c9f591d704d66dc022cf63d184bc9c8f47b92977fb62fbd30f1f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec85f1c349db9ffbd0dba6feb03027c36c78454d4fae63c1bc04934537308273a952da89271d61c2c73adf85239e244bf301ca1e13f60020f51102ac609ed667b9881d3ec25cf2ef5d279bb11f38cdc1f6df05a6b8b7e4d3dad4332dd9fa91f62c8f0aeb9f3e426b3cc8174d3df78083ec9639ef2c8f2b48;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18750227a050f31b3d0c804d2cdf7d84c7414612d46f3cba67bdc5bdd9aa2e668935666fb8c569af894791c68e22f438f3f333164b5baae7c8c3196eb78f4489aca62f2d15cc675e2f85b71fadb255f5df2b2a32c77afbaa5d072587619f5fed15ae460b7a50d6cb6544066c87436d24549003441baa34435;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ee0c4cb8ae6ffaed33ff07333fbf7e442297b1eb650b179248aa96a6220b4e04c230b5ba884ac4cfe3c2b8618c489723d0c7c18167a42df107f45dc4a5300b9efa4b89f67be7bfb9a02394c70f232615ff3ccab8db789592fb98433d7e59397718d9a84b31fc3af80ed05ffd2f5abce35d3c0a698e5e016;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52018613118c7c836f43ba468361b364b413ad2668875344044a8e83d2855f828f69638f50d37d275ce2ba3e5de9339d0fef2497100341cdd103c13cffc75c6d0dac66ac7cf561c6b5ce3462bb649611062fc00435cbcf48023ff49679560a0fdd2ff55cbb78b483220b882cb0e33b07446b17c9173b212e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116ea49c1606f518d7bdb72904f2c68906a401f0258a1847121804f8fe42eb12f7a528a4e887bfd5fe091387f2faebcbac64807ced664a6c87dd0d18d94000a5b6ec7e23b5caf7b7f2132555b2fc7b71743e71d9fade06a39af7b925e812f05b61a2b0e4c2dc22f1f8a164294058cc5b4fee0aba759aa9697;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c1c745a5c244b3dc8aede02208c44514a23c83925ff74d5bcca6a70e38e9f8ea1d1ab628278cc5eb3911e462c8b61a7faf4a82c115f74aa8d862bdd68226ebeda47c26182c33cf9baf32631fd8fbb57deae8fe3adfc900709de35e5e6b880c27f4d22267262e2b8f235c2d91df6b57b701899cabcb87230;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8287b774aa9bed6deba0f27288b73e2583903d68cb91862610000b0c65de7ea9d98101b1e1b51fec506494ad2844444ed2cddc0bc14550e2a6f81aae65b35bceadee4b250e0bd3ba7f99d0802d86f4822f3f23bd2571802212dc3d2ef61d5aded3968b7f3bef48c7b6896d61899abeb6bf9ae19542b6d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf172bf42261612319b68b50e034baffd0f5ccc779c244be5ab35cbb4e065114cdf6db69bf0d5ea0c8316f13a1ad5045bc2d1913c3d887f2821fcbd860b8a19753872d84422ccdfb91c57aec055c26466cb00863faaa993a0fae3c91e1e27223e3a0075e7e20d8f8c0983c6a4c46499c41518ae13ac136789;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h176033fc001409ef0736b0d83ea24bb0051b0df480fb6ae1e975db198b38f637ae1510d378e6312e0d8bca0b9b39c5400d44330d9652aa50b7cd9ac14a1a42fc31f79e34264f4bbf9c4c9faa56a6f9da59b8d624f682b772e04bd748b758b973bddb1d8ec2af63bd69177327d7e31888e0f6910321ca46a7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h85d4c85311a008fbf25217e8f53d7914dfa4729374e858162d5724ec178a70755080e25d6145669d5f9a6b35286a916a270e603dbda253eec0df4a6b7a3668322e247ebe92718362feec40398f6b4c9688690f2eb3d28709f501e68794d592007bff8f6d189fa95d924c689366dd5ca47b7512764f1b99f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18921150740d8e10750b024702ff0b63e3812c05b2cf1653e7ba5e8c3b8dd14cced43d6768eeb1f357fbc666e404a70b89de5044633ccd085cd17b0b854bed3965021be5f4732fa3807b40f67cece5d09a2b1b3e509cf18d84259177a08dfd98e9e9a40084fd27c7957298be38bcdfddfaea39279c742b062;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ffd19eaa6d5822d9e191778cccb4dbdfd6fd93d9dfe529d4f8a884e1bf175596fd465bc754be66a142888fbd699d776647b8729827631733519f1b508ef27686748d158e0d7c4d986720a91f316a6167ce47b2e3d261ae623426643d551d2c3512e339fdf973c2f9af0d264f2ce3ca41306e282202a5f0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6505bcfcc6b18dec31df8a12b68fb8e896ad6d9c061bc1430550e870523bfe552e1af7f5d89525c73f86ea325fec61d00542347332f5517b49337151b66cf9a28e82d570b914c2cc4a7175e136fe443cc561483de8382ee392c66b04a9615819c41193169946f17a635a0632936088ddad3412e0ef4e022f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc650266cf4798b59ed4c0e0fc39c16cd299966121e0fb84e52f46563918bc14388bdd6ee2c359795624c9e58a699a376d0d7e3f8ca42f467c83475f819f3cd6bcc8861c5a157d2561ef5ccaa17f20e6629617b73e3129e77bebfba80a7cc5e914ef0d3a55b783dd2b02c3d5b296ee5124945c0d5e8187d28;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f502b9635e57554048181535e83d47a7f91e0914bdb99974d8463e02d026d85cdff65364c48cb0a765835abc58b19ac229d24bab844c9407cff7e4d228eac6691f9b9b4ac1641d62643871c25f0adff799da9aa2fbfc66138fb6f246c6f47ae171a66a247b73cc066cfd107ec3fcf77cf87a189273fbb2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h119234745c3058e7b4b8afa33555e4b199a3398c0f9dd7f24b3b2df3c6a86e12b9e7b1e19fb1768b964d193f7330cbf9057888e998cce3251691d1be8cba85840476db61276ae10a98eb222d5ca6a00638b728338ae1828111bc1004fe45a3576636f800b2929aeccfc4c35c8f6652cdf9f709a49f4d79d7e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h556be9f468034ce6248f0a66b82ba373aebfd156d4ed91335a02fa52731857b81f75855391f8ba2a82f8019e1caa3644f2ea1c635a06012d5f8ae6c0d63a757f5a9be5c18bf08a89f328bdb9302310371fd7fec3778a4becaf7cae14dcc57b45a055af776b8bf3a9089bebb5a95cd7ee59afa20533146770;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6317aec0dcef040539baa43013b6525418fa03f100ffb61ad79c073adaca5638ccad5b72f82142a65ea9ad51d795ffcf9d489bd5aa90cb3673542ccd32b68dc6e677e672dfcb3f6f267ab1773e852e93525f0db0a2f2f66cad102442e4573d8d94b06bb95dfc67337b9d43e2b3a1c65222308b2eb030646b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115463aece37390acb22499413d628bae24fa4c04d2b781c248788dd524e893ac242b7e8ba8b1006b59a49229bdad3e8b37bf15ecaaa6290506eb945c4d281c5ed87e9aaa4d3c832d5ef7dc66a82ad85efbf623365be3e4893f5d1e3c0afe946635aa91c00754d831d3d24f6c38038e832ea05c0b2c21ad6a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c1a97184d7cf9f1ac5d3824f8dc9c24a7ac51e8603da03a4f304105e96904e42c341da9a768bf0c631f8aadab53fe704d5445ef1d47b812f506f93d3d6d0a592098872cc00e85155d61c802014852e40270d97249b51d7e0678dcd8fdb2a14269ab34b78081eab1b7a1f992bd9f4174b7b0a186880db05fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h46ece8e4801b941178b21c74959d1f6956645a8af34c2e8f7b699a1a8d6fd426cbe19ba98ee54bf4836d263f810256bedef60e24b697ab2f78d5fedfa477d3595abbad0d889a1306df56bcc99b7c07d23afab42a4b404237bd3527df6fbb3eabee0970b2906f50778a109b5ed3a777520c99c97820583881;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d3914b8c3f4b4cddac9584a78b0cd2fa1feb13a1907a9419d3e807c8644f20b8a33afbc05e8d19a86e6775e901ed6eb4579e6b10e5994f54b3bcb8bf51f4ea5cd5cc807fc7610cbfa9adf85da03c749bf93c6bc6bf2416d287b56455141c480db163dc77c0b26802478a8b9ef87ffe7c365b500fad8494f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6bb38fc49aa374cff5b9a142ae8efcda43b083282899f73ec4835de717f03097bc4270637e54cb4ec11a2ed4a0c9856a8ab051902964279b458dfba1888bb6cf2ca6deb1326522dcdd0441deea2f2eb55d09f933adc5bf16ff8c965f41524054a3d56bc62beb8a122b5dbd32bac4e2679673e23085a2afa7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae8b871b76d64ea29cef896059eb6a77bd308346da69179ba907e73c24ce3bf1be22fd0d0c4f0866a301e03a34958e3178f1b0e47a61c6162487f832c89f8c2384fa6021c792bbb3d9629f3e1e6e261aad4d1b3d2175161572da908a4e4adf57310a791650314171a19d11d3125cef8d2599afd715b8baed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h417e9c9c345d6132735a7cee1363d28d99cc8eea39f6ad1d32d2543d5fd532bfe0e457e4889120e5c4cf2c15bda65ef66be3788e0e1f89bcbda2c0b0df46462db85016ebba5b8bccd9694cec5ea2faac3e8a1a73e4978df79658d5bbe38c25ba3ed9def60ae9ea297dfe0ccaf1c72b8dd11d6216ff55c75e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13d77499d49e5e67d3c365e2d9f659953aae5e871ce0052a03aa1dd07133ed9f8ab600423432d828885f49c016c74728afbf3754c3182420980639fc879425933ea3f049d9f60eec5788553386f660a0a7551dcf6f8fe772971962b06e41fdabdef7231ab320f1a50d6dc5705e8526cc1067065977c47847b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15071f6a056b8546471e80c224ab0df56a254db8733e15cf0011a42f81c9522aa323195db38ea6e59974acdf26538e93f994d88d0947502866ae7a517fbca5ce879f30469f085d1954a66bcdf715a9ea088d6810373f527a5826d5aeb27f6341cdcb1072951943833892471487558f3c5b8de4652f46db3a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4fa829d0e4adcedab425bd2d37fc8bea8b2fddd6ec16ca95cc239c20bfd69e5b9f4e65b9194db4d43f19db17fba6437e1f641ac8ed649037919b74285f5ebb70cff0fc5090ac03cda37df0af72017741456cfb675d7b4ca462aeb7d3552a74d3c87d97cfe0e7682b193a3abc9f09a8512e273bd5b855bb2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f53e751cf427a8ebc4b835192247a4fc12afced16a3200eb3c4fe30c7fa8f1289a1111b6a615e0afde9bcdc44d7bf72003eaf74d299b962fb06d2eee2ec8b90dca66291a0899ae10919a9d445ed380fb5e7527705d1f6f15873c6f8d07c1a8d6f58dd62467dba6ef32686f1d1592f9f142bdc8d2f517285;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h183ed7984d96e2e71443703087a20bd7570b142347aee6e47101cda6e60ce2e7cfcf6965b8479998c87fc5f45bd52fa9bd229e27cc062fe276d5a404b8dff02b36667ddd659211cc892de93411d3f58ccc3d2129aa52d84a4fb1a021bf708d46b5ca6d5306293edb6c49e122d40f458c5ab5fe13dd88b9355;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1962713a8d051c508feff4b3d37ea36467f6e90e9293b0b9a92288bc12506a3c64bda6e9534164ffda6d8c8c99572ad67588667394d1599f79a0046d56ebd82df7b0ac7bf80a0d3ef780a8f311ff27fb196a6039c69898ca1760bc0f59862bf14472b924883fa489b253f5b784ab49d3b0a69d9017077af9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b07edc8464482841361efb31e10380a7fb066961634876a78d5d413e2947cdacb4e28e61bbab5200ff95beb5f9da811c258e5594e3c95c4e5849adc4492e89d949f39abdcc25956337bfc97b3d7956941e73b09e86eacb20b57f79f2f5d635c61586797df35243e2b2ca3a34a1f25f31f38093a0fd22679;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bfd886743f81e02c22fbd67675405e7581e12adec304db924d66e03e8e33fcc8034210d72d09e3fc2fd966e74dae6a79c2d1ed87b30112a1e5f615bf4ad3efb512f5fc32d0c145b92ee44f1b722669ead5aa540ca8ab3eca7d853b4297a38ae80ddbfcb427bebc66e75f54b10fb346627bd3814f5f2d5f8a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd6657b0af8cd56c37678aae4668aacb8c62378f3009c0540912ca40cd0f80b8507985470faf651100aa169a5d067e38e620906b4a157df8c1e5c4df31f0d8671816d812fbc5d9c316562336b84a5090610e5ca58e7f447363d7290db24975964cb6a51d593ba1a4067a0eb5d7a36295a86c210e897dfde2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2aeaa154c6ab413c39aa52b49b2b6d83957fa67c0164720f22bd8dc7221815e0c404bf6d394c9439821f5bb349a97766c1cc95cff11b16de49f10d51a89b09c63fc5c1cf5ba1dcd1e4780e57670b65c218f1f1faf49da16691eacbe685010369f6f6392709c312aa6e89383ae7da6c180355aaa9f3f72483;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h95688dcb1fe81200e062f5df3ede9b02f0594607695dc67f57e5b91899d1a346c5236ba47de08d0eb35a3837d6dc03e2b1bc212ab107476415dba14ce41a0a8b17c2075183156440fe1555ea115d026e8b28a4680a3ee81d3896e2516d0cf0891b4a70e93013f63c9a4ea21a2f9f12db582b1ae7b4fa0856;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10b0244516832e27a9cc449bdfec215f00661bebb86048ae69d4232e36e24927b2bcecf593eb0120f9932c7bcd22b58660bf51560132650743c7ae3f5dde1d2d320e2bc834389e693a608d54e6819a249d2e46af8c888ef72c3e82b37840f9f930badbf391aff9cf8e818fbb986bf336560a89d9a9907c637;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he3e563b54f4ba5774925ac49a383f6dfef9a052fb761ad9b4fba10228cd527288454c1c33661b2524ac73d87cb8b8554e60cf01f9226f3add782b619e700111c3d0453d6a1f5d766183680c7bd6d883b22c2c7e43e1045ab831df802a2bea59c09deb1d8ee87937e7ebdb2b080c4a779ae604dc3a042a34a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1614fc16f85371cee50241d6b6a32771becc4b2b9509cf9c8bf4e10fee5ac3823a166ad3e94085a6f4fec83f5d175161a56fcca36f2ed0d6c0a6845ae19dad06a923e656604ea44abd6af2aa3c93efbe21afe8c4a3c38ec3e846a21e642d7c465846d7390879dd36de570d3f0a8c1cbf8c1314ef7b31120ec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e0a90fc20ceec1428aaf4df8015fd175a0f16b8e561b4466c577657610268f0052d296633492f2d96e266fbc18a968b598fd8f0823670b10125527ee65ad8edf333ce5de1f2e741c50add8f00c3dcdf4ddc4737d03305b076ea0fb9cf8b56b689a8e20958c6229c4b2fa6bb9a4f1f884fff92fb7a5e40ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heade0913089bdf3af99613ffadbdc6e195ef038ddfe47c314003356cca57e966ea4140dd69d3fbf340fef8eb374bfcc0d94a8e948b9a917d1a25efc5bbd44fb2cb5e03aa8aca3b8999587b19b3f8c5a3ac9204be79444e1e2b86eec8ef43ed314804ac60b8c37d35e369fa2429b733610a65b425ce7da5da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h160bc3e1761c2025c6cca07e715e413262577a578f765ad7c69796c20525f9cc9d17684b99402ad591b061f7aeb76422d70bbb0f65882ee9e1a9e28810fa0d2fc20836cdf6c9d91e71127ce9f6cc92c20d32c852adf70180acdf0072bb2ebc281f4330b8d37eff4f07f896d0f96b58ddfbcd210be815a1e34;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbbbc7f9eb8922ce6b65fbcb86c3720bac012794bacaff6e43b9faf5e1f91a4fcc3a714589f8f6eedf53354b4f4d76b84f555004579423c25e46ca407f6925d1f7456dc8d10b14adc2240f896bd8edb5549da980436166576e62dee6829c04d8363b2e211eeebbd0810d480273704a50a213579a548f5434b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10dc85294dd9f39e88b342e36118c3c3da0dd90a7cfd1c674927f4381e355fb96a3ffd32cddd69b6aea44591237f518d8accaafa6e2f97dc8e3966cf37eefaa1be5efa71bfd4d57f11f1c7fc8997109cd7cfe77c8e8ffb92b6a683dbd0358e687f29d473e37eb076fa50850cd4e15e36a21b034cef3c25c31;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb87f91fdbdc1535ba263c0e9299bea11936ef3d1b15a71c1cc9f9b020b842fcd1a0fa2b23a0e0b1499d1b8cae980d80faf767713576f3a4427a1a3db669ae3d3f07742e599bed1ce7c6954e86d09a1c79ec2254f92b06beb65d727591516b76288e01ddeefd300aad92baa6a83cf93432d3b68571e390569;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17013a0112cbe2c142c224facca73db951816b4f54a5467622128485d92e37c5dd1db85f911dcb112d9671a233bb109122ee728b7e153a08fc2b40d559428d04e2e702da6b81a3fbf1db4d497ca84f8fdf8d3821c22e0cc3d7e35f02d690426379d02f23c2a3b1261eddb1ab9c5d151be8596b6a8212f8ba8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12c11c75b5439c4af4fc346ca65fc7b751a46aacdd81e6c6c674f28992f9aa4f50eea3aea2232004037170d68710c000ad3923c0a2c760fb909cdfdaef0c3aedf2b011364ec8c19320aa6c343cbbfcb0a9867394a175910bfc1865190c9793f41a1b196958562cf9079d8c4015d8f07d17ba79e74c54fb178;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfcb8e068acea222476c341950161b325034226832444c9735fbd66d16e8da685474f934a23311f5c9b477880fc9b2c6522fd8210afb7f07d0fd5ca665e2fcb09910230697b8898ec6fb047e5bd74a566738728f03207525fbf44c757fb1ec4b62ae59353d6def00478042e0f1d7448d7196e773b8251d8f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h926187b3cb084e7453879145b10a6979b5d53aef2abf36012daeb8e20a7c560e059c8964a9b6d90165758609d5bfb7bcd491b4c1b1e0569e327c2dbfc1e0b68e004f9329b31ecc338b81777a4285b6572e0fe2b7bd5585984ba07b9c76f37b924e02658ca3b31be39c54c430bbb7c40b223c19df7a3e4d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7ae602942f5c6bdaed072be7094e5e6af5fae6cace2be7033200739818d62950a3342c174d70593a6d36263829ed3484730dd2055919315e5c7bcd310d4eb389962bdcc0359f5e9ddff7c8081958fea3cccb7855c3f516de035acf0fac97fbec10d71359e14175eed3065f132cf838275f972c6d6072dbc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a4361edc2b2b54f9067a2022ab6e9942288282858a20699f253b55354bc8f45e5bcc24064dbffec23533e6a61c4f9f76d547ba1fec76a9e03dc626563a0f110a8a620ae36d0f1d5510bf0b7f77c91025ce4b09133a1120eac7df0af17751b96db2f498160604881e1c681a828222c8490d66e2b464a2abb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7031de7e6cf4dd19145afd190a85a3aa59ba4efd61a4cf6dacfc48b7b520d542ad2989b2d9bece44a4c514f045141990e4317993291bf99ba6b2d9516f3e53ab28d98eb863513acc72ec90f17245b4d170bd7ff0eeeb45c2d14845c681a116dd0f8bd8b355b00d0e989cbfa5616f44df8094ee5d1863f61f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2d4df28e8e6343a67f7033c0193fc1a6e8951b1f85b683916a9069c028a0b372aef1861f7a1f8877c8b1daea5c17aa11188fc144eac8fa0e7af9123806059e898162d395193c13a2898c07c0c43d8e552d641302de23c13393971e1ad0f72834c76b1a162367cc5cd7ef37999e09a903b9d125fc7a9b02b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63dd5ac2bca9684133da413f0fe8c2c358c90d0cc6cb3c3e527df4a312260612eaba8e6fcfd6fdc05f4d79aaeab54d1c5393d7409d920aa57c16dffefbc0c1214fb48f887999c216f6a426b60fdfe9e9723d5168ef05ac4b26e5442de5039722d776a88ab1940dd7bc9526da7e14af0a1e4ca67c28d28ff5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h163edce1663970cc34c1c1929d33d8290b554b477e7f554f0229bc446cac9b9e1c64980c727215a71a2572cd6a2100efbaf14c90b5976d2a84c3d0c9671aaeb25923b5d3f12a1ff152786c12e7a0f3415910e5cbdd73d879577e631133363a393462207f387fc8e726660e13870a71425344eb5c938672c52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h56ae2d3859d64bc7a12a02bb0a586dd7465e74e6d749e3ae2e52bf54bd66c5bda5acd770b4e95ff258815985effa4e08a3f565f40d0631388efd6396b47699b55faef9f29a6423a421f63bf5402d533dcdd6dcfd6314ff0c06fa9b4d6b12ba9576590221e158e90b40f153e12beb8650ae425099ef1e6174;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h995dc0f452e6f9b0c6861acd5d18a397b6d2772e749e90bd395995f675668c386730814dab38a137760622f0dfc1b9faddee608815aaea6d425de2d74f364b32ae81914f568a80984d86c4d4ec4e8239e7efe1f53d9c020cf2e510fd11fecd8524f8d2bdaa1994e22ab1a3264348a374c1a5ccb20b73723;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e3fa4e35bd65a6a4f8c9969df766ed4a28484036c7ece53b275ed2b9c9b9d988ab9aac47b9180ef6706583f171ab7239840f2ced7401e557f43193cb0e512e16ad8d2bd7460f68faee57cc19c3ba2339b4080a3a79405af72fc0cddcb65f240f69e053de3b074457eb26f455353c3563ba0f746529544b41;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14c18de5068c03153139fdd929730482e6d4d55f95c54ebd5d0673da4b59696834bccd012668bd8c9f12b87f78382decdba6388958a8f970fdb76174af5f8134dc0602e7f74551ecb12201718a895d67b535b75f56e70617f5dd5eed137898f2c269b286d1a56781fa428e994abed97d21f72d6f1a27dcf25;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6466f996f8945b745cd9e00da48ef0bab20e00534159afb11b914a339b83544b921ad22dcd35242c0084538de4cc21c7bcd1062057d85f6fc3e7c68312f8660f5fbb9fb5fad5189904fa4b10b91060b73c859af1f221268c49a1848e365188770a020704a6de9acd82d7c6c6e8e2d719709f36f410572e09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heb04d19a788f4c3c0438e1ff5a8dd1c5a94728226dcabf9f8095f4bda5de626b4df40cdd54109aa5be8349e096a8626aad277f7bd894616988fc7f0f8482fe39f5aac223212befe1baaecf4d1268dea30019db366152af8545b3fe1afe5f2c3e927200cfa4e405e2a7aea155cb410f22c2ae6817ca452354;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2b112c0206c89dc03cd885a090a5113cd1621c0324cc4c0e5709d785afcdec309e0b04ddbaec1d737cc39290ba847dd2359710fa81370fa50f298cc49efd52c177f4fc49bb0f36b944aee2c60db753b674800aa4f7dc4ad45e4787bb460b43a34566e8cf24e0ff839a7e70bedba5c5b704de00b9c31e8fd3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ccde9bd5bc11e2770b5b25ad1ed32781944a758dc582ab4bc3031fdd6164eef0d541fa94f90913335ff619f1c590f42c0f5d0dfe506fb5e85af38f3083c52dadff104c66d50daf4376b0e9b0d98c3ac150ef323a2454a0bc5457d1082cca97b8b161dad1d2f23693ba4622d8bfb2946cd7c2dfa9ab9ae05e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bae7393ede78f247858ce9c74175887c533aff5bf7e6c8e21d389ca0a56b1a3a9faa33e82254867b0b2309a37faea93376a61cbbb32cc36782ac72e9a2d9205e8546503f09ca4f6e9d0559b87c5696584bac91d01fa71510a4cccaa24faf0871093b11cddf9781c78c4cfcccb2e0c704e80e7f134039190;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7bdad6a6eb3c1e92e725b29a398d7b5b33e8ef6e467519bc886af1058306579e74bf3ce18796efc1d67d2b61311e86ebdbfea1edbf84d26940519f1ce9b13a9d9dc33f0dfca84dcd20fbb3c8a33a79d66b759050390cfe6cbd9ab0c7302a918ef9aca983353ba9724118426eed557ccc10249bf5e4b9d997;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117213368f178d96abb3a2d587b8e05be3d9a50d0e9ef60ffe886e6af0a9dea2b06c88fff087de9630b953b9b26e576831832789125646f7d1a39434fc0c2d5ef2bdf28a434c9043cc77cb830c2de476109e718b8747349a2f1cdd6e82b8bffd689b315854aaef2745a8c33a0e1a9ef2bf299039f2526ecf4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f427c577adef82cf81610c6006bebf96c867b71c5f6fdd87d63ff0e897c6f0d8ec084d95d9d34fe57441ec358dd1c33331504c56b952c2d76978b673d7aecb039e9f501355236803019dd7accf2252f294c78a558fa6b0f98018615249d3307c332ba09269914a50d34d62655b2d9b9ffefb0e95dc65e81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf262d1919bb0339b01c10a1c9fbbbda41048c4062185ffa62cbf4030332c4f96cd618b1a8537b2dd11b81aed68be0b65ca1f89d8723ca30ea04eb7988f7485d705ee0d19448b4e86c878f74f050e02fa4de80ddc6caf95699e1131a61629eb8f5e651eb449ae503a6b2ab7854ab3ebcb82d020f4035c1da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4fd70dfa058423b75e03a6ffc8b449dc529737806ddfa4c5f398b00446ac1b9c3a0b4dff03fdf4940a8ab30ab2aeca3886d23d40cd418f25d2f205ac42e474e169f6884ab5cb7c9f634036247bde2e49ad1d06f5f4f3786a9d10d1af835ff96b9ceccc9b389113964a59c779283ebed853876e12cccaf2ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h93248f1ee246095340344de7f0d53071ac96f7df097abc4c2083a3178525139c8064ee8d0cb167777367f62db70df129a366b01699fa8006749c4510b0edb52089c7eb69005f15dbe30b245f2b9dbee3b2c48173e591332f30b5359e82ff8a0b563d5b2bf4dc562e8b9bde174a4749e3927674bd00b5a270;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b07393ec25dd710fa9e4bd2ee0119712e7aa6565fa4e6d1731bb69ee908009c769dc128553bbd0c4f355492724eb73dd3cd54997ffadc74899060af8905c71b4d451d5d54b493e91b5aed1609018a56ffe83e73342f653b9f7d13a89d5ed2c68978e4e6395568afe59fcfbd31ca1aa18c1bb1522e25221c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e30c5047bce8e96657ac407f77c0122f9b566d09ba231e8c7936c9bfffdcb8059c16db0fa420a54fb173ed1706decf0d2c15215e06e972e76795b749387cad3982d09fe1a34c622863d8c66e73751443b38b816d6e381787ea738bbc67f21f832c0367d6b0bb92c8564a4585d18f734f435c59f4dced53;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d75e1d21a1510f026324fdb2a712aea71d5797096e948fd126b6aaceac845e1fae3aa4f95abcd330d833fb0a23b0f209a5240920b9db227e749806503d45342b1014a5c6fde2479cdd1862f970904e1f85099f845837413320d53ce731d777cd193780df49c56ba8eb6926018f0632bb5da02db1db6bace0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ec700f2141a36dba68d77e09d39f0a5473ff880dcb30442e28456da0d0b67ce12d3d6bc93bfd1a0917291cc21a082651df06910d499eb8a16732a8aa3b4af00c7fdff3eb1f9d8733a39d09a081b1f369f89c5f02f72d5f66dd2f32e77cd3c0a1cef1f57b88f0cd006a52146976663a6c8e95044988b6b26;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e35068133e7a6e8dea953c15e32b85b743ec284288ba09acee522855cf86850d3ce8950e2ed21929e49fee4305f969ad065a33e9888087706f78ee6ff2d58b96fc1657e185e20edb3cc485f02d0cd66c395c0d7018ec058a8ac2aea03f90f3a6db0a220ac624dbff4c34b2fd621b4c51e4265dc13be8dd1b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12c8d5452201387470cbe0a5370dfe13e4f2f591a841b4583691f9362ec2d6cd1e93f4674c1abaf458daa140d1d9e172de66d0c90d31a300f7d503120d198bb7b93db75f7ae4f3928d1154258230e0442fecb5ca637cf6a26d1fda7698a8b7c18a9728a37c8008fbdf8c54fe06fadb47507c132481071930e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de57bc2ece11d35708fd5dff9fa31bbea412de705608cc8fa420a4a83d08e5f6afc85d52fff6021d2af1e97816341b07cf6f0f35c4724643713f421f11cdd907e8955cbe19d1e0e1ef8e52a028835cce39819256eb49049d8826a0c9db5b664332363932378c9795d35bbfaa75526502eb0dacd532c2150b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13947d45fad30c7fc931f514688ef836c70c9c616d21a1b5c166d29af764446aee34c679a1c3c923563cb3e80e90e9da64b0d089f65aa08d9c1e03b8b4b56053b443b59d656bd5c0c3294672b67fc1dd0b297909766068335c01a36311ebf528d3999177de660ff32422ddbb3973baee7ecefcbcb67c0cb2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h135a04e6440598ed1124713e4b741ff3399aa925a5585a6a2281a7f9ca927b9f23725bf8b6897dd55ab41d606bb707772452e6529992c6385a0ca10ed77b24a2d20a4444ae3dfba8eb491cbc44f538c0986ea8b0daf07e58a7461e55054b8d1419d1b92e02a52a83657dc7d9fe22e7f0a1452cddf4c7c7306;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34fe6ea7db4ecdb0b20e3f02bc56c1aca4e9a6ee873b8d6bfbf59a078b2978c83047fa40bd3ffc57af54577046fb7629b714ce80bae906685ca9e2b6b664c743c0d48b68b52482ac594ad7d7e9eb22db409dcc226bbede18b1907a165e04eecaef52a296526d0e0866b5155d73d1643e7d580bf25dcf375c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17e6505c7d41339681600500263befe2ab5f69dba18dd25ac87a97ff6711f421c2e3f10b8729683609f0c5eacf0cda1b3f49232dd58acea5527b5ca0c7194d92c46903ed0739761a25f3edbfc9a20700e5e944c5a306c5231dccf7abece90cb3b2c30d12a0c12e71749fce79eab0fa72b7bdcd41823c43001;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6adef15a3ea91777d429d0f2c7ec193d2f856745eb10e6b78fe00e1ef93b5cb7c148d9fcfb7ffceeb3305e5decd56b3d5994ebfac1b9debea3228e637113fecde9dcb73b07e0804dab97f89331f1414f083e08d7f60fa572626011c07be5b6a6677d149de3ad30714d54cafb5bd770a4f3fb630f9f2bcb65;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb35d94a1b7e33b5ac4f93df835fb05ecf164a731ac67b68ab57c22ce68f8b7509861511739b59e0e1537e24c1bff54324072277fd59669147cc73578fd86722fa52e966b076a7ff43cab1b3856c04243b2c67fede95fafbadae3129688b3a26f8bc1df52f9e4a8e6d7d99bb4d4411b6eda36e7f7941e60c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h145c92b3acf59e4012d30c7e9357fa2a09b3f15dee31a8abe86b44501e91eac121ecc40598a485aa164a62b43c6b5a2a8ecc5aeaa0d1c37ae418e1b1fa869b47c64180e4d0408eeaf6d8b1b49d3f396b3b2806a2d1593333cfe2fdbfd1964df47e1bf990727bd459df41a3d049800783c4e639cf8229c9697;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb758e160e1755319bfcd9ed4577ff16d193c2887f97f6f41ca0fff6906a7c515ed701064b92770cf1b7cbaf7965f72d13d11fce417640a700c74b4daea51eee11c509cb792b5f60a0952c84a905addc186fc8e37f955899481b3b3d6f6bd4005c2b2f5e362e54ffa53159325319dc7cb841a47aae1c5d46f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5677964e8ba85c7e9b81cf17669d5ecc1ea562541664f67ab4ab37efedfcff26f621ed7130f83f0fe5050064d96b1d68e8906de22158633b6ed7c99245ef697164ca54bec70bfe00147af45477f638e182ec53ccb06ebac2f7dfbaeebfb45abeaa34653abe49a38d243297e381a997eab40c63d607219f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h171eb8bacfc952f609833b620ca6e8dce9a6d459bc97026db41c8e9c7275f472167cf08760541987f803ac2354995d6a28d5e3af24df70042ba03b9f83005c656c5433dc7e473c2f60e4ee9634f7ea92aac07e9383fee2fce5da87de7afacdf7e3922fb549801d1d0c9be52e638c83778a54dd2fe3773575;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cbf44b1a5703e2a424712f8519289f7167631880c1383cf5e63688915e9b4f31eb84226fdc956f2f40ad44823a3c32edf6d4fb0d70090ddc08e3f384ada52c1ccda0e023f16f43a49aae9a280398c794f1e43ac94c7c906dffe6cc441f8686cc09de20b127c2859a580531988059741e73c142cc7e775ca4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h856c978014e01b6c315f6ceca5a9db5d89f796171bfab3fa21a39f1900373d11b3a04a5945b0d47232a0dea5d174fff170bbd926b0e2e180ccc9d91f2b571b9147bd6d49ab3ee9c004352952db7dd753a809cf55ffac1dccb743ebe8074c0b78a4ce82c55719073c2b5c41a5eac4b130a58735a3f4f4626a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc06d276b079d3b6ccc96130c109c816ad568115510464d385f553f973399ec7c4c0cb0fb80cbdfeacbebbc95bbb16395a7cddd8b4f7cbda39955d6ef0e52425431629af367beaa08add3d35d509d1517ff7d92411f5da68b6091f0a962e79bc319b3b435d13bf92c8aa1b6376b77c79c99b4ae047b1b357d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h178b1d7e8c7e9edf0cc2e94fa707f37ddf44a5e0cf95368f598e1a971926a6562fb9354a7ea372e6376417274bc417d62d472333027ef5d396c9bb3ace6a4e77da4ac2b424cb384f82269ca20f4a7535c91aa61e76ace329f097bec4708b3135c97a0fba422d045a4f37737f708d8cbd47c028982a3e6c139;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h72eb2a31dd9997ee2849ccee5b55784c6baa70bb1a65e1b770ff049fcdaa09e2f845f91bbbe0677f765aadd0f0b606ef859315746756070b42defd12dab3f01f2debf3693afbffc0e8ad4382a3a38c577cf28cedcd8d67378f157575b2d98578f25a574ceeb492812dc0fa8febe1bc7e2aa8eed9f33ed2d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f9321dd66816436630a5ec2cfcc90e0407b6658ace4b575e56207620f55f81f10befb77a89071626d6ecb72aa564346f0e24bcc62f4d69bcb1c2675871e612fc28816fe4f4256d54da48764eac018b27c915f227c6009e46b3ab7b43490fe4c4b3473282e328ca2a78e9385f0d40b2c93ce6cf01f1996e97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h74538e3676dd01951f1899124b415490c758f8ce211d1e3f3e767a35a514f0d37db54cd2d8c62a737caa4f976192a16abf58d031a10abc4155c54f10866ecc19ba42d5700ce687a2b716c3ca5f91f4b76c267d6377d91b09c138a3a78ef8bb77b2fd1372f1749235a76575f3f6d02673824288d008645a35;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb31d71720dd72c4e0537b0410039edd6d3618e495a2a0c9d659f26ffa28a8eb9c959814981e1336050446f89b19831d062439236970a5000320355b2b5a3a5a4f7ff81294a1cecc3747147fcb0c34b8a5c43cc6141a9ac2b482785b30532cbcb41c5f1d4dfba8c1bbb9f196d9c3a5c484c7a0e109ec36ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2fb23589421d47e48fd3f1c6e79f44c738e666667060cb586f2be9688b1d454fb0ad4578d61aecc125bd90130bc3007ccf65889b78fa22a518e6586b5a544db6ee4175ac75b9a282e377fccdd763caaf9591d9d5f002686e007bc4148be0e0c3896804d080052b50d0c3290eedcef57bc72313fcdf4666f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcde7159a41ca0771bc77b654e5b6f23db294eb25c776a4abda2378e11879f00b64bb34ef2739dad459676e41c0634d0bc55398d97afc886feb079d56ef1f5785ca92f3ed8dab11ef7bcd3d390c109285c6fd9170651adc5e7fd403c6b509d33f6c3a4cc1585c9d1d29577d7803514eddf5475137c222dc74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168d2a40967dc80904566981b3605261c3b600b9762dfdfb78ba82093a5b3b6dca1ea3bd05913e90e78c0bc7f9fa0001d4d022fd4906e726087b9189432c5001e23d10434d5c70fe58b9efeee6e8fc9187786bdab1e40d02a5be1f2c0cda1e867392d1f91b14396a67cbb82a0d42eb80270fce6f8afd88f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a69b9ac2e3e471ec4128c01c926ee7e487a534d34390e3a2a28a719e94e5419637e654713713154e5b201e665980ec271f4693e1b180c75f66d7e5e1862361fb5c311190b65b1f70b2f4674506eb9b1e866d566da195eb324e7a2449342ba60172ff641f34dfdb8998c27e52855e74a5f46a23ae616a0f50;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h119338b08bc3d1d48fc817aab48d59cb25fdea420e37af67b54a8b5670489639aaf7b756178f57435e7377c2540bf15a942f1129ecd5f1cc66160fbdc2eaa1badea341d44ba89bc6459efe2ee7f5f885c400b3a92cb8dfdf2f2bd24a2443b043ffbe8cb7f9890bc525504854f9e37471800013b9aa1ae3625;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1793d567f6904c61413dddb237421e975999edd0c8714c86619e7a18eff3716f3d12677730b374c1308e23816cd8502bcc089767b55d807364c612f74da24705ec383cdb7a83507825dab661a70a6f6d042a32d2433dd7f74898b1abe0ae3b144bb6c8b82faefb5fc67d322a0619bbd470a47af139c99f2c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h43b2eacf1cc34056b203e2652b7fcacb8188838841e94106235127207e4fd128d49f11713e40b733e5b875887a5e83e5cd163f2b785e43c69dd27c1fb6b285b48e03723eba360fee79f2cb4d79c0e06756cb984512040dc520b83829222c458723fd63e83155fc513913a637932e408238c5090d19c7e92a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he2fb0ff70dbe7b26bcd863fffb7f466ac5daab233e58fa991c8759e74a8b50b12563fe05aac6f49d063436af4a213f02559f14fddacf21e956373c26be2094d1f296ed45ea8b0dd1bdd1bc14478b47359b2234d05d69a793f2079ed963fc3b8146a93bf7b2212bb7aabddf48c29a7b9974d72bd58257f8bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5f7165f025660fa9788ceb4a61412bd8705ea6432999d03adb58a2c212250a99ee0cedd307e3f7073ea38d16beaa1d9e7e82601eea6fbe81bb178bd48745119f5230366e7728c7a3877d8ab022f7c4ccf098ba75d614152fb5ecd54ed2ff75ad3ba87a3482db88b39a7627ee5a6ebe3fbdfba06d9536c7ce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1569df685d345b9b5d1be77cdb0d630ee790d23055cc56572a85ef13ff0aba7328f25e7aea657832b5eb00610833fb3a26ef65b4d93f96a9cfeb1b83112362fa113bf24ae215c11751525a62ea633f62ac5c1160210041f32e190b031604ddedc43c709a4cda12d3e35674d171b8d1406902701ea60c24619;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf33e61b559ec5055c608a3cd62e68949597d7db83caca44f1ca68fce03215059027709353d8672994eae6d6a71bcbec8469386cab3151c30030e5131ae7a98ccd2fef95ccd439eee845173e3db56267dcbce8a08c7eeaf972dfaa396ca516d31e2aa09a2a9c35570b8a13cf15b425030c09a6d438b523d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5c808b03f83958010f04394c3f52f29b81ddd56793d2817df8775bb6eddb5efed6aa86fd91c0cab64e0456e78b56381ed100a403208e4ac1d47242bc1182644967ae592f0a7ae2823052ff68f3cb93197f9af9931f5a055ac554fbc29f3680a64f9c5eac14d730c9d4c6d6bfef9fd0a4005345d97614ba8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc88de9735f3d80be0bf2e6082da6780f224b69fcd2edcd77be24376b888b533ab5a6d1e7dd1e04d6c4abb45739275bfd1d49b139f79cea2821f47a41963ecbbf5ec1323c2e15e54a23bb327b016d2b03880dc4b2348b274f193125fe2bd83f43f48ba47667a2ee2d17fda18d2588ceacbd13a15b85f06d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h321847dac7b7ac187b0194914e9fa81854565312120c4d42c37f5f010ab6c104785d3b4ce8f80b49485123134fb0b3ca9c9d7e5c063c1ad048087137409425d0c67e3e0570c7dbb1b7c4cafbc72bf080613508492191c0baddbe27e6f9adaacee4ba90bd3b88742d993bf95bb6762c2d8d2747be0d112e20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1873a61e75d23acf9bea1368f294d56aab3d3615053d69b7adb095a0b8f4c9c0598a64dfde9ac33c4775e8fef0221478a4d173e5cea492be3bd25536e9b86e90ba73d52ec4caa17e5153d60312c26fe1bb281a110567181529b34307099db8fe3ed6d303d908a218f3c287bf028b2906525813e1199c934ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h348b43f656d96addfbe3e3cfb7ee098dfa4937732ec8177498b51ccee7ab39cf2cc493d1c5148faeef9a4d44e4cabf082ee63e5461b97236836321add1ae49b1a58e857a231c0038d57914dd51f659090cc4d732d06d40a2fdb7119d65e2b55731110b1825b1dd5c3d3f60b5684c31e18fcead8e95da0170;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14aaaaab93c11e53b5e50d56a374f7dc9cc0b5ada8b599e0413ac57a46d7182f7bd7edf0be1c874a2c432de0c54292f4172210bc047aec5aa099d11d42628ef43b88c58017de3ca2bbbd6c12fe4e77b0b5d401dfd1bd2dc7056aaaa0f01da37fbd357850da19fb704db70b6a1b15b72118048ffc06be30d2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3641e917c2055d02a019734d49702b8a1676b38775af3f3d8761291810f78bc68c47e1b9ed11395506b96935b3e1981ad304292031c24d8c96e9285f43a364a563690f78e08d8eb40d016cec4cba3471ef02983e16ebfc799e9d0e5be6114965de2c800e628c71665436a6e30d7028f6b68d2d4f07b2a3c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2219cf474b60838fa591e9eab05d30b0cbcf1a19b25618d61c91f4c42ed78ce179a1fe078cdfab9f31b7d19298da464b9b475901342f7d90a164e50877d56b899d935efa4e8ae2474ced166912a48fdc4ef6c41cbbe11d2ac8e06162e0d291b79237216a6f7aa21b196f69fb7594ebdef41d6a62df03c650;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h449225925d53f2b12e3890e16ccbf7926671bb0d88d56fa997e9264609d84efa28e64f167c4959509ccc9eab18620ab039d6697fd39b09814177aa1af3ed16504850d71a03a9909c50666a550411091247e791f4e25ef7a0b35370cfbe98afc94f737ae0bc68314fbb1435baec260454d2cc24e986cac89f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1741d746e4cd77e31fa8e08d1ad60c49f3a0496b418900611569a63350f4d39635ad33d689ca312b715c1331b5291c260c8466db763f2da6bd3f56f20215cb71c5f704f89d0a57e758dbdb2a4d5d3e6b4151d922e0d288a5bbf46d7e391f2993f27f95597aca95e8c8560e45a3cb56e98b3a78bf98aaa5ebf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8eaf5f3e5d2f95b1d9db56a6d590fffdefdd401743eeee11342c2b554433fdb58f2c0047a31586e322d9459714ad3339548f36259fe6c43df0e02700b84e03c67fb7145d8bbb70a28f46c8e3478c9a4e469bef2193d5c7a41112d3546a9be3b83b268d5e5f4174f465512d70e0f070d13b84684db0e46356;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18827cf7bfc1aec827609e49d1243a4d0ae2cef39a49f8dbd14e3ae8f65a40c4c9c0d303c40142f8f909f4f5e77f6f61994b6521e6b48150fa8e21dbc48bf37b3bcd951c8aabc9e20a51a9dd38dbc8cf39e328dc8c50e7b652d623ca6a5b8bb2e5e288b49b58ed5ec228810abf09f44e687562d26b2bd8e4d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12940732a3835808a00553e76bbdcd7b1eb3514c23e4f0b75b00d3612abcc283966ffabc511a8cd7d03d97b1b72ce6fdbc96aebf706476cdaac7a20e2d87bb89fea4bfaa56d22283485f70c5eeb71fb5a80d4acea5df8e5191dda162fa601fa5556ead081b229ab957ab491fc8226010ac2556adc1221a036;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he76cd542c69f3bd3e8c68f3d8555b33ade2e104d81b33e1e122fce22d31fb80352a31fb75c96521acb48d1deb00c58e8f47f8f408e83ecaf938fb47c52ea64540504bff9b9b70519fd32fb09a0cfff5e53b67424371fefdf99bf2592134154c2c004609184be2c89e666b2cfef1cd21da930be96903fbb7e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1928aee7fe33f184e8ea77b7d36de3836facd7e3e54e77f6b93bc8a54d1e068c1fda27222ced0b41397abeed2e366e3e0a7c8f56b643397ab4d1b61c8a0205bb2c457502c510484cf5f1b3db5b3e3dc9f5628bef1eb13fb1a0710f03ed6a5650ff9e9c7d56d56b68d09b35ce2482c8f1c5d171591a62e4527;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h682a50977f937b099284572ec60ec07f39719c09b02cc29221d59efdf8fe80957e3a1ee952a438832de3eeec183b296cd1c8561888f85faf5c69c38aff96981175b226d5ad81ad147f489a5e8f1d33b6a049ed928aa4b7a2e2d8c37c8386fc9c2b8a7345b2a70a3aa655b4b46a9cd95535f9011a155a573c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd64d5d1b7f6eac50f5e5938cec1bfc14007b5236892b4460ded0fdf5a220fdfdfcfe1639ce4999280cded718dd0607837a19912369c28598897e29c261bed90cd0618146dfb50627f0c179c6796ec0f9b2f37bc9bab6fbf8db814c6bc5865d53db8eeae6999f99a0640b4090b61008d7e4d93e8d565200d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf3db38dbd4ea8699c50ff50fc2dcec3c0504541cec9b00adbc8d7700be8e133bf78a9679b71564d944417d226367b94c3b0c171d1b46ddae60802eaf22f711f9280b033b971201b35288f5bd355be0d8b88846b5c50aca9051eec18d5d30bf8cfabb9eb5b8e49573cab54cca821922fc6278a6b434451a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc44183f917d31529be6888c49cb504895365d3ccaab73af5ad58ae1160a77e91bc5bfc868e24bd388b6669f4a042f821e1395f1d5dd95014331233b0f1290b9a77d6edf06956785f84cec27ceb05ddcbe228b68ebe86b892185daabaa06ce75d20651bcf3451f21a0d0a6b8bedabb43cec530a284a5dfae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dbeaf61e0948c86eb017c880b7d0d9284a46b4f7592d23b06bf9445f453a8b327810bd4fd4de00c8fc3e46d7e175d16633231d615e3f0577c5cbef5a6177dbbe3e0c1dff110e5a8aad255c2f67386e0a84fb7d77e36d826febc7014b6f8de32c28df27f92d37923a85549ae994339ab3aafcc5a6e0674838;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h528c6da4f68b6e177b0318862cc728601887e9cda12b69d3ac700b93e30a6847be16b85362103d6d215d19c2d1d53cbc3538794cf7359ed6e1f4619b06ccdb56ea1a56c09f600e47d0833db3ad58118aaede66cdcc3835f0c5cc0e9683b4445a887d7c8475a2f683bbd2f1fde9fac336c72c0b19f6808bd6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a526cd18ca6d798fc3703907aa5c72947340ce07feef03466505398c456e40d84bd5cb53635fb304133fc8a4f054eb8b62cc5d939c94a2c01edc35c3db8999f4c0b8872feaf854230a9b24e41701e3479d92eac35a56c095a7d7969da00402b88a3d7308f4a9c495e0b8558aa674a76e95d4d43d11bca62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1726bb0d6c56eddae802d30fff44e391a08979ae5ddaab6e13a34749152f0b69e8a8729e58398858163db42bd51837b2bc370c4adcacec598072a064325a7a862f14554f7b9e3f4eb4aad17672841c58acdd01e252400682d954baf980bc02e77a3bd44c9214063e884d6243bbdba64518b3643de0c12b94;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156a2ee3c253b04a714ac8c1af528eaeb17b1a9244b6b3f59c2d02f54e19bf82f05ca028430679eb113ee15e0b6052233a87df78141e9f92400a804b7f391bb24bf4c7f0854cab15cd63bb3085c341356863377f81eebc6a1281d2555be4aa572257f30d550264a3d40661081c6d5f413ecc7790fa15c8816;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f18effcbde687e7b068aa4b20f926f05a17e6f9e36318d40762b703d87e95c8a181dc35dc091203274f71d10a1a2c68b346ff4880c4236f0556adad15c1680751da3e9b973acf757fb5689fe00f8471c8f4276f67cc808bd5d1632b077b59e960d06894b587cbf0e4f92c86ff6a3b894702cec2984c2d3a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b287bd91195fafb97a0a0ea4e5623a3494830b65f01cdeaf79ba8b0d3ea829963eafedee1afc46e539f44baee70e7c66d956c7aba5c888a24d61dcd4aa913d7b8480f731df70d0ec50eac5e9f70ec54bf604845d5bf69c1aac4f8a2a1b73decb6faf9f8296723254ceeb0c3d645a8c7a58339dfd0aa89e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eb12b5c5ae87ae40b0a3656e5898fd13631a431fbfa0eaa056d00436fbe1ee351b0f4cea19aaa13410f426dc63f5ef9c470fec594b12720634461fed0ed4cb334ffe8256bc011f013e15b8fb0dd3a50a66551afd14bfdff201aa786b417d64c7082421adf0be93e76e672f28b440151dacd94480771ddaec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bbc7a7f6777e3278481b81e7278996f425d327023b3a1154282f813f6c2c9ad32d5c0acc9922d847102e2f3e887907d12458eb1d108786e1d3b2654eb527fb4b24b9596c9e59b439a1e6ecbd1f0dbe22357035fa29da40fbab2eca563d016a67ed9b99869c65c58ecb3e0e875220c3153cbc4f6b4412e827;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2d5973af39bfe0f41d2cea53f90fd089b73036fb1455f7f06ebd50028c84130df40ef4693fd369e58c566ec12b3dd97b0bbdc6adf98c8bd1155c344d1bf01ebe8343052a81bd1a6aad948f3e60d7e60d1dbf32e43f7b040109502cd766a972c4bfef7e3058d8e24b368d12d7af6dc3b79a4caf9a72ac4e8f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1997a396d26254a29f1678d7bdc9a362bb073bd93e94ecf02cc558002c44e738c264dd99ab34127cc725c1b3fb5e096c29b3898a5f6bc3c1009583c7d0aacc9e461cc2420222ddef066bd2c03342094d1710d8c51c4f97e4dbf7d5d76cc9e437aeb4b5ae359f24fdc60665469c38fd91a116f15799d4e0eb3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h466f28bef432373dd984b7898c826dc4bb7b134368d87bb81aaf011ffd51d77d8fe7c67582cd5d8ec8bc8a2cf6aa25734e522e81eb86c90fdc831f0ab6d0d731419237f7bf2117b6fd7f2832ef146c20051a1aef7c9ca2747dc1807624cccbfbab105aa129279e40d608cc159c0853cf2696e6b4e571b766;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdbcb1cf41a4dff7f0e1fef280e816afab7f42d7eaebb4d35ecdd603159f789da5f188a3e57368fdd43999d76931223ab6390c28ae892725f93ae2afd6fda458c9f6200e7144b2e2c31bad0b69d6cfbf8a7ad52d503bd10c6f421c06a3b03ab6418a9c39d3352489f2f460a3f0f66f815d5368f1694670bc7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f727fa28200ec29bf3331af97c179a0f6e2e616ae804a1767ae735cbd72ef183dcc5ac36d867747e52036cbc6821398187dd86ec68c3b5e88d3c00eeeff869526e3174c55a8246109c19ccdc1018370f7f6b623f79db056fab7a02097fd2729dac7fc30c82baf4dcdc6f782d300e333e59d39ea56f6c7153;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h138d465ee6085538fd29a7c48add23b5d6380d95e595db02222430f856384965d7fa09d23d826c2825b4f2ba70f319af17443e8c6b7c37c57b0c4d527d5754cc570318a4361df9fe3fb741a2837d089d8dbfa54abc30126ff75bdc541509523e7c28c777772bb2d0f71586e9c8faa5b6a233dd5b4beb0650c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b9ebb7b3863ee6a54f04c6985dea4fb843dbabd3cd448bedae862995885fa318618908f76e373e96b497fba756d087ade2117c4e7dee6be748a32af1ea7f8669b1ca31d5423dedc95832359df92cf5aa82dc9e3c8c0e78ba03ca5bf3cb9e2eea80d1d8cb2fce644ab8860cef6b34529ae4fc0a1a6858a5ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1f75b37170ad91ea56ba479b6855538f0882f814d46b4ed44c3d3b3d18fa721889e9fdade174539ae7c21a3c19bc80beb5c1db789491954f4d0735ec8defd0ef73044bc99eddcd1b761d72f4276ac6a9bd353708a91f0c598e62a7bf3221873d935d41ede6be8291320cb381c75e567cd2fa6022c9894b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h135c4613d8fe977237c7c4172fb306711b15fe38ec7a5d6dfcba5a3c5d9e5babb47412751a82f55220c3b6ac23208a9777afb91360b3d3a1731a3d5bf1ad9e4602abe5d7a49a53513e976358f79fc1481ba564ede6176e29e859441a8e8d50b3b566ff670297b48289766cc81690be92b2319a283a1fedac2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10b872a3889f2b31db1776c2e5938bbb0dcda3b69cb00e0d0e00224eece54ac12eed9cd70cf1a7ec8c640cd42a49c7bfb6fb7d754097c3c7861ab980edd60b173f87f960d10778a920c8d11d00a75700aa9b23381183fa61c993b138c6eabcbe895b6d863096b02b134644f126b22c3b09fda1b64801fd86f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12357820bd91fc389f39f7ed60bbd1566d6d0778464dbb2fb4a4d77d5606aa2ae0517f15f503157fbd20e66f42d7f142733e18069ca5249e859d5e5508404ac938e920626885ff0d2d089808aa3a58c9e623d6a8496cbfe940d799459ba8bc4e81c69db15436ac0ad7b6e166c7f15ac225238b544759e6e0d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1bb8b255041f6490464829742eadac68264f0cb96c9d1069b5f29b88122742cf1d0a70d89c8e62ca88c10ba3300d959955ec742a1134fa595c1654aeea680d14b554e39889c6a512865c581d0634bb24950eba2c5cfd0d11c1ca1a5144b7f6404677296d7890d4825e4540d0567ce68dd256206bbdca970;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1094a3a360383d7dcac09d3f861c5df20e24be60cf947f27a9e1e6fed13e9d5ff87e190d3cd5d1cbfa444653a2e35f6b70e0b540f105c9483809b327effdf66fbec93042a8ad45f147f3eaa1013fe5d7dd57876ff59cad44d6208bf61694647ae331b8d3428638040e9d88d70646796146a19232ed9bb9ff6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1beaa683ebf9dfd7095dc09b15bca4b5a63b72430706a16da5e2c610338f4ff1a1639253a964c2839fa20da164ddd223f00eb7abcf394176e62e7c33adc431f4c5325eeb748b11f73b91e5ee18eae33b5673d9d858b0fcfbd743798e96da84d6a99db49758e79fac7fd0e1ed1d091200e47cba31b9d0fc31e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h103ba5c46560565bca45a11139908f299b99b71a24943c27afb1cf5535d7792ef71b9bc82aed880b656d16d02d6f118bd7eaf4cdbdeb178fd228533553b2016d24b8a9d2bfd1de9781a40d9c89003a5c5d79bb9e99bf6eeacc36bfee31831f258fc2a9e3c1fe57db73a1dde9da4089cd244835e26fe28b872;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hba82cf5ccff8789df03996764d4677df811a66b957634505c7856a26865d0126d6931a1d704c6426fca8a93010e688a4eb69476ddb3823c8f0f6e9cc54a1e8b7121df844ab80abbbc68350102a2c1390c5e2ad98a1c6d1cc000b81a134882dc8f0f9a6ef19233acae106e6570b3b5992495caa79471487d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6678505b8320bec4f2bc1a4a8ae84f320ee3a258828e07868a7de36859d0d46655d074beff9f319a138a71dfa7186ae3cc1a9c41751b846911586dbf9cb87b5fe6fce624d693bd9edc952b82f8e8dcf5746c4b807198e9800be83587b7fb6f5fe255ade35b79f7572d8777660f92535471442e404b06eed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b06779c88a14854288614ee38fcd4872f266cb2d4aa9caa360c5fcf4f454d2de67b9388321f4252e9e3e962ac86c18dc5e8db43cd005716a4be572a617a3f5b004552ee435215f8239788ef4539c9c69ad747f22c7147fb1f3342be000aeae4da477ff0fb19af7ed2ec445db4ca153585129fb9e6051c221;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haab740479236f2d6090ba55567f7dd871821ad64ee6ca7758888e2c195360dc7055e26d8d126536541862067c53e7cee49659100f38b8de8364f00d8be28ea9fd5f657303313b7ef738c3a9248ddd61274c440b072b10c862198907d05320cd7b2b3b64fa2ae3bfadd8c5f321a6331cb07e64751a81df34b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c85d43f3ebee1224205442b47a74c5b8f46ed87d7896fc6e55acf3b4a102c8ee25a19b9e36042f9e44362137732a53c70a702b69663e3cad25841fd4d230b593996900c623f381a7c954741ec75ecbb06ba0bf52d0aab76fe1cf3c2af8bed0ebbf78bae9d00abb8eb2e73197914ae39c346c6e439c6eabbc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h179c028fdaf68325b9eab5e835c65f9f86094edc642d4d7a01968e8ba0298e38a20a13a367d3452a54fd7443feff3fdd69d1fd7e65245be40d1de3967572e1cd814f5990c354c9ff27789763590c172d03dc164af7146c35a11f0a4d1c9960385937fec44d563f8e1d139e9345f430b384024c966372410cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e53c9e9e1f63b257990f795f83f9adb084e1274d63689a083f0ec0ca668ba6c4e59de003fb65558e283977d373b50950706efa91f999ae12241c1ee6cf433326343a2cd8a05528181806bbe4b2be5a4edac06c071c1e39b50cb8c9e1fc2568f71d5034db13982751ee57d006d9c9c47b47b90206a2e2ace;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16d6d4618cb1a3e7687539c53bfadaa29b768b9b0b17f3fbd8ac701eb732aafff45eaf27df6ec67678d23a2ca82830f3fd8ce70bd7723a5a25b908c9bea49c978be7004762d23e7d924114b95f8a4f1c4f449745b3106493050f710e3acf75c3e3b1c5db206de99ae153c030647f28d17442b626590562e6d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1599dea653743edbd2a20c74d23dfbf39defcb4b52671de82f6cc986c6a400b0b8c15b5ff6bdfbc36a9f3041fd13fe3be1ca064ec2045390723b001034dccfe09276a9b30ec174a3f7945a8dfe9d565d1329a78a2c3e2ab529c2c42283e2e44efcbcc0c23ceea395c11b4d75b98477a0efef3f83483fed96c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79452664ae46694c82d0d540b7db590d0b9442599674bdc71a488632a1f283e0137b28546997078d629f4846fe005d47ceb746877dd7454408856b89b8638f0c9d67c4e8898f199adb73c73d2f6230ac40e874468b6d70cf112b1602e36d4928899df54f669efaed735b1064e973608295848c6b4225e18d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168f6c291539f5991755bdce026012ef83e9eb28c8c99c5361014198a48478f62e47e7ff359a81d5c5c38174927f9fddc68cdc5613d7c1d698d746f014470974a631f218f1f37cff6b29b7ec57d1ac18af345c82813ebec8fb6736361047449ec1537230cd6bc31b5b68b83a84756f362f546ab953c256401;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ad07dcfaa551b50e720cca6dfd5a7517081e87363820d7357b7f0f5423193353ef022cc5c5e4f2e698d36276cb2ed405588770f04de44618e31a0dd2f807f422c19a71d352eab6cca48a9551dd8658250dbe728799d5e3fc3bb90f908295300e52a47299a6d81bb4fe8eaadf8c89b8fc295c32d1115293e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17d0023b7cc84d59acf6c2090fbf83933381f80c481702557e2a684e4ca6bdc8cd5ba73a28ba2976c25b304f487c138c4291a083d93d949a966f2c7eec96ad415069f66594d471a86e13d3d5e3b5c159f631993d0bc0292b0e138f55f0e470cc89393dbf5cb5b6ee2b59c89e75f2044f2803a6ae7e9cd3395;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h403d08a97ffd6e99ed37d1ce7f96a06706cbad13b1d0c805b5b70eb6b1ba3387234e36a1cd2a771094c45de65d6e41111f151641b451725828bec7a49fb28c0766cc99dc48f4bc555443ac492b6de193e1dae6116ae73f93202856a634c37f37264a93bb2131ded1c4dea8234621fc30443c24b74a2bbeec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da02cdb375da00a6a376761756877dd1a1d7e1e56a914b2b5156e9b743dccb70a21eb32279462c5a36844260d89c83ba3ddb4892a0e421460448b0516f1fb97d7c450a98b0eaef4495e04062a970960e71c34cb8741191d6e1af1faf810cb980a36991fdec77c5981d6d0c0a1ec23787ee29fc5a3300665;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hafaea1a857621d9f5a36d5ab7d3e50f74d06c30813db4489fee751fa5c28a7d3e1886549621b3b544be6d8f27169fac68c36d0a4978bbb609408b0bc312651c728755a808885e869bbde4adece24ebf30e79b5cb12d39d77d39591375643934332f06e3bf9be12a413ae1aa146d46a2187fc1e765028a30f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc156aef5882b29bc61584f77b51bd911d658251c5c3dabec7671b28690c89dab965c7e16e9e30507670a7fed31be3b3c31d91f8feaa9f303c2063f36905948e386c8c4f298a089eef5f811eff8f83e72eab6e74f8bd9f9cca91fa0fc3d7b54c1ec788f0ce01907b8bfc137aa63a6951a8bf73ccf31a50aa9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d710488b3c26055509a7929a336703e0bfb70795ae5f8d10d0aab3dc7d0c8cbc86f230cd019350426f0154ce4fe710da87e4116fbcd7353ada697bacaf3dc5c680801480f5d0979e17a339245b6882b80624c0c015f248556f0dca441d04f374d0029af28be519cc194b4f2f47fa775eb490dff2ef8db1b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b31953664a030db92b3fee3d2faab56f80085ddbbeb1080371741dcdea85648d953926d5a77ed453c69f00ebb12fcb6e1c9fb5df917e4a8b8c2453370945f9ee9b6d0279f9af8873ce4b174da706d402b0c6deac358178fbd5631c662ce628aabd7cdcb3e2f41e1c2b9178607e9413e1056de85f81afde4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ed86fda56e8276a84e4a9d6f2377069bad3224e13e77bc3648d5fd77531adbcfadded269eca6a631981b87787f73040120d8b6c0a26f5affe2fa911cb4de4dfa9f827af470051563840c1855de12f65d397807c6dae9935d5a72f29f9bd359fb1b927e82d8615551903492d1448edab78bce5d689ab28a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1578c00388acecdf7a78d62b72795a81c46f7fb8ded89341bcbb9215aa25737638a812e922773fb85a844a3e2e4b93ec0751cd73f70c32f7ee78e990447af5bac5bf74e1dfa58491237cb6a83b4b8b2caf2469aa7c4bab1fe87ebed9312a1fc4abca81d9aea1259fd160595dc87200044b5c2b28752aed44b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h144010e8fbd888536bff4d896b688546c39aea40cff2877b64d060cb2d8ee462e2d28330f4956a770c3b059a6094277b5cc1231be59d34d69a13a42e0d1a4acb3e3dd434f314eda6881c24c6abf6bb12abab738f764ba9cec320929efd65c24f1afeae64c7f12d8088572890f8594cc8cd8fea2d928ab0fe9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35c334883ba51dbce7edd45178ce8673d2e550a890ae35082c2fe8512367aa8308af0c243c27dfa0c4a393979329dd3d76f3451b62880864b9f5f4d006932c11bdaf3da2ba3493765923df694c191b021611eea1db5622e700928acdedf2463a0e36f9788e30702cd9e12038392cea62248c2dbc11c7bca3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf710c3d35474b4f553d98dd25bc2deff9b502bc668c07a566f2e3d1f26c74edce4e9bc3fd1accdbd3e1b911caccb52695e99dbc0c8565644746061786046b15da7e91e2a700e51c8d4c29035f0d2d23e98b90c48a77e5c7e169384a52cc0a858bd619f648a136f229b35683998799d008ff9cd86d30cfd58;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9cd2f1b74ef001e8cd92536c6871541c655d79fffa47a288147949d46505df2a01e56590c6e74dd6f1346f1cc8902f4781b4d6e13e083f92087a93e51453922483a0b37bee201314632dfb5f6301c4db54c480ee87aa036dd44e6c314bbb21f20704a3ec44a2e69a3ba6aa568d95e2145546d5b7ad9176d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h127188751d257fe40de417364b99af43abb3e2a47b0c6382da11633376460a0161535bdbf452ec3bfa0a5dbced9e8c849863b6cb5d406fc6be9278800eb411e8ef5ca9c931c4d816255e09e9d321a56c85de9a61fff9fc5a22c2a72b2c57e0cd81752f1991772f03f459ab691f891a2af7e4a393155acfd1a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2dc017e93b3e140d4712cd6d44b204b7b786b8135b407ced3a04352c1e3071c6de3ded15ab582ce950bc90497c8ede69e8ca0abc5cdf6ab464b56716787df645609f1ecbb6d611db2c13b5fcec887c4ff3d23ccb5a2f5171fcd332d94841b1fb111c324b8bf8774a70a0cc644a96c01e3abda0e840c237b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b71d900812f14d9834c4ef68802bbe696e84f9fda6650c0403f6d44ae73435752df3b3382099be2f5c0f72066a68969229ebeca950a5fcd44983a61b33c8cd356cf6af79a855dab070de8a165f72a0d921545e18a890d795222ff80de2aec0cb3250b5eb8870755a11d4fea583afa15d4e454290ea8682e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c84c83fffa08fe06088f7712b6059fdd79d912b5214e613f6182d7569f23b5de24589f3bb28c78ef9f4393708c9681aacc780721100d87f3b76b9807f3747040d4261c111e84484d41feb775b3dc7aca5ad6880c745b5cf500f21d19cd50c8134456510990be8120e61993ed7b816e567184157173409df2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15ab96d1f4135c8cf432991a05c14f71e0d3adf45b99579df9b0e0265a0882cfc718e181cd8cc5b42f010897437d06009adb21514278a7a0ed63c5d0fe9671735183a7e78df70c14bbedff915927a400baacce8646e4292c426d795a957f1811e93397dfb59eb25695000a042ea2c602a63538e8c1e8a6b0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e3a14e29635cc7a71780411320b364244dc0f99992b95bad7c0b6422bd838817236a36b5bcbddfc5fd8e404bb171b429b54df61b2c08cef4a7061db5d32cdc2a7b33a72f8be032818cba062bdf4c65cffb73ffeedc6f46d147b79cf436bc761ae4c27a983b115a1112851125efc6d31c1663462b47bb8b06;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb1ffca2c7fadc1ee7161117aa01f2d34eb66329c5f1ac36e618bd75af06df079f0520c0679c5036d739040ae595221ea3b568edf35562336cc0c0336ee49467d7c6f55bc3ddd0b9419936984ca2e5ef4c33066344cd8e9586815d39e4d1fac5510f1e561e226f89ffd08ee2426e7b10135e46d5532d3a211;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2bcd6756340ec15d383cd7571b3ca50b4c105dda6874b5e8e2673543942acca0264e18f163388a74ece3015e2a1dd03fc0acb7fa8b7a39b86dee090390789015b193bce503be6b2e23071327fd5bd1d59831db7165b3628a67d70e24869c3ab7aa4752854cf824098bda80086aa4942439f39f86066eb08a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3996daeac52b3677eec39ea958373dbd0cd18ad99a606c3a36e9a1d24fa0dac16ef53a91818f8298e73aa437f1ad243f0bf388e8e9837cd0abc02fbdda40305cfab83a880c1d1f8222564bae10bb690971141a158141e5003b641f8a8153aa9dfdd090ebeacde87b73111fa8c5e023604f6576630a0893db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a304e5564b6aac4c8724a4df67cbb0464b422af4d52a4c63d2788a122caf666104115ce647e5cd9acfe3f2f2fc117756baf5dd0699d1a30f99eb7a3563274caedad2ae88300f98e83c327927242fb490be0bb4c5203f1a6aab5b5bb9d31aa5c5e88a47032b4cca562cebb3f220d3f0e35a669096cdd2e0f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a9b98263739e0aa6323b52bbd4b20ed9bf8af392e3f0296c43954467f4c91c5355b0612fc80c5cfef07d58742df28c1e6a4eae3f199e4e6927be2fb5b149897ea10dde0e67027c9d701383b90a73fce8f3f9ed20e538b6b6b264bb6cf893756b9fed062807ba14bef557bad6fafb04d8807893da0c2dfffb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10fc78054cd50075c4d48a2be912181ea7d3f87146a33a8f66c691d4db8b5c6ef4fbd14fea08ea5cb2d90bf9cd22ab5b37bdb2098299494cc01a37b279c22525e3ab5b42a1c913b4e538f86f6f373df84f4071068169f3ff763daeec300dab16225bd71b19aea48df6fcba01ad32a0203ed9125e57995fd05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fbfe947cf2fb924a4ccf295f71231f8c179e77788f9c63afb354f45f786137de82945520f36bbfeb4d8d965e4019fc3b171faeca060cd2beb95f254a5afa400c2d5fd9e93cf0e4151d772fcdaf1311b900264cdf47291d4c39f70f30ab8bd14d33cff0e00d97acb550bb9e9643174033c79090b15cd82f78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12dcb170fe7d26f650fca9bf2076aa9f0186ee1f0d2c5d8cbce47a80696313fb18d810be5fe7b84cc7fe78c166075c90dfc54e1f0660667bab4a22975666a0883dc06d62e334cbf2987eb55ea4ccc4964ff4f696ee9b378b13bc4629db9dc74e69fe005c0e1469a0afa29dc06a4f8454be417362ab6ae045b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h161f4c7c58c22d3361a7314ef45b5c480a14e3c1beaa375e8d6200f942924b08fde86eaddf711c1d0efc81865060602d433f2bdbd07a79bcccb374f3930fce49064b3e78e388bbe6eb553d2474dc0576ec4109471f6f5f4b8d97322c5d67ea2041067cf3dfbe144ca138b160c3ea2d3007155f1ad0c2deee6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h179b7bc2a88e3075e8ae30e42a2d18d169d40002d9ade816e7c539294cfc505c7052a535213b304d37cd54e4034311853bc48e70461d6d80e366644c47d17794bffcf7e7cc301b147c4b97f4409b77321775d296d5d13b481d0e2fa49519fe03081900fab505a227594d3630aabbfff30d53a8fbac74be6be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h39b6fc4b7ee31e414d29bfaef82dcc4b79d9ebb031adbecdd1fb312c058a041f8e53e836e58051b79610c08e00ce4e718db0773459e125315cebe7218aa157e2cb495af176e89b945599c20c96d49ec038ccae5912d39e6c1e32b80ddc41a4d8f7c71476675d327017c7cf0250a8ee4c5f47d1bb5d81793a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9adb7608e7461504ad8ed7744d0ce9b7f4b1274aa3dcdc5ac8216357f300a38b1ccc3f3ed288e59a63e4a46e0793db77ae1aa31212dab586fa580e7e132c690f988a99e9d1b14865eacb4f88f57b04183e360a4343ffa10b4821289c5f50c1b21f8917d0e3928b534146f7a3dac91844cf607dc7c059e3d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1445471a9e1bde687319a763cb018c68054d05525fba576e4045444e7008f038651e3b74a3e26f0573e2da43026512da63f9756e773d383087b077dbee855732606095f0172f6e35e2249fb01a1194a0f373fb73cafc3c6b56e2a7324b89384ae8d4d4115450dd8e682c255a1586cc8235b7e8d9116e32704;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2a3945733c23dcbaace634bdee2375640e6ead57c10c7ddd1e31ed9ea49628404bf0360fb18f15d09a1ae6df8379cc3fe93b4ffd318c2c4b2f9417ece2d5e2088f1cb4f70dbb27600086b9a1b6d5a6f5f37bf68dd3df7b40245866edfa52a0e42eb8b7a8f15f4c6e19f019e8841cef6454cf5281f4ced5f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12bd0dcc82a691b2067cfa20827fdb4fe29e06bd9e68454767ae4508f5f392331655b2719909a77903e6efedde21131f44c3f7d53583f49948d9558a856919be536fce8d004955e73226f211028f5ed3112a4a2a6f077996ab9fb0eb489f2d68319a43d0cab437946ee46eb23c5bc3267cb2aef1e6274fe5a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1bc256797a6d506936571922ef21165aff41377ad20ec29049975abeae6db929aed7d8c239cc93fc6a280ba915220e4ff14e152ca48c3a21c7f075156b8250b3858e177fd8c1b61fc42611509ac3a817e027ca59e610e0a59522e3f5ac2706619b8c1f7a30e7c012f29d432b91269259d7551a06b03ec05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1055a20d1df20726e33b778eb7f3e5b84b5f43993ee753dda71a9709232217bfa6d000630b4df1406db44157691d44bfac0e4ad2a34b2ed99f8cb06fa64e8b52cb9b6b51ba6ee011f501b55ba968acec025245b4410088cdc94233177a209218fe6a6a2bc73778f3e6c555a51a3fbc89773f6b12556c0685;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e1168f899786d450ad1ff6b4951e0a33b1d9cbc272180f3f754f74dceaefd0729f225f7a3a89de6562b3966868cbfeaac20532cbd6ed05c8ccc9a69099275ccca8a1bd7244307ab8e4764911431cb22f8f8455c314fb778d08d305b8231baa2a79732c9f0f0e9d8fab028b6826195a1b56fde310d42c37eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19cfa634e17e18cefaa35a8f318722246edfdeef8a2b33fffaafcefb046dcb595a974024a2bff1cfd1f0c0c3d90e4d3fb60131ca8302189daeeeabd5e64ffc6d3909bf55921cbf1cf011d7b71cd607019cb98b522a687d8dd8f136ce098908176b23cf88bfcb78c5d20aa8e4511ccca15d7e5cde04576b3b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h588b8bf71a3b1aec98201c800387f47552875c00bdf3774ca7fbcf29bc03051afdae730075449a09a33830bccededc6e6f367dbd3634b86c5f63fe085605808b3d0090b63742b2bb2e3bb361d01013b48663a9d3f96cc074cbe2b788c6be417adf54de90792c8660ac71fa053f9540f9d319e8d1a4d8e714;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1393a975a8aa6b5d5173c8d77940f6977b0dffabe71d6cf67bc36cca74f6b9052e9e0c15380acef96df23c3feacd30050407025f95941feadb600473cba25701b725300f30334d913087b7cb6ab4192b96e2cde1d3fd5c8a9c7387edc8233cd3f8d4b1ae0c9c57b322094a78a3a965ef81673c721f1aeada6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd70b4a53e82f587c31d05d81d734aa4abc5088b24835cb4ec49ac5490002b41dcf2a608f4d542125cbe6a64ed2af99a134d30baa784a565d70af8107f9ad125437d3c19ed4c39cdd83d0f1ea3106ee790968e3b2d82a2082a7fb7af969a6a67e7a0344eb1096cc0c170fcf05935cdc35f01b80f6d9daa20c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7deccd2aaeb33148ea11d2731501bd3881c6158db85b14d8a07a366d299524af0bef0b36652dcd9167417c2f3ba89e7e4872795cc96e5ca9c489269c38f0fb31f9b45267b39c0c2d299148e50add2f61fa28ec4477cfaf6da487316124a30a01ec4d686cbe5dbfec683c6279b43fd8d875625a82932cd51d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11c7bc39625c2038164f23d6ada963ff2823e00f8e941abe8cbbdc1284dd59c85314ce50a229432b4cf870a8a5b31bea4a36203ea7035943afd036d6756fe02bfb884a4bad661f8c7623b51a92f4dd1022c192ec8f9638bb21204860c5bc89220ac56b9182ea98bbab8a43a4e9962a44de0abb7cc2e8b249;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc089521b16bad7d384aba87d310f2ac195bac54c30c88c50f9be486e62d531aa3e1ba314f4355eb3a6cda2df34746596db02c9bf13778d6ca9d5ae17dbdedb8da330e330c4ffad2cd196ff37b905ef77608cd9c52cec3ad6d1cb1a1db1ecf6f277892abd6f78040103074a013d8b8547bbf6c58f09861ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15ca9d75efac397f2580295d8c70427f7054954ec972f41a40d07c5448e04c63872238646e288e3d2e081be7febfb354009004c57d547f38ef7a240b20579a137aa1cb46c6692f5b67ccef1686224912466b20c47f59596851831828a20044de30d29278d903bfc862c21b5727835c7485e4f057b7970bae6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf3df8d418bd5fb7d8931695c3b485b81e07e2607e07ddaf6085c1cd77c1bdd07e215820e73617a5d1ee14fc790e4bf632b8d8fdb6b50aabf73a6d5b79c9b1a07c2c9baf552c53474bbef723219a2019a16f4c2a19fa8e7cf397b03c5cac5e700c740b519b6dc8fee8e5295d74ca07744ba0d87c074fe990e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a133fdafc53cd09a717424bdb3729e0825a9eaf8fd7cc91a40bb2bbc7b2e044a506e981fae0da7e06da0d3e65e21540308bdd418c8c3aabf7b16a030e76becbe85e3036eb849440216732e9b7658e7475d0e37335c888dd979b6b6947d0369d4b865a30ff4be6a7f4146f212d15195fa6b5d6783bcc48f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2abe70045a36c9f017661ce548354f5343130b43a20d0db635927dc9cb49b721aa9a9aa0fdfbbb419f2864cff6c5f328a42dc7a0439b5f1a6c9743d1fbeb25200ba4e482a962e1780e46fd22c30de28d94ad1a187bf0c448162a59baaa02ce2e7fdd3417bc353c1040569b883692b768409e2d89c242be83;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d3c389579655476cb9d1fd5452aea9971c8df3d989d3dafda3e2a08b84b8e1e419ba8476b71a0b2e15dfdfbb84f56c8142dc38f2bf051244282ef427ed1954da2982c84aa805326e7d791ba0b018a48e258bd5acc671e16c3dbae81f40a728d21779a62351aae8c6dd0840cdf2fa027c062b64468f2fca7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc20356a8f4848a16543e4f07aaed280518850709b4e3afaec2a68ed4950034c7fa82d72ac7e09fb4d6c6e54da541b204c7dc828ce4e1078a6a3f3430f7bc3b647036c3b982f8a71728800a1be64242d1e30e0e4476ee2845d3df880c824f37b9fc36d52e182395c49f0810e561a3cf4f75075c944544b32;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15ae76029bdca2af8278d149d80858c0dcdc748879ab5bd1dc316311f2a78671567456841508d17748b950ffeb1c183fa7d2126a3979ba86fc6143e915a01c5e04518af32d469a79b0b0de359ad2a8f7bfb8b539c098e12ac3eeb97a6d34127f2b5315da74ccf684512ca0b4f20e1104b8eb36d865c5c349b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a8c2dc5b9ed08c296ccc2f9fcc5f6f3f499f3c41fa4cf4d581d0cb7258fe9af439c15c9898ea74bfee0b8257bdd09ce38e217274ca4f3f1091f1c8e61cfa76b834a199045cacbc75232c08a3c07972b7c25a33109085ee00cd1be092033e882028c0eb838b6a101db0934f39f9db134a81fba4272fcb086;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10dc2788739528fb65aa24b86a0f94099d98bfb376cc807de2f879746dea68347ecca43ab8b545a3f24f3f0b2d16279ac2e46c553ac2d5cc15514b727bcc9fd7ca46fcdd12d434906f803665ed7593cff60bced1ddb1414e2206f1f1a8eee641e71e34439dc8458c90f6d17ea2bfb0b1a2b8ac96d07556d19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he2b950c0f4680c2175f1381f1a8f2df259d8d14a6693f430083f898c7c7cd014e5d65c7b167fdc78dbddfd4964bfe2fb9310a184539f3925517a0493a7e6ed25d837cef645cf8b63c11e9ddb40efb705215a3f73437100d557c30791b631916cf44cf4b34c47678ec0e26c8cfd1aa1ba3b75307905e37d67;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbd8936ad4e3587e809c8d20c582e255f45bf2d144881e78ff23c59dfe5740a192c3f16a49993d9bfd684b27aaa098d99f76aeb7724ce1159f7c6ea6d2de40e36a2514fbb50e5c3e0e9be3af61ad8dc028325cc50c83580d9cc5f41277efcebcd0a92bacc4876027fb0dae97950b0bc95440722ecae7725ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19735e29f6101d0d0993809f7dd64491f182ed8768d7921cca48e1ef4cb3a0a37b7d7a943e4e0ed4866d9042182945739ab14d485f49fb3b8e4a01c1ed8b98886b2ed774299ad1bc85348b976a2311b06953cd36d4e85f721d4a2c62d2e149fbfc2211c349dac452ff7adca09e051bd0d16e4b9a95f532a5d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117f7f9d647b28c686935bce77063bc3253c9e8a840d43e66a7436e79fe8358ee6ee9e3868fcdbdb1cb69dbe5f74e7ef171fe03c93a5176a5642461aceefee1d3726b30107977ecd2bf20818a0cd1975b9d01e4f50703542eee4e74ad23d6f527753db1d39ef48d2aa1a56041bfc5e98155b6f5399bd9ee82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b14a6406b3d48fd65e1edd5ae23b34c89595013818cc00b5a592bc563a8b3a0851177bd60c8b19f8decdb1bba5c81e5fe73cc1dc74a065318d4c012489a2592595f9253323bfe595490a231253cb88b6c530a9f71bc71d2efd7d2061d560d29c711fb9e32f25b27c13e47addfc6bf810953dcf45d7390769;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h325684869e88c02a6f0878e9e2ccf4771dacbf14fa0c2b2dfc6f1572545504c8dcd30367d4de471df6b5d227769e2dfa62fa679a142f608877162d4c5d018f955bdda5968d1b41c92b44f383ea79f1f521a1a7b22f169404b8271d248930de838307acd098dd655aa6370cff6824c0dccd9c8701a4b815be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c126d608c179e66d8c6006653cd57542b1c397709c0809a65b95d66cc13b64b96e42cc38f94daad7d3119c0618088d322e290b7eca62791eac37bcad124c841a615b57c38c87b84422d33978ca3c6062e216fde742a84b6fae44f4dd2a5d9de8695bc4dcaafb2093c924abb1de62c3a86ba7c876609e7036;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4f277bad467cb430298adc08522ed1265a857358209a57b38f286bc77e262a167246a038742f03b59428b562b6993ccfd582281da9e3aee8c154d7f3c20b777af6bc25bcf9234e2a6d72e3ba94c4fb0716413d2435a992a07445981f393be1876f30f8fadb1e3cbdd587e66933fe049c72e14d2f89bc7eb1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a7f710bafe910b2a0dfd261b2649f59d098746da2eef62aaf46c8fee001fa23822056ca7d545c55d983e9065522e3dfa7853235c4852920f99d1232eba8be72c9fc3e988fb4d66eb1a643a4741df9a482a66534d722ac9911c77377c8afd34c991374c41f606fa54ac93e5a3dc7c1834a5cea9113fc9e86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f83924334d0783a175078ea74dfc83c94b15f09e54053fe25e047ddc6de371c5038023dcdd17464e88064ce841ca67448d9c00f341c7cbdeec79d9839c9f3c88eba0820cacba478ff31637ab2b644d7502fab7bcb0b3475def4d35976953ec00a2d014ca875aa22c5bc7428a52d1a172e7ba05e99dd0500;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h283107280f986a39c4ecff95ab93ed511aad135e8fe913a1fb2b13f7c1c506a74e928a36b30979097ef04e8d78e0d92a09e83b3ec086e12a62cd9286c35eedb772fbb26ea036c9eb02397172a7370be35358ff6d47126384f0f6b425e97cad943210cbd8e964bf3e020e27ed7e8e0e88f593dae1baab093d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c7847fb8f8f9b36d8c5c17b0b6ec243125909cd0c683c9c2b17e36a1def0add436ba87ac1d78e436d32f99aeb195ae248866a3712ebcfb692a359c457b2905513ca58de9ee128b338b36ee9ae955c4dc7e4ca507a9b33c62c0372176ff081fd1497de3c77d5b103afe6e462f513dfec27ca0fcff318c50dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b929e66440b1cee2b490b992fced9070409e91813bb663eb0e35b083e15c553df198538dda31b7760ae3481b1812e96267b83a90e6c34528f5e45f3e7c56dcdf9116ea2f03ecee3774dd722b685825d646da5817aace1b19dd6f15fa9aafda2817bffc04ee658fe89b3e0ba3384b165a85252c5e5c44bd48;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9fced69c4a4df39f53cb126eee41b7051dc3da7ba6fc73a1c52bb9087b50d94be03e2488ccb353f1fcbf5148195763dbcbcb6440c203f3533cbf9490d7e3a832786267f0594caeac9c83d5c0ffb9209c418d401078eba86ddc7ff693fc4fad8c5427777524cc0e2b4f6d49cd6c06f15e46296c265e0be17e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c5598e50315270f0501f55f47c563ee78904566419645dad3b5690686afdd163afe1ffa4d7164f1fcb1a6bd71088cefa938a976867cf0f62fa6cf4543165bfa8e5b1377d0b194348dcd334b0eeaca9ac0753dac4cacc84beefa06a66a99e06221476c4a3ff8e1cb3d24fa484ad17dd55d11f965f30594225;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bbcead35242dd934ceae170acb1e8c2aa5916ad96517ed057a7e3f2e7a1165389cc660e1507250fc6f5bb684f3a675fc7271fab35b48c77d415ee297437bf529aa997f1e84dbb82ae875dec3dfe3a6cd75bb2926d116823f92576d6866e5812f688f7b5a4df95c830aeaec65a221cb9bd9f508c55a2ea922;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d5c6913cb981116a77a7f5cb57da88c312d265bf9bbdb608eb7d27aac919716615efee656de39623d58349b1c58014b730da65ecd0370aedb0aaa43af68f38601fc675b7626096e9874e488af7356c19639fa3db9aa81dca05848f2409cfef9814a480137df0fbf0796d8a676716a2091d0db132f6738476;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd04296df9294e24363c8b43acef5909146bd882f591293b040d86af409fbfc704e9cbc18defc7635a0aa3bd39c214e75ddc51840a54ab529b7c326797a33266db9a6e7db71e2824aac49cfb042ac0d37ae13c6126c4608a44f57d24bc0779a313d0df5e30e992354021d0aa201ff73402e6afd2f06ac247d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h97cb922ec6cc51aad660ea1d6c3e02b870a9af86a79a74cf43bfeba44d82ef2ebc3dae7e25d90b9fe96ad37bf8a48fdc07c85e241aaf9fdf729c9a5d24790c9b6243ec113584b3204964629c5ee3c7a5198e21bd633639b4a7c5b25c451ebfb8c62ac468fce1612f213b5b2c897f296cce98aabe4374a555;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb0f4fe6c3d52d84abb5678c022735282079ad4077a2326abada78179885870afd4e19d2b5611c0ceddfd203f5dc2dad7aaca23e7e0ad02bb762c50137c79f4b053ca8c514e1284d0ed0b7089d4560a0b92539c6066c5cd59535811fa2c0a77a7acc9222e8a30dbe940e44bf60203567d717c53f65352141;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9e9fa9a50edc0ae6546c12cf29a0d0da93e6f34c1dad65593269a333c0972ff39c8367d6855e3131ffea2bd4c0ad3e1a3eef44be7ff43e3427fc514ff2999d125cdd79a2cdad2146b0d8d90a63fa8806d545817ef9a3cf1209814d61f7dbd70d79e2115a8efd16af0fde24b8b18b951047a42551a0dd3f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9df146a3208357202dcced1190e01f96d4663489b18d4c72de06067ccde22f890469da127e07d388d94f70236bcf06420cca3a7c712765c71a036f0583094068c52757a44ab792b4e160a089696f05e9bd893ff4e170c01808a1e115ec66a806af60b85d3b8f126bb5ea19a85937ca22c3eeda6b228a99fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa25a7354b72eff3cb91d44be0898a4baedbfee32ce4c148c7c5ca824dc99bb7ffa4317b23e4d03966e6753b859dc986516a92d07dd1c11fd1b8352bf6669eb0b407dad0b7d908385d0a6f6cfad750117270e49d4681ed0e2f58f1a027dcfbac42bd19cbcaa5be23d0b263dd157703e86592b05512884930;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf4473a96b9ef8aeb280a1cd91dd0e680438bce3d1ef36099427707e5dc595f6a1bdb8fa9d49ad5e55ad9e4ef3f94f9da05890005f1dbc24d700eccaf7df598a7bbe8057ab8eaa8f44076b7c51650d616dd340258d71084c44e2af97af6770cf712c24b3eca4acaefe33617a7a739cb4c00ed69621113d53;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d17b71786b7a3798a0bceaa59c9983b0489119dbfe9af490584cfb3cf30d4a5b8c781560643278aa8e7dc2dad58b2106730790e5cec5ddd885b10e6ba5cd5238cb4335720ee1e9ee6d9e7c238d03de9e1f42e8511b6ef79d80becbabe18db2420cd962aaf4de578d3b9a60ed2f0fdd06953fd699fc48097e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e1b3baf89356b898987b3153fc18dce5965b06dc5ae7db2cac5ede3f7f2a7e4b4408d9a3f6fc6230b1d94da1f25b50aafd595ae66787fd04e2484fa25d25b1460fe816fd4d1f851f1272de21d0eb5097c71efbb023fca11e4d48d20fac879765138e12867c27c6dc9e1ab9a7bdb7014e81bdae1c613808c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8bcc3ecdf71d5d98d66311323de5573f0a37e55a898117ab3000484f888b20b3c4b75a45e7bb72cd34f034eb40d23fee9b3aac503c6827088f2b6bbae2fc65afe1b6b538b1d28b46874d1ed7726ac8a52f0f00c84625442cf26c22687a65a1d2a187be3986c2c6dfa8e092caadcaa7d560e03458039ec87;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d93e2e1544048efc816b726cf3191ef4c42738dd821813130d27878169c518348b5b1961a33ceb20cdb99c61385e6c67ed15ff98219840e545eea00dcad362dc6777e2f1052e0947ee699ab2d58df9ca65c1bc85a46a7714501c88f6c6caa026184624bb4e505d901eece8aa1686499296ab953e2fedb700;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h157bed5d871952e2294345180a39a571a6a556e4bb6551c46d40145a6dcc4ca26ff9543d4d3ba5635fad6456dfa7ff4512ac72f500c937f62d882f5468f1f3d6af9721df9d3d678d65eb0c2761d2a97c0abe2cf59865bf8e580f24f83aa7546304a9cdc5ae6aeb024787473468153a91413c1ee7e6d83137c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5215388d6117d8b9d3d2bbf7e81606482a4683267fbb76b7d2f661ffa0eeebdfec65285ab888641e77da70355cb77b489f64b7fd5492a13938915bd8f2433f940873f7f385799c366aa40509f05ea9d17c1abf04c1f7a00b04dd55c1a5a147b0b0ab5ce3fdae97c7f226459d0ecd358802d5612b2f53fe3e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ff4eef06fc3476b2b98ed0e72846879145ffc8c65b732f5ae3967b8df4594181ce6f0242ae035b873f8029389453727d61921b4ba6a612befe8742c1411782cb387319f842f6bc6bc6b46fb4dc7195167b2df39c45973e550ba11d6835dab7931b6ff6fb08679779132e54d20b56a70cda2f080b22a1184;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18f14dcdfe89ad362c110af48bfd5048bc142b7d1b0fb94d8b926686603a6df8d04bcd8b6aa6371209da13a938b1203869c6b996f4b3e746fe9d93ccdea3d1eab11959f7ab3e3c4a37b2c1d5da297a6264a7c7f17e4183375d73f8b6bf92fde3beb82ba26595e054fa62c506456e31d43e384631add206a4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18439a528699585da9724fafea2d41099d3efa456d112014a86697b920fc6d08dbc080434dd4f739b87a09e3f22b021c33fbb95af83af480654361f053f844dfb1d9b718bb89e945142df9620166ebe036f09fbbab6267e46d57e781f94aecbc6c8255206c9f1355cad115034b1dfbc3085f7a6315a42aa99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h182af2388ac38a54d6038ae1a41135041eb5fb676dc86621e25b976d98e0db36666a0b6020ed68d1bf5c56b51bb1d57fa4f6016c84bccfe3f31c5f81bda18ae791ce7fc0b29c058e994c0135e68bf68c347682788d8902bd8fde0a37b8835786952e2bcb3adbbdbb1f272e569c9c144c45212f7de9c504542;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa3967706577ead27faf03fe2b81eacd9576a5839fe707343d14738390775afd92e702609b3bd0cd3007aebffdad0bb6055e6c75de3ef6ff0c3690a3736754ab6b7928d14248afa0a9d69c3c39889b3376de378416fb2b2c79a33a189a346054490d663b6ddaf7707c22bed892c28ace42429636744d24c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3dcf8f6e189d705b561dab4bd9d4bcc76f41c91ad6b0081000fa25a7f37a8f8a8c3fbcc4c169c6bd01d15b18426370910de89aacb715730391ed6b1f1f4a2d4197839c3a55551e4b6ede1da8e8a0c6b978439c0d2f787587712f09b6e47ec2230d36d74db41626998186158075ded43faaeb48805ba0c7b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13652d121dc562df064b33e975f3c1980d4179d463e3de1cb446ab424425ad7858a34fe0f8776a064d3618338c3fd3c21d3da2b93dcd7b055672eb5890f3ce09c643eb9a8cd6d7481f44115224d9b197275b2a62b99d21a05dbf38f75f072f7133e7edd1b84326cdc0a967137da7d6533837e98c51f00892c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f26869c000024190d9e6474787dbcec9d03674dd66aa476bbf4d40a9c891cb6a2933d01d3d19537b1d6d630d9ad93e71c4d527f17ff00438822a2ac08af67a90b5ff2c847e4b63ed3264fef7096b4eed185cf3c62822ce8ba2c75482c9949e0cd068f1bc4cee48e03599b6b005b36bff504558f5153ae4d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb1292f7efb9874b316f9d3b28b80ed3f45230b1e2d480e61b741147a49e2cac39138ce5f200f94b4b633986544eed727ca43b078a5c0e34eedaa2b0e49738e0fdcc12396a072b0dbeee11c86f9a3ed339996404cbf14960dfaae6ed5cfd24bb9425990fd401eeace8408de030bcd9e257be95cc6efa67460;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4bccb701ae8305425b300b54543ccce72b9d43d378513e9aaf71e10037b30197d01b98e8a431706c5d75a9ae5721b61554507125c321b896a2c154985dafde937aa3eede0b0e61da09d415e45ae54d01b2a4d868a23a8979ee3870c11533d808d8efe1c54bb0a8828d1e73a49872b26a170c2e38804d4f74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hffc7ecdf872994bceabf81c72d6b09ac3ea3065dfe413d8eedddbe793ce9e309c032c278d626394021398cdbadd199ee58bbc1388215a19a2066697573157d1776d10157eafa95144e7cec0ce1d16a8d91334aee9581bd66a367fe211fa43e38d2f19e57b7012ac1951584425ba98c82e9cda362e9c337a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h161e85084125f78b7685dcaa7e3fb6b1ba786bff213327255841c0a0af1e4fc7f4d9bbc20ef1caffd29fda5ce6077a41bb166850d9f65cb0e2a2fd24b13cfb0bcf1c876756775f0dd7e61baad02ec409243d28515c7192e21862f2da9aa30023cd1cfc32b64bd61c87b70baa781a7df92e047290b3d84a280;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb2391f91d23b4097ba8cab81cdc562e463038297066c363c893558e1fdb97c6bd07eb9b77c56064c35bf655b072ca062261194f391bc19f5039176bca816fc74d6ec4d780c0b146e2869cbd42b228cb63a7e98e95228211e93e766c4fd4a0500ca1ae7f0740cb611473f0e2f508686dd3920a2848900bdd8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hadb1f9f95a47a0db0b3d57e73e8ad38df073ad8a40f7a488484410820bbeb81be487425cb563f5f333ea2c59a517742213c433c20b73f67a2d06fc204087bfa0664b03fd3735e5b9975eb2cbdb1fd963fc13bcc6d41f2b2cd89571e9dcff9038d35db4714ffe3de82e0c18cdc458b1586f9210566c2fd87c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hea20552f5a01adf96d35485237be32dcb3f3840b63563451767731cc8e36939563704e66fb609d75d9638ed51c82657271c790efba2ea3e8702580360a2c326f66a2646d16b80a07a78b435233cd3477df9f9b2f6eaeeae433983eb0de3dfbeca69ca71e5d608b09436316a26a73311f10d1237faad0d57e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f8357353faf096c807b11c2663b504ba984dfbf0c27658f5057e3555b395f486b0ba6c45dfeb6c0bdf4c9e6a0e489afd4893fea6e8790e18574e2c8465d48e4bfaed5651b9cce6d73cd003104d46fe2c0f0017f707932a3fd82b3b111599a1ce18452a45bad55e1796b7957e514d2c98df3de2cfde7a49bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c06031212b89bbc02a3eb5a8b53bc4d33bf415446047444518ff2d725f05070ea3c1e1ced44391ff23c36cb0639f774f0c1754f096ba244748068498dc2ab651e52ca5d09106b5c4375ab3d3f3d4c783e33522b6724cd8582221a4e3e690a1003f0729a26b00e1c25a4d13392641121334e8640ff8660f38;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8543f6f1632bf09764af1a8ca75b773c07a7a2fb7cc9f69da0c92b0e7beb950cb15eafcc5f5956bdb6ae3021e459b55cd586cf005e0fc2867a94f18d3b115a5a6364742e954016d7dcec365ac6667158f0bb0a8113d67345996da6092e10702ef8c787821901f45ae8801620741f79bae5de77de3b7a196;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h122a0b8aae72212f8676c248d23a4abb11124b2fd5362db297d262c0b604a53b616ab97aa7facd6936219ce94b0d02f664e29dd97086232680468263c29130405135f42accd5842b81603341cdd4e02fc2ccfa4484fbe3d2c70eeb74a6fe22ea9ceb7eab087b432bad92bb109937bb09b7654e2648435fe8c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc6db13b99a4d640943f498fbcc9b7ed87a19ba625de1d4fa4022bde2c6a4eefbc6c97b1cab2b62ea350012b45a174ddbbe856c45317438068a3985884a0686155bf78d8bc6985415561d6f7d6fc4fa09c29bb355fee87397d6562f9850bf47c1bfb8295f57aa451238e687e476fef2654baeb1f5228c316;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5161031c4327e55221ae84312d2cc24acaa5b5446ed1d1d3ded8cdfe66d7bd64a632023601abb42e4487f221004bb58daf96c469190ccdcf993b003bdce78ecabfb5557655a49539c5ac3fcb5fc2d03a6fac185e449e46705917daa65d4b659e7e78c49d29f0c83871f38bf939e44441a25b171e5659804;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc32a59e9062c91bc5faa198afbf095e24c2c4a69e5157c36ae188624adc5d743227a294536c6efb616ebe6d6d900e9c439efd35ea4eb9c31c8bc9ba838f822167bcb5447443a7894dd61e3786c805527616a466d2b5ac65aae8eac087352c7f9e85ad3f6c3b356d445ce6b05401842168d1e3077e262cac4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bdf15d90f5485500bc750aa6a9fb89ce647a4592deb9d0da8f4fe28f95fadb4c8a7269b66b45a9e8fc4e220888faa5322a5d9184dbaef42537fd591f143d27ffc4ea89f0e77f77f9670ec9e3908163b5d5379a38f2171e8956582d08d2d80d711bcc2a0a8d828e60ae0e607ed4601715075d63cfe681cc2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h73253ab3b87eec963b2768be2ed44c466423aad02716c7b0a8aa303ee9bfc6d11b26f263962ee1eb937029c97bbef45cce9b06785f4ecc0fcf597af0603665cdc9e77f58d5fa657b8a40e4519a40ad2a2debd9496ae8ac70ef246e7e36df7231019e63065088475ba5032485d0ca0c6ba16a021af4cd033c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h134931bb8c3255ee1976beae86a2be31f624efe29b12768603ddb28107688cd900c7c172b05f1aed171fd38ddf240963ed21b3bdcfa1262f660e36eecef492c12c5d7a646fcb9d3527046217faec934d9b0adb1cc51e6bf962f10daf5f6d700900e8ca73eedbd719d5d58968c7b0388f778f429b978247ed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1874c876b809545bc34f21cf77b961433b077c9393eb051e7b2d70d076566fb379f9988d138ebbb2eee99eb877731dd6d8c716f5a431bbd6e8ff0b42284e735d63e7c38c1b44d0731feef60a3e957c7113434be3ad96a923a92d553cd7fc77556343530fe127125cb7d1d68540895542731b1a0e0729a3643;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c744a20c608d3393c9bfa1e1744bb86871c433538506f34ef554864fdf2a7571ca246d551bc2a8378c4c9470439190050ae3495f712a9f84b4c890612cb839602759b86efd5a3a3b7ca6abe6bea3fb59b90b92de09f7b50f231489cfb517dc36a149693d0d88c523d337144cc786828f893ae46a4824d9b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c45a8aaad7351d943cffc41b5f8d8b917b8bdf40afec66053fa46f31dc9fae0076e1fc4358c81b3e841ee4d25f23e4dbc7c7b1d7f8af37962e10ba735fc83c39b5499b16ff90f26d2200f3e977ee5553b41ab6afafac6416baa186dad14c11485ca6ff71efa50e8c6569dd364ae356a1e7eb5fd1107096d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12053e4463ca60badfad68a6a1ebe684332a50eb28a2aff0dd150560adee30847ba488038d89c3ca764ebab8036a92264ed00886587dcd639d610bc4868213434347f33f256a0b1f5702f4bddf0e487f9ba49ad54696714a4e5ffda1c584f76a8ca12e52e0bcb6b78a9c000099c76842c61442fc26dc4f0cd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h148e1d9d7d4985c3c485d1bad8be82c87f0332db9350dbd937727f7a7b68e8a0d2d25c1b9eaec2645a8e3b39106fc89c17c8e9f8edc1c0da093db62c33910c3a126251c84d0d9546687f503f85c6e9ee8c2a669dcb9ed4ac9e6aedeead1b332d8a33e1ce1e23033d040e4188a2bf3b217168fc194d59040d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1529dce6b2ca9e9a70245538f8fc472ae1e26e45b96630c35162b4d9212d68946002fd2c0c6682bc036cd22fa48fc7789fda3ef04975ce7c839bc7319ccee7460a676c5bcac04c52c189d7a8acee35cebfb1a205d5703cca5553e0fdcd11d8a8d285385ff30e8c73f09ee80caec7d4728066fbe8609410f6c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7f53d8ada6e290ce21f723f39d448d3cd3d05db89c8d316394f7eee5ff8eda4ab849679c2b217d1cf4151889801da33a364f67975103ff4da0e7f462c0c7bf0c1a307e47c395bc41412a1227030d6f6d8e57003920d5b85e7d270b7a5017ba4aac25ec721db992775bba7b568aa10037da878f3e4ab25855;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1c5ec12b36e6794e6e5fd78eee3f306c6f3a9451b308b33397301ac98ba5e94b0a3a9606d81866fd55bcb0f8625cfd8f1f678f9794cc18c91a2c415fd6b0c06746d6775094b585cd5672ccaff5a588fdb28dc4af75f7c5aaa2a1c1096e20199daa786210099c064ce743dbcff42aed4a1adec11a456d87a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h24955ea7dcba838980d91d996c135edf12343daaf41ef1a6b4eec3fb2ca5fa1ac0ec7570df29b57f2a98227567ef27d5f6df1709d8eec7712f473c1061fb78b8e3b7d076b7c812d678f099e240f559f5237d2f762437de42c4cfb86bd4cf6e327dbae0812dea5248abff90b431c19fd9a99885bf00c59cf4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha244ada871ee0168f28fb6b53a1111d8c4a49f80b322ec0f74d98b27a83c72a1d103e43d64c44c4491adf75751f4200b438744926dfbbe2d022f8622d34f59bf5e0f69267a64a7777243c8689dae4d4c952a721b4331479a7f4ff67c59e01d29cf84c0b9730c0856ecafe07571be148db6a24411511149ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f3dce8ee7cc322a3ae5e39303c25e9822a89dda1fcdcc3c8ef7aa90cc17f8c5e10a946aefd84152e276baa449b76cfb300ef136d306e486b81a1bab000bd7f89b812377d37766579c2dea46142f15ec7ea6678ea2547274471f0cdd8f075ed8034e2dfd62e8dd9dbabcc20dbe5fa68c2f08098c30176a83;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e7f5ad3d0344ee388ec0f395c6c397096adcf828d32204a184ef7ed24ebc6985005ea0dde687c53aaf58eca5f1b8c0694b1f24b7a640be8d23ec65eda9eceaa3af911bf1a1c9ea0f43a0227f64df03fd1de6ca379e6519ed67fde05672bf10199f84d3d8064ae859421a033fd6c021a1d978629d17a8c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14cd109f108355e7b4002bbdc0bc6db8d9d20eb57984aa2b4cf6a33ff5db33f485720991aa4d4c8d2f39e0b17209aa78886aafdf5755c7d792a1cd40d9dd69c360923d8a23e49d69c0651602f7225325d327b85432bfb40de2740c3270468d896137b738b88e71f53e4a337c5fd9125f6df02c92d5dfdce87;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e506447160958ff344e8e47d16efef77b14b25b8236aecbd944e57fc6f1bae45ae1705ee1d2da694872b06968006e2bf682eff90a6f2e56b53bf6453ee6178c5622c6443432f09ba90cfa996e52af9d40c2e9aad0786d0d48efb9e39048b75c0d99476896d600a7931a2c9a801940d19ad7c1c78745c3bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae543a8cc93b5593380c1a0ab603d3cf18077db9396509d12999252f3824d8dae80868b769a6c7674d06264c9cc9f96df5df97afc8f29abcdbd496b2df98e0aef43b099ef4865816a9199796b228c0de8f4e58ed1b37f3fbff5404ee8055bba929fdebc35f05681a761300dca5242fe31f252e0a4278458d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f14f7cd95a316636b16986de6e94eb8f135ef9830999db0491efdf16d99298918b46a5ec061d4ee3bdbb6760a060de98e96c3cfa988a9a94f2208c84af1587fbdc4734eb34184b2a31da8457804687e75e69e970d839b9dff31c80a2b449c2e0ec861aff3f2434e3e792df12a96c4e21cc7b76a2cb7ab66e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149067d55647937449c7eeb47d59e99f9e751dadb6a155cb28405e147a4a2f5e907afb57c0a734f88fed3c222000385555134ead3f44f5356eda4d914f953e31f525c846e3a0ca77fe13515974eea6a279ce6ca2e0718e774ecda775c47aa3ff7124ec994a630eb96a8b5973496c6e70eb1be1e9e1c24541;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h125848f67e00e1fee0702d821cabe7717fb94f0f4f8d34cf2b3b2b88a8fae469282b1524780af4ca73f661ebc08b41e72e1e21fce7de606ce0ea393bde396abc2047a2113674222ceeb2997b1960a6f71c8b07bc45c3847ff1b4a2121c371c1dc55fb588db73bad974f327b1f8c912590dc60a43688e6a9de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8662b66979766d41041a413b2fa5e6e0f53dd865abdac6afc46abc040c372d72cded28ff3225a4c9af9f9efa7f1dc0378cf5694d19d70b9aa44d085e11b5f5f7f9abab55381ea1948f7346a26a4fe6db1c73642638c18e9de122052ccedc884f12199af725497329c85763719317d9e2cd0cafb5cdeee346;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h28d0351d4de8e4788f0ea9e06978aeb4080bcff3949c6e9e17d62ba1b53d6f6cfa16e1fd7ce3a081215204beb17f415b169a0c6cf8da5f808af7ebf7ad46f741685ddc4db678dab82485b6b54ba21cbf1dd73dde4f42d7cd0438d625c6044ec574edef5ebc899ad10c863b004a72d2915eff8a27652e391;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b22b6b63e3af4436782c690970d24fca2555bc8e66a6b5a081207448ccf3d18eb4f277efc0d6d47358684e994dae57aebb287d196f6a97730e70d27c9d89ca34f186c64467eaf72115b6befa09063be69d45864b3da233dd279061338f335aa3122ec635d17fe232090c329f6a8c91a3707a7f13962e875e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11906eada3ab0e7cf35cca34401e40bb6fa60c70a0ac3fde817c8a5f3ba2e3c27094f8a2c6ea2e9f90127b2c220ad66230e893ced75b9c0612df20b237114b8c358407d85267583e51b87734874d8576d2e1f10700e3eb5aba8ece8b9922cc96c8c0dadbd88d4658cb16dd04442b6b31243feb7d34aba9c4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f38dfb0602288592cbf78faa194d468b8a041d82d67b9284797fe5a9157ed5752b201283a69c9f2141e7fd361ae49fb09ba9c095bbdbd3992a8fa255f23285b500cb1d3ba943cd6ae5405ea29d2f9eb6f323f05c3b87d9bba8e71b0d4904501723d085266e12312b6bc25ac89c803a4b1bf12de6a2544bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h32004a5afa7d7f05063e09c6075f6999f6fc071d1fea28042f16764a93c8b998910f940415db052fe53f94b63e2266ba562693a4bcdb3607aa6ed3f958a9e471be73167c024017b32bf6ee43958865abfb478c63ed3b3f01a1f8b49ded8a5acbb09c02b87307c04ebe6ac3f96964c8782d3a33288c4920d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h135556064d0bdbf98f9b89abc533c37c6c9428a18cc44ee4e20a9f75b3a5733eaa36d740500c8ddb929612e98208cb926c4edb5ac520964f3848ab925fe1de513bdd6a0e67852a4625ce369a3ab151e91a70e693d8d5998083ee766b5f8f0239e64fde5ab2953cbb163864ebb69cc113260480895abbc5123;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1005830de2b43a9a79aab271dcd8e5a4e5b7aad2539ec31c8b1b9fdf497d1aad913086e0cf126a7a8394145254534b3690956888d9309baaf2e5831e22a20155ca021da6a979e2a16a7b58f3f98de64af4c85dece3b2dc05150bf21b2e5e119ce1332e46fdf491e2fef3331cba16628a4cf0bf2b86817d4e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf148aef7ea72903dac0866a932dd8b2710ee105b42ce87ff079924cc3f37ca3e9f50db54c2d302d340b0298f5689315298c1c20a185705933d2c7f7f1f105e2c858ca55b37f88a98b9d25db6cbfc4ca2b2abdc6e9ede28e8cdb4f9000a48ac4f30ed80788be0119cc1f3ac59d6e0b6bb5081a57a51fbd079;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1522afbda151c31d182e8f222ab8fa5c41795593fab89dc099b916f9b5623a0de0ee1a7757b0bec37f5beec0b2a2964d3dc647bf35da66f41e3bce854c68005fd82f1fb29724a1dd38e5b20cb53926ae1c0cf93cdcd9f35419139364c73929f02a8002b660203d1784eff25dc860a53ff8b99dd585284f62b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a831326d272b49902d037a9f36131f93191d5f02948fb9ae6c37a3e938942ce2682694a67e9f7685c5ce9c43713d7e7c92814a906361b9b78ab119d5f008a8adcefb83bf2216ddb86a5e50d76d6c25d78848d3a2e0064d19fcde39489a39001184695216beaf7658bda97f7e74e85edd292a6efadc581631;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18b35b2cce033cf7cfa32364b735a611de59ee0ef143ffd72bc6ffc5db123f45ba84d3c30f4902a03dbfc5c9493ab11ece1471e10183b172acb5ef6a3b868c5a90d2cfdfb657391fd907c92a042b0c4e4cc4f52ec4aafc6bcb7af471f7d02ec4fd94cc0228b39a7983070eef7df860534fe1e3fb8522d0522;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f779c512c49e5600dc52d772fc473f89000fca16fe126d0f5d0ed42fa15a0316736fabfad7a09a8ade0de969abc6bf4eb441a8e7b19a536b75de6a6e96442d82a8bcecef659835ba9e0dc32ad9974b3cce379317a5385263369a2fc899ddf300da27a0c567c44ceefc2896afd9e7cf87f36445b7e8c5ff4c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c700bd666286a9b1083599df4e43b66b0ad59e31c074312fd71a388608a703985227cfe7e70e724363b4efba066f7226985e935ee3ac8eaaac382a8e4d36012dc8edce41e9e6dcec944f6f5d82316110d19d3d331232e4410e245a51886fb3918c479b1cd4908928e58f371aeefdf65e062a9c82542e3091;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f3099c6f504bea8a137a48ff2290a610bc233ccb7e250d4054c066ae592c88deeb9ef7d70a95bbc2369db0c4bf03ca600559a0b5e390e407e3e3e3057cb3b1687aa93e31f94b55bcb131a02144e1dbfece36243e71be27b3f6d7ac9656eb40e5306cc7127649c9337ce5f47ed2545c1b0adbabf0ac656c4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88e940d97ec3533af63166740d699b20e56eab3749c3c4224b2034cb9f7c0f579fb0d089eb3ec5f816c1d36d8f1ed7cc533ceea5adfdff7179cb7f9c362adfcf4f480bfbd5aea238b3c2f47d949e934d4806ddc313b785c2bc27d5315a2c149f80e543897409ccb75fa846d9c9d29af08f45ac3ddaa3e187;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda60abc890789498250fe1c7a9f1881b176302d08e4dbfcfd7a37ff26b5bd31d00259f79362178b77a372055ac470fbef8f55ff70a25c1410004f9dc1f4369ebc4c5181953d2e3d23a2b54e34bb3e62365ad716669014e660f91bf91d9fcb090997fb5f4bff042077008b3aad9562a416c1aad24560d8f4d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6628d1e92bcaad96ccb71ac6adff56f1cf09659d88abca3060baf6e8403f6bc0a422c8acbbd124a0ccfded816822533148a6a6047e06e642f6bdb3a2222ebaf7020b23d480e04b14a58eb9890ffe206812fd78f7577afbd33eae5186380be08e2581d58c4bc3b687fb9768fc2d7c59cbe3675999ff5da413;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3cf0a5bd0b1470456ccefd6326a3e6edef7441c242d10633b26b1019a2dec39179fc0c23b39bc95f1222fbaa1011e4f3e60b1ab0c80f4238c7b907122e89850e7d4c14661d73a0c31afa587b82d4daa1b4e611c8f038bc538d158ddc2a184e231ec6cf5e1c7671357e5467e6cb3f2a0234dc213da8d8c7cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1b73d8e290d187e30c6d3274b5def68879bd98f9f69b9076120f7eb8391de84cf440ca2bc53989813999762098e68198cf07d5a584ca280e04144b8965fe726fa89679ca6e503878822f92b33f24cc828b338fff9b90e8e9e01e9307e0a831914ba0e847f101552a68c86b56e6002d4dbb3abbb7735ac9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h85c20b6ffbf60acc6e3b55a0b28d0bc0d7a08bfbde40fac9d8ae072c6391c23813bb58a75811227c93ef822479f7531ee0b10b827fe1f23dcba41957015e8047a1c965a957497a60fdc3b4b8c26fd00ba5fca3a10ec459f3818892fe68a73d7ecab44bfaf11eb06b800d7cca36e39d1e1a85cd8940aacc1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h167f56173cdb25d8a01a019b7987a2b6f363fe34a4accd699b258d085d0c092d1b2d07755df514a0205d82fe9a63dcc3de0ed38246e4bb10cc35023848eb906f529e245098b6026236c4b1e6d927f7a31e4e223a7420edc6d6d2d553ba7025dc66453a9947004932dbb0788570646c98bfa8c8e3b1ff46e86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102dd63a469ec5a66ae4fe79daa49e2883046b038707f766910bf35eceb5411fc910d17c26033932eaa7a09272084bd38c513c6210f35162d10937ac0629258e5e4129c1411c4f500afa7654d1e0876962c3eebf8fc4cb1f66a11614f6346fe7c80f17f8909c5d4d8f128e21d85a8754d5d3dd8f0ea6b6f93;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5173b0b1700698a653e68721efd4a5b6337b5c9d09ce141ec55139557cbfc3cd202e12e4356e86e9e7ce11deb0b057f2c95bf8705609c31c4d0f393ab9c727d350d7725a9caabd9fc0a43348798bb54523124c8d4a43cc1b0cc0a6c6ded7e711676cb7a7ce337649f102115699621ae582986dd1863d70be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h59b6f3818c2829ced0647bd48465abaae23172e7296e664fe3d443061ca341ce754a2f39f8e344d414f861870fd8e0b2e02792ad0a1788bf6606812e77511fcd732ab13114068a5d3a45b8a2b9c24313af949289ef41613031f6a010f37889f9b2859baee2af8174b7682f5d05a10b7a539a2597d1fb1054;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ecab4a59a49ce69c6d122f7b51f03a065f9f5c3cb2710e1bc8a0554675108cfd6241d50a9715ca8c2ae655a6dbb1d9bf7aad7edd8807e1a6f3901097b0d31a3905752ebe565d7b91d7c72e7524c3a45dfe9d3eb5c19eed728e498c400ce3223ebab819c98450fec1e99871099d371a7b40345d37d3d9a3cf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h96005d4d5d62984a6efa758b75a58b60e1648a2548e53306b13fcc9f6bec30a8aeba44dd66974255a247764f66f722d1c5025bbbc64635819108d8b408316002698ad4b2bbf67e39d5bd9bf600570df02c42442e0eb18c9f025b1e0250a4013717eaa7fb22b65dce9315ae635543420249897bf959d24114;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe0a59dc92728bc5c8f874af999768685e209d394706e2bcfb3b5f3b86877f54b0ffcee2142fd14fd1e7411f23d58ec301622172a96cf2f66e43510055b90bb08f9ca88201110fbf79f256a98840f61cf4f9b9640a2e63f5fc44db567a0e5392791a4c27b1d4120ac10808d94242dfa6f9a000ce3b6c92a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aada86fc57328c72e174bf57cbb5699b3d6220b78c52c01ec68ddd418e61430359233d1f474ce3c01aeb3acc771ccbce7b3867eaf7ace47da93f58b1fbac1622424ddd6ac4dcd4301d954a36e8f478a3a7e131c5037d3245b93ccb7083bc352705f6878408857da3c04435aeaa4e1a020cbd5f61f52f76e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h50c2dd06462d4fbc774cb846947989bf0e2d996a5c678dd7fbad0601c25363fbfb9cc094d322b7cdecc3d415660e221ec9fb97067a6954a545d74a51d5d43a5fc428d210bb81dc9cdbd228930526f1f01cf53da11a733e83ea06545bc252e74c7bdb8e478d2e878c272fd54234a315750d5fe8267c282251;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14636c4bbe0541c82aa6abd9b7d23b171c827e82ca51374379df557fc9b281f9955e86f035d2cc7e082d4b77238187f26af026fe7d3a697ed2f93fa8039105b57603792fbbac7cde9c28e0f305b41227436be6c6346bb9fb073c468773439681dd94218d047ed324f172d6b82d452bb6f31169ee937e23044;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cabc93a4d39c4ff09af3e8c92a0f0090de7454c2025a58b467201ade7bd298a621b9880c8c6ed9feed2cb7db1d1f4175b6b7d67d3b350ee0729db3660df3e566c6a34b92b2a0ecc15e45f994c7c15f3fb2eef5c5c41b608c78c7fde00824f27cf003ba764c5c28a64986066e17109f4e2a718cba4f6fe8e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0cd55ab1c156b02cd20751e4d93cb76dc70191bb617eaa0bc551de2cda1c43adc9bd60254dbdc04c2dbbe091c6e8656208c384226ebe88f71fbbc85d506d70546e19d52fa0008069c0ab1a0cd1aa370905ffdbf36f8b49321eb0b27cd95c9130eec7c9760001a32cde43be29cf03119af45300ec8bffe9d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ab41e313cfac13c7f8fc6db69b5a212bbe63a9db0f937a8964fae5cad882214b8c811295d99991a55bab907766ae5f34597872c8db4446a2a9f7a99cd567037c1fc4613a4f964eaed20d79267501fdb02b51a48ea89ba5a2a42bf762d55a40cbef3c521d1a111d4f3d4b0b862e36e2dd2c6a72091bfe65c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84a07f769742c905732a6be7503ad63355bcabb1d46d41fdf272e75595182d4b59ccdc0b75c9d5848ccc5e2b5ae408799f70f61601fdba188279c9f941bbc4039291d1d51c2c598f610bcad70635860e3a43137685aa4fb9f4c5bad1c56815d9681cb1e2fc25cef7dc88088b33ee41572d8246920e8d5247;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h36d58770114528ce45f50a5a9f6287daf25569fb630629045d1f48efb83c3000083c47fb9c2d4b413849fd11eb42df7c091c1c92107bd89235f45b887daf2727932506e5bf5f991152ab441125720406f7c1e9d33e96c5a7cef92cd3957c98c30a31e1e4ec894660e6b8a3f0703f623aafedcc1788cf6c28;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h300525e70bd92ff5733c8151bd031efdb05a491c962ca6a26de3277efe19c4bd64b04ecd7c52ce7c053b45b4ca56a3a10ad15a7e171c7d72e01ab73a2c4c6d3b8244b8abae4ae64ba412bcee2800248a5dd11f961a115cdef4fa4462116d8194aeec57056a6e15fac7c635558adc710fde5789336852ee22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7eb7876d3b8abf7c72ad97105a76be13c04e75ba17cd103b55350d79a0ce5a26fd104b2fa7f4c5c0237230f9878008d4e047b95e09b3af7f6368fbe139967bafcb576dbb8e36e8f66bc9fdb13b014e05b1506cb541a334a6bc21bc9de8d71d3975d50c870c40bb1d66826d8777ab0f4dc82bb0ccc06cc6f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b9b1e1f5ce70a250f3de219bdcb23fd8298e72e2373dbffd5474299cdb53391a612a4f4c8fc2f5553faa840a8e0c7145140ade2a260ee1c4c95627d434623c93462bbcc817f359e1c8f71c3b3fca3aebb735cce922e41b922be840e1a8605102ad12abcbbd77b79438a1a79b2e7e86cc33abc779614ecdb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf44359bbed442ecb8fed7efe1af2d6a170e7406ed6f329e8b36e039a9610819aa43e332b790699605c79842e116766c6698c2b24236ecd5a82952ad682bc30ae1ec6684e399c44db205ee26f2ba6c6d2dc6046320b88977bd24e14a2c620436afeec4782b557ff29880fdd0cd6f2cee58571f8a19d8330e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6dc0a4977ab163e07721d6767302a811b2a05bd7773b79dc951ac7347ba53b84a79b09b0c2a6da163ea2bf1e6335be3d86a06d94a4ea3129400da14c8b5022db2936024c69405d29c7df881d4d0f116a9fa895586a7830e6da5a58b4288806df0306fa151c9447cc71aa5b8d2838bd66990c777d7e5102d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc20daa69edd5aa38d5ae440fbdb0f32c6cf2447745ec34aab5f340cdc917b407d6252da4c1ce450c983573791c69b9d26d5a2d1f4e0da341a411b184a0cbc4e90fc17348f30e027cb526ff699ebfd074dfdb06c6b523b6dcc0135f3829672a33c9ac2b07ecc332efff4c647b5f2559287bb34646d57251f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c55bd9096b056ed80791663dcf27c12f7a2223011540eff44ebe65e4fa2bcd9679ed34254ae805ebda92c446c72aff874ba9bda55c99fb9fd60de58e8568ffadceb48cf246760f479f84b6a2919674e0eb15c9975529aae6c4c832571a00a907444f4c30c0a399541b378cf958053adbb787ffc197e9f0c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h182530af822d8747d14c76cb0ee27d747b4beb4f195ad73c142450b20269a193423b0cdbd47773aabc8dbac56fd9d6b16465e3d4b53a3f976d3cc9c0fa0a64e56918b53078b8b314968065b7251aa7edc8a94273338fb9d089d8ee09980b836031ec7760352faa5788370fcae39c1b65f8e810556bbe3bdf8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac0aa6465b9e0d251829ec79f228926797a37f4280c9530153f1d028f05d46917dd06d6f156df87c9cb363c9314e8d33aea9db68391293078f2de2a0913a6f73730e0f58f22f62689d2df545497632e7ab5255ec009c6edf4e155c91b13817f29e8336d01e3b37e1a2b01d2220c0115f3d4951c6bd18d36b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd93dcef0d5716b98b9421692e9478decb73b0054f7b118ec36aa4d457ceb0a40c5831572cff827d96ad1137d1edfb57d55cff28a965210973bb6a29442058e1c9ef8d10b63f5825c4eafb019d851d99e20990f29b8c9dda500182cfb3e36e4d138ec786a8f99e041475543c44bf59696d16adccf7a37bc5d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b9c863271d4544025d6dffff51e43ac98cc7adbe1af95e0bf3614d0b157d1d5fc2bbefd504ed5dc821f6bce17a2e8e90a099b9326d315fbaacd9da0e8d6eb5116c5da0ea890146373d02f394616eadc03b5428b987ee7c7185e9bb2836f4e032cab31b8cba8da06e9e7a8c984b8094b89b0485c1a74ff5f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd79eb14e8dafbfe60cdcb5f71f9db3715ffd15891ff641f978a0d3b3188684695c3567d3ef0c53a2afc2b50be1bcba2fec2e22f26e50e2541b50d12f0786173cf4a93a4caa2f932910cc0ca7acb8ea04a7d466dd23a3d8b00a685a8cddf26309999444eef8b18a9fb5e6bd31b98f64391e24907cfdf16e6f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b22e79ac0ba34298faff2659843e3541cf91978fa5d57b9c8c32dc73bf2f18b37d5fce49a41a5fb19df30a9e3f687dbffcf1ce79f8a9371446ceceeeb39f9f78a886ecfd9bc114967d51775d5126fd05c84e67e9bdb4390ba51768a1c6ea6ea0f535b79cc61bfc3e173ee7efc104e052c137b0bf9a58f04a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h129093a408a8d19a013f93656003b81b71c5bf76be1744a58eae07f8cc8cab55f263901d382cf9e5472eb585650860a3765ccd7847119e2c89ce2dbcb3ba407572511411133639dfac452a49da82ba4876203b5573ad61a9f695a834c13c542e62a291e18a1f7f0406a7958c9f56d5ac5f55617adb37a696d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1301d64555e9bd60d76a4af7761d6275a8dd31defb7651b781a15d59127f7bce54fdc94809dcdccd99f2e73c67ac72b1f4c5701482d095a27d8d3474c64645ca4c6a27df895a878efd7fe92c2810afe93defe3480f7ff8874d6c25cfd40fdc4d7afba16c8fd5bcaa2cae062119882d212805bb6f88b241912;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1af23c1cd1ae84db0ced0946d7ba5d64ff9e018a526f479837bfa1019a406cc57640432398d213c23cf58f56369d2b025df1ead958239682fc7107a00b54369d83004f6fa89ac407a5738c46e00c41cd9631e6ae160f9e3a4835e5b2c1a42af6cf11683db0ee0b45e59a4376be3bac852d3a5574cc8eb7863;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13fdcf68f29c8a765e95405464264bd1deace0b8ac6e951a69ed03b7c47b3c94a959fb86ebe6a6de9cf84720461620ec1bb7ad7b08b247c733c9852a0c75d398cb9b99c0ac79dc96396dffb35549ea3e2d33bf149ff8842519ad0da4fb898b453543b8c844ac048f2f89cda7395157ed06c85a06f7c49e0a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa00794074a9dcbbb302db69badc89442318f64f3c917f5564daff93195b2c986f60fec461ff80df870555aa575f2da3e2c048b22ae36f6ef54df0f4f5e06a78367c9e9110b83c69ac28333fdbd51fcb7084f087a611badd3c0e5a41a238d7f01887fea5a9f6e7b8d5aa790a47001db6a644ec8b4847856a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h894514782ccb92a47dfd5dd08d1cd36fc295104e7c3922213fc406ce65eaca6c183f99f2f680a140f59dbe21656be841d2b78b4a990ea8ecb425ee74eb21da0fc2ce2001edde2be10ca15218e2fb6bca19816a0ba01d09fe281b2f2a058176d1c4824ffcf2db53ccb947a3c9284b9daa4201ec6974ec1346;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f82ae08892dab870be67d39cb5f28bf252fdb516a75aca59ebd9505cc1f06e6bf479731b8209486679f8400197f73148d2ece3011145a6e80b9209a1aff29c1fe320ac08e1207a126c320f545c006a9a301fa064333d0caa7f53fb9744ad39a205047d0fa65709e56f2580559ffb3b00c65b568865dcc0ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d24317a2a825eedd532c26141f1d007e48e1118eaae15c3ddcdd95e94af6c9a55abaa0fe4532109842fe466165aae097d7dbd88a2712de7d751b708ee813f790d4295cce026215d0a0211adae65e86d221d74875b4911e3be6de6c0fddf275a87ba303712ab5f566e042aca3154fbcdb4e664c1fd29dacd5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10c5c74b2258b9a37e13c8755cbab9e02651cf2647b40e085ed84f0cfd3fa21ce1df3a40131748a9417328aead46a4eea84ae1a94f832bbd86cf0fb7d90ccf469a98b449b3836e516e56aaf8ee8d61030679377db54d9b56b53dabb68a8ee57b5bb2a6da3490235565ed41b59b332ba0e9c92a5fdbe77f504;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c43ad1adb8a3c9a8e967e830c17b44167757a7455bbd6f7c3aa45b3257c53a1a4be0648b2587660c60a1961b830eef1b0acf1118399b77dfa4caf46cab2deb73b606d11b3d532b376ba9db29ed37091f309c5bfc299aa2917f74ba9cbc788d1b7379618af97a51cf67ba9b4406a6c423beb9de661775196f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14e57eef4ddf8b8463ee99e592d7a056d5e525714336185406e1bc75a44a98d7f39a0e96766b6d859660db15b465f200783cb7e6646f5de559074e298b71d33699aa1135506517135aff303ae50a15d5d122414426ef5a483839ee743d5df076d2bcddec9332d41e0258c55b4684fd3dff3a6595ce53ff212;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13148b8072859873703258df2d8d70aa193018cdbc766528985d8554b4a917e5e6babf27d19109c3663235b15cbbe4eb3a2b118b0030f82251066c4c24b87f7a21b84d8705a0b0c09e643c14689abd8a576e507fa45b322e46e215f30ea28da1c16d33f8c8c1064ced3605d333b63d16b6a788b4f854a58a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1122f2890c5f9c02104ae633d153b9e0031a75f2725fc4bb80b106f9a4577845f8b73372978018da173737d5f677d2a494201a36c2d46a55f8a44f1999771263491e139a1f172ccc779b1b8c0f12d8836dc8f3bf9e0a59e11bf8d704a0a7ae5adc2f1d111aab4b85510c06f3700d38d3f42ec6afcdbe633d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137d92961ea17f4ed235b67d35f165a4aeb9564f7ccb7561f284422edb4127b149adb8aa33c577108ba865f00310defc8c44c7d18181c890fca2ea362951ae30ebaa27b3ee23ec129a81e7a27e9804d66d69111199ce5c4bdaa3863a6fe1aff3c666d86f47262c3fee56e6218d90aa5d87c458c8843bb171b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d281c18130397d8b911d251def37ec96ed8dcfce0a64de76f6f94663c753d4b1d1875dd5885935a19e6cca7d51be4cd93cd46011b16efe400b10e64717f3b14d98374dd2dbd72343dd31ccdbe0c3561f73bb4288a57c18bc966f05e473725028543a8b9d12992d085de41e6ad356237e02240e059475b1bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae75efcf838f4f4622dc960b9448a2efe387662a516e936be1038cc9b02acdabe347cf699e07c19042995ff6db235ac4d19ca83f48afe0d8adf1768083b88f225b279ec4ad3fbb14737506faf7d4d1cd1d027f1d6faadba89b335f751cabece2c61fd7193f66301237ad02b473f8215ec9135548ba2e1854;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e51c3a126816d5ee92f7aeb7cbc4044427eed88bf00a5b0142b7e36ec8aa59833322361a2ca26ead60a1205394bf5ce533c1df13254dc67a930126a9739a796f1458c19306847464423e927a84826c4b60ae6a1ad19fa880abbfc433529a5d4e12602f8a19494c713ad78e746556b10cfc43de73723de63b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h176e5e0c0f5e5a15518f873e55d2f7a3f395b979c798ec42ba0acb53b6079ac4924aec1900f0519e48c984d0e0e8e9a6eb108e5d6d8b5b87d366f26f02c151730109f2e779f6d6e01eb0e767148e1de492fb2679af7c36ced4406186590d249eff4c71936e0b5a5f69593a8fcef1440424f56f7d38ebc3992;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d4c8c722a5f1ffc6e3f91e5a67fb318d4380e0fd453d2ae9c18c1ab55fbc77e6bf0b338b9f9470ccd8a655109264748dbc9c0f5e26ddb463ffea4c1290c3dc1db8a65bccbabcbb0e83c58b82b345c8ae5300ca29c9ff95e562f829221d6cfbea28b039b1ff27aa83f80a7f6f72face1f02f2da982d9b90c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h368e21978e66c730d6ab5fad6954e28b5592458b50b7c5bffe690a75ecdd3c19ba52e5329245800b72880245f26fa9a1bbb0eef584096ecb61d9213eae5294dbcfc2136d2e2cdca49e6d781cae6a3e2bf4544b3f23745d4a87784094d7cefc41edf06ff3abe2ad46f57e2fd2a1836e19ba8484052ba6c9f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h28731c43d5b585e41f0baa971506b7c948214d570a7a2a371ad62f10738d297396dc7f2dd7f1e38e24177f9a9f7a8fc60a6da6a73ee05c2be09ceb53e1297c1d7d23d0cf12ad479bbaf83fa1ccca7ee21c365d0ee207c38f31dfcf5dc67fb0227e34f04ecd583e625de2a938342130aa10547bdc14e7c1e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h191eef274de53530f75d151b4f0c4ff4fb0efbd830cd6ca427a755c7590618a87273a1f8a01a5c8541cbd97bda3c7f476173a42f6fa7e0902f19d0638a5611d11acb84ae40e583110071205c9c9902fd60ab17ea770f754d249cb2bdc781a6a85ad9e0232724217771fc369ccd6437d5d7ee40555eb7433f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf96e380c73f30b17c649e82b0946705f5c17f0d2c6fbe59174b0259f159ac25034db402fcbb6640abf7dce4c0ec65e9584c055ca798cd16c9fb8cca2681aa4955d7ebf7c192ef33bdc916efd1a8fa437b8eb14fc3bb7e612291db6240a6d340d92c8c50b272d851643510047cf41cbab4b22debaf5c56e00;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d7e02257f55fbba096fd16246b71300fe2ba13e735c27cdf2cc63d6ab86f0b4625f73c19bd27bea0318d564f94285b34bf14484e242c2a2e9595a3c3e756b83b3f903f51f498838bee4af7c38a9f58df0a33f7ae068856d6b1ef74592fb02e3fd361da438452c9b7ca51785a6a524b90ee429e64088c561;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115336a097760dcfe2b7d5df13d9d3bbd7dc3b38f79b931f1e8ed23cfa8be49cc56a85147cb51b90fe7e2dd9cc33302595a80b6e61533b3affd640998afd6eb16ba04dbdd96ec317aa22b30b517f084658d4465d86761a4f0df9955634961146a83337b0b343d9401dd2272696d29ef4f7fefa96d5e9ea1ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h57be1de3e26ae718f0f97d14289ddf9ee1bcc2fa36a5ba91a63a615d51baca52d6f26a36120ace041be19cc2a149a7c45d3e96b3de5de38418251c0e3b559854e1889a41d4d66db1c89b4a1ea057f8b67eaef5374c6147f3dc45b967b6c1edfc66f006af9676139172a0d28a56da44efc832f5dfe24950b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b9a413bd1c517959f47ad32560626b9912de00fc25fa807744dfa376ddd9e97ee4fd34f057c7047ed58d35d2020f0437c28d04d894e8ec70914f6afa4b285e109c068e03d2c682ef85162a4ae54c139cf9b01b3e33c8dfece99610e1133c0a491021f3a5456dc6857a602244ef6febbc47f60ab518172f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2bce10b81b14511026d4af8c36a9eb98b178461cba3ebae7a8bc6547511b7b3561f358c9580140c4679e3b0cc420c2a4b72748c2994be95d242fe999695a7f2a2db8d956231e1b366d92039f9c3ace5364f596a4668b6c5a73ef869ca690a1229e3204d2086db2a51925e6aba8ee8200799dd2d672a748;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he93dc2a7d8521aebcb06adb09cec1cf8dc40560745e2bce9fa29d93ac42e1a54e93c2cb9938d8aa526bb923ebbb822a3ec797839e2f7aba76a2a0f7ec3aa40b568d6f5c4106efd7ad94ff8e4fc8e0e39379d1e171cd022a0de6e432d644a200706729c645f76ef4f78c166f8c96cff259271d6f00583cc57;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14fb94a8725956702e1643faddcde4a052e5db94d3732b2a41b68d77be2d8c0cf632eac96fb708a0773b5acec746625cf0a38fe7c106b721d868b55132ce4610f4e2383df419e812fc4a1f401f21196cf2b396a5fe74d079fc419a8b8810172072617887ae50a1dcc08a0fdeda20abe7d0a67429ac5435e66;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18fcff50b6ac88bd567ca7ed8c1a1433d2f5d10d6cbac23f24a51dc5659ed9b43fc0aab5d57d7fe93977011e8774e90deda8cc75167658950d945080fa737ea69006718e5f2672f6d1a139afea396c68da3f8c360474ca6054319121200302cbf2a1596ebe622728ea5f84f1e76672712d8fd9fa437b58453;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdb1d05432ff419b9d7b76288e05b5527e19c1f99cd14967a69535ecb4a9bdacf0121cc84abffa6d341cdd3d1e48057f181362279ce7d44507d7ef2e22d4dbc60e81fa576e34d1a675e213006cc0914ba18ae5208ade64a31b5b14bc65311e8441cdb5f9feb08ad089d3fbe84c1a0baa670a8bb6339237d23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd04f151a5f3c3f6d86789b3c997e9ab8cf6a2b7b5a7b021fea6b9277f104414a31e482fb7cae595f259a6a5471717f00cce33760d638d650ec154952c700e1de8c6e45f9e13a645fdf6c704f4fe8fcfa6b482e7eb92ef1d73d66eb6ed2262ef6748ec4f8732ff4783d032fdb8d9e3064ac0eefff165554c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h464b1eafed7e5aaf61c140070681bf461da25e8ac1dc046734e510f4e9d1799041d1864fe6a2a02112a2cb55a950538b7621614b56791c7994615fc8250c51eeae5d78b13b7868ed0b8d8188cc648c915c89d42f48ea18ba89f9451bb65dfdc63b86c37327500767915c5e29c057beb376fb427f1d51d972;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117bf1d798b5f8a3432cf0fadb0eeeb561db21c0a656df2734380e72f2ae5e8d36250c30a66c9b7117111eb59ba232f7dcfc27a3f3b113b158c4735a3e2e571d52b68fb84e193dd2aa79c7b8f33a0edb737a5f0eccfe029166e16518f7131d4b030716f2691befd5a94342ebe7c0816f16ed2ec6c7aafbbc5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6f050dded06efdd035feb88b205c0869294e9220200c221649b0ec3a0ee8f95c4e9c55326f15e8374cb10f6c6ab97e969c4635d347671d4bdd93aef611473a3ea30752a368fd34b772425f42b1c0e5af5a09a2f28fe9536f411dae916cd05c9d997d66e81a70fe1dccb6ba8730446170e1eb86ed2b24674;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc097dda8a8b3ee20a734b488dd650f29a7fe1ab1791bf7b63ef139a1cf6142ba75cd929b572eba6e6b4f1eeeb4c6278fe39003e6ff8d21f7fed9194afd29dfe4a70be9de36343f95f277a8a268a0bc2660f854b2b3448c09d1bb3c7d56456ff4b72592d4e34a6268b021eed44d350191ff1aac6d3bb942dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h701e2c0789a9089e0f2f7cc8a0c8650a81ad7f5c95e2d7c9a390e6e23f9c5d35eb2527e70d0e06298cae6d5aba2492f2a9f4bb3709e7bec874137cebf508812f57739973e3d4324ba08b34d718578b6f50e905f2ef741f6dd88d8d0c2f5cd51522ff6ea91f104610d9dca77deb58d11da26a032a6cdeba6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfcb498edf9db1cf254b487173020c0d8dbdb8c4b3a4f0c519d139d9b23e165af6c643f2ab05dfd9ac5aec3e5809c55eb524620c52a00acd0a7f6abcdb97a35fbb80c5c92d383782550876c17000ee7a679909e5393b858143b41d456dfd2315b4673789ac6913d3fd56b6abfd3ab6f406b8c25059312d1fc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd9360ed8bd29d7a58be98fed0266ec0ce0cc402c9910df0cff52517b2e3c7612e1063b4d744e9f2e081975f752e70c2c706f4a8b75d09dc7464abcb916b6eef27d3afb6feb0a293a10ebf6262bf207326e2260542303124078fb1c1cd73a2ca6cc5a42eec3d831419db82d80c4b5035a0294f12ae67f8aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h767a624357d15e5a6860b1c931458541b60cad2fa8a1fbe92853de563afafd5fb37fe8402b4e4cb7715421d1e30f11d22a34d5fb03b6283551f8ecd1ee484b8721b1b113eaacd475acb31ee344e9c2bd158039e0fc79bab7dcb47940eb13c231bc2ebed959418df7ee1b2ab5e2e06011fea18ecbba946547;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16092e53b3cb0c1d6a22ef6c933cbd8649a1178c0b1e9e0b9b8509393822de51f5b66988e0118ebf91448ba4b529853c2d49358fbc363858f78e8cb66ae6f000eb2c459c176ab9198277883d5b83595a94dca00089bd661e18ed14337e938bcd27687cd95c9e93924de903cb37a75f5909f5aaef58008314b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hadbc496afbfcf1915dda923ed09f84ea36c5300c0daa73596ea120f04df403e7619f59620668ad255f1a536745f3ce3ad5f4267948c82bcb112a2d01330eb468e9082e07a48e0d9bc732467c2d1eda3df70afa2eb2964d659d1c935091478a3f8849434108cb0a13c642e897cb71f8eb205c130a99fc729e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa26b2e59adffb5cbc833f6ebccbaac88c3953bde33363cb9b4e0fd4fede0cd118a3bd489670b11d381e81519165513a23d88fe6fd40ae05110004753fd5fe805400882f964a8c8b12bff3d8c7302aeb16876ba937785b9a50e98e575392be667d5f27d789839e766ccd22283f6cbeb84db593ca89c129aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19a7bb5fc5675389156ec6faf8424ca42ad84387d925a5e495d35c5578fc725e2d808771af0ef98d7be8bc66af1c946774bfdea9b433cf0f25884a0063c46366e43e9cef32f4f36cefb06df5180e5de6e8a0817cd6041f5506858844b1618c022730eed157db62707613e3857acb516098f816a0d81514a23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1671c1abd223ad0c692c8f736a71af270c70bd04c9b6bb7be3ab8470e6d9a803aa57631475815bdbc39f9fd8687c6addeb274e3756b716eacc95c1e2308f56a00a5eeb6bf6c590e258cef2b7c0deefd8c1d8175b19ce0d202813f070589879d0a7edc33e88330a0338fa247c24e37b231981e56d06c043;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha49815e88d7881bd8f5f2f320886573971d8290456d9070874ba24155558104fb54020c2612caec20a464d3a10e3552aae34c54a8eabd090b6f3eac44cc3295e9d547e6e842787d567b839740beef648dd55f7cf5b9305f0b2eb0ae1a050ca0d8ef9bc1c9f43eab9ba99e71fc6bf62f13b4bb9a14d30e812;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61207f73db73783f7a27635396ca07127aefbf224b540ef185572fe2c27533fbb90d7af9e484edbb1771d911881e1baa0feb318d6e04a7ebe47022c3042b4b85ce2da3fe04baead3690a377885eefa3097130b9fabe28f39ba1902a9bd3d4f956ba8a504abe7ed4dbf44c83d52ade5c6e3d23971a85fc592;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f2bf4086a3245950ba573819249319b22f2de05bb26223d1ae68925281773915396fae83667ed8eb2a35d778009d002570ec9fe34158f070da7913ffa5758e2d73a75161a8dce56b8d4097669dbe40d45daece06cc1660ec9491a6ac157365739e8fe8f64d3638e493d04963a0519c7a33d55c35c174636;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1663889d405009c2fe3f18e9c7dbda670d755d799cff7ced8a3fd49169e6d62a2aea43a1649c0eeadd6366f25bbfca455ff47ad9f5bdee63a1143b7c6611c1c9839c617e9d60261150da80ebd64cdf1553dc66f74e3cd6aae7b1a33c6caccb41de5f1d1d24cdf9b0b089c420fcb1d6ccb19f6d83b0318e391;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb7fc15369431237e399d4ed90be634086e981d0893e936b584bf416cd088b651e7e6c8128e047d76ce953d3d1544af9f16778e2d51f773c7a5ee99885ed31be8760d64a25c888532535e9395bcaf7f78745decff67d9a9b9ede27416a49aebbdc206fdf19bf6fa4018379dcf9721f15290c23d776957f806;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h948782a0bb73811f5f02490e6c8395941d2c1260f8d42599b230044df79c3ed79cb15510a165aaa4f5f419a9e9dfdca4fd0f4c18d94d0def5d32043c6fca67c144b22b17efebf3c0661905b4c74cac65eba45c45361cbec23ae55b132a6dcb94d9d3a618d982143a3a28cb13bdf8a7a3197d985a2015d9fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h781dcbc4795d95b1f0728ea74e02fea1b9235f96a2fb0c0d2cd89b0da3e70e150c483bf500a9b5c837042d0c3e642e5e290cfd75c93b79b72f0cfad177358295c791eaa4fe1708df5f351f677d2d3bd2f94678c6ae5f85f22c3eecaa3c12658fe927e51199081c3081371ae6b20c5e52967d770221f2915b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9f08b54aa8132cbb209e0b0b9a23b8932f5d05733c7bcaf772937d52e37d86e67f264ca9c2bb9939cb046ca51ad060d62cf89e289aa7e702a320d3d0cf42e694559fe9cc0c075fe0072645eaa246e45695d611263cea502e1944ecefb97f72c64b5dd2a0a0f95a8945ed29bb07026a7ec3e177986107ba92;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bac4fadb649876c74b7646f6198d71a769116b2250db368edc16f148c587cdd98d197eb956df1c1fcd00e06a57cb62b3936b22e278327184edc751531263afc2f7d6b40ad8fbddd5a9c11cb367f8105ff05a0d106ed92d985be3372bb2587a30fde47bfef2dafa618a103483c6228bab673556b5760e49cd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4c7475f7a6fe3998aa98b5bf434c3e7e59dca989f05a3d25949b240b03c035ec0a39eecc2d79714d73062034b14104bde4b7a8111ded0a7720c6be0ef5acf0c0ee14541bdd72250519f57fd4bcadd85d3e747a81e481a1cbd1b7485bbfd9ef407912e495a3f98d78dae5fcda2752fe05ee6b0c76be7d56e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd21faeb28edc1f195be957d960b2e890377a6a2cc2efeab382442581af5628bb9608cd53a31d1e1a72ed54d65b3ca0652d9044a6bd3a55b34d6cea97760e7c3b94bfe1b2fc2b34af7d1d1c47107c990c983ff494803e942c9c192c7574d4b7b86b018256fd72b452950c501fd239d0e2dc4d958308861412;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e4105520e50cfa662380dc10f7ff4aba5e48fbe15ce3e701e04aa1bb55e2c110ffa00200ef7810c05f111a28927e7744e361580d70e645aebb2c2a469c4891583f1790677c2c388a78a976de9de651a23983a661fa01cef25472c7d1f925b254dfe7b2cd4faca08eb131e05cb7c5d48ce1ce80a3958e8cef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10bc6ec75a9e3fd0bf41214df36e5551dbc6931954c102bd3d9f6be11e90e8b562c9bc321299f81802e6ba1dbcd2d3a50e459d60e3ad51ad31572b2858f214026a1e1abbb2b747df8ccfeed34665f1ed6365eac1b30454bc9d31af88bab5ce934f37091b0bfe8d6a7cf53544ba77c3a8b169774578b4deabf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a6d9b69c1ef6701a96ccdc5cd1a2816f3bc3c1b21b61a914af374890ca466863f72c00197b8af76acb611f704d5f90b383e80c0e5baa9048320664ca6ab59191a894401f54c1866cc0bf1de8e76cd4c0998d8d4c7a3537d09f317f6d2908d31d1bf4becbfceab06ce04868f17693b81dd1c0e7f8c6550e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18c3144470472a45d01194b83f8db36e8faa437d4eea9190d67a8eb9befacf65ebb6040b9766a76558ff4b2aaba637ffde95c8aff53d1b3b5dc17193d9c58326b21a5c2145e25f9b58e876db856d256733c74f51421adfcbb3981e63e7c071efefa88e336d4ee2b8e59723c4efdf036f6815c4b4387630890;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf1aeae31ec800d5746184595b9e965bfc12000f0ddc6db1b7ca8617ea1013d893db9419213c081747b7c185ff9fe6428c350705670128b7118f591c8456643287579efc17f8ce1e35ba43a042cdf43f511890f0647a504665ed1e841260608fa4e5f15f981477ac50fdf1fc475c174d975e1751d7e4cace4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he6772d7336be69ad83355d70454bea114c108d03067d21cc355a5bdcdcd42e740df15d4c68a3974c811038df0846d36e74d840518988e307788bc987c5c158b86da0fce0a21dcf7f579cfc8f64c9abc9c99b1094277c8ad5612d5bf67007d145f5fa60e766a456df074c98044c3184c1429e0234e9a2b514;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7bc63b808404380cdbe7056aad873c24ee6daf4332c75a74eecb408ce2b43c8d436e19e7aad89e3259239b3e7f9ac0e27624892e44bcb1850918d0f0d3d9eeeb18daffa8a91a98578bae5c0d7def7de0860801d4deda2ff832c47820cddce526580e3b76087a32642bce098302c673a387f125751ea8ecf1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h197f13d6a0ad0afd54da93fb1e15993bc1a871b93ad974afc961c9b98aa3f02fc852f80903c29c2562c7cc7fdcd33501c7bca1a5bbe6b7caef972055ef087922120fcb2373879cd70a17c41c672d7c910d21f9ad4d57e6f1f00d99bb567d41e654a7fa9db7dbfdf01e52a1f8b0e5d1a37f3b4d10a41d07058;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd1cafbcb121a984c33da644ca0767146599e8cd9a5c6f3abf9920fafc4660135adb2abb74f8f7f11e3e2d3563b58f26a7b80b6ac45b43b08296d32a901ff899eb3ebd173cdfeda549532d5d5a92cf458fa529dfb22056997286b571c40f8477c4114f35c44a6c3ea9cd42954db74b83351530a68bd1f4068;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e7b581d2b74a5dc501cb203cbc59d6d08254f4557938e2ea45fbb0d6dffe25a1c2a294d9d81e30ec20c516fb642fedb36d6711fafee477afd6419934085a8b697dbecf862cb283a7c9fc1e7d29054eeef66385ea338055e858e2e39f6a5103e6165cb7641417369fe57e81198e9a287f7c9e40f7f0f568;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1990e4b877c23fd45d69b11619506e10dff7f988a6b21f55c82ad759a393954b85ba50c4f9b42db51cd7c211702bbf07e9f16e1ca152f9377e91100e8981e75aae1344ef5c3ea9a671659605d37c981afc1aaec215f11db7eca5e2f9da37c74e211a2f81b8d5f42c7cfc797a43ce110c10d556202e6839716;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17002f51078e4045ac8bdc0b9bf54acbb0f17e8a4f0ea04a8deaa7c239072a9da44671697585fd9e63b2d73b03822ce50c5b4d2bad4eab388310048266dfd353417375ca47392291f99082b93123e367f1539016705759605226acb39e300be5d556750f55f1d8d3bdcb25b9b2661974e126943a5a5a690b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3ff0d489fb381522548f30a2ba7f70161d912487d68f8a125780972d2e40f8dde8be71ace680d8ce0bbdf034244a92c1f53207e5050520f2c06aea994b92ea2e580276df9597f617ac742a8196cb7849241f69e329207447f22bb7b3b2e489ac8aff4af6ce701482bdf4bf2d6833619243213aa3424bc8b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19dbabb97d76cd80c3632d5c78d332d4e5cd7c4b4f5295689f667ceebc261c3dfa6bca07baccd4d1aa8abc28340dc90929abfa012a5fb6a86b2ccc525e4b563cf299ddf46bfeb079c11b23e6736f63af7d1a9eb4af50504de3a531bffbc557cced31a948ccb710185eef22ff2259c89b79ff2f761c0228761;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d4765252e72c2d448b796ba56848ae2d054e42b660d9a379682186cd4e53d3521c2f060d906779e44367e303192bb05773caf56dcdc4cda204af9de895b1f6880d796e17dafef988fc37953bde1eb2edca6a50112d4b398ce4251e1b84ca16ee422cc5c5a398b0012746583c8500da140dc8a80afb32086e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b12035952867b3bfae8950e6c98d24e01e56bd20c9d0c606def90af049151ad568b8c60d6c80598448e1b5f19867ff141153b0096afd445c5dd57d8ecfd02a44f1bdf5b2c9ee24a07b2c42d5d58eb85a2a0c09a1074d67dd96fbc5e965e42c37751b680657cec22c5c123c34fe909f02ffb0a4a29bbfa684;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h144fbcac851f6cdc5abbe9238f5536ebf24cc272f729f5d2dae3a678fb25c68aa83a7aa22b2d10af8a903aaa7c65bf8101fa588646c08cc4a0a5bcad8388569fdf672bf5d7595b4463fce48c252f371da1fb927bc5a87033faf5f1bc6b3161ad0a9c2734f614449b6a170c086a9a95164d9b5ad8772ee39d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h40a2cc59640951738b87a415567e1b5372f58a6e07899b98900c3208e51fb80248d643c87445dbe84ef3dcab1315a789757127494cffe8e5668264efa4acb73f3fda3edfc241ce6fbe6e994441f3cd9fe39b3fb6532ae3c9f80a0221e6ce69091f13a186a098acea4e1b7928f415ef96f9a37ed82233b3d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h331a7ec5b6f34e446471823882d0d6d48516e00bd2b463e69d96b64096440050e8af985ee83e83a67150d1e507c6916e7615dfd22ca0abb31e2020017b4bfaf14f89567d19acec0028252d3868537921b78c0fa3179b8b04996151fdf5bde391801974e25986177b729384626dfa44d80983414b943e6da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haead2291fde35f8a6d203c790945a98d8d5d340b7590ec7b51e467c0f647bc2b94d70c576f804dbc0f5935c31f8d348baa0990d4854c5b1d51202818bb50ffa83036c65191b961519c6916832928887904299ef3d631cf13109bec405a34968f7a98d39e01731434b228cf884fe123d15bee49bc3dede9f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d4b9ab9152c1ef62a3bca08d5633c8ff9aa2180862078688826caed85897275bbf8fad25d5fdfee72b1aeecccda92d74ce2e95bc2342a838452427ce2eea1bea422ba132dd9dce18c9bef30ba56dd46ef536b2ccd8dc229aed9e25067cb1aa136dcb747cbcf745c11e136fa9c599633dc5c7e2ff6868b69c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c875433c9b136e3485a3cf4581d89cffdc01c03ba54fb3be3ec8f13ae39ccc045da64c249f5e8483b3c592fd4e8f6c4b4addb887c915ffac1ccfa14cd890ecb6141f05b56443ba44e3ba9c90f485204b0e9588955a70a6b74915544bb029e47a92c0c64a4bb34a2b62f69cc13f4f75e2344caa8ed4352f92;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc46edd747aaac3f8df584d4d2cb4c67de7e3bdae4b9de4019a33c0724a359210740534e87f31302acef003dc0d0aa7b93c6ff555fa8cbb1bf7ab487566fea3b0ce1b05703b699cb1ffe28da29675ed92c67110069f1378a36f2833235fb12fcb04aec805510a89c1b741eb4ea8e19465966d56825c789e5f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha1b20b95e18fca4b9711b68b0e044f1ec9817dec0738f8fa49dbcddf78782dd3ff94ff38e5f06694eea0a3e215c851f2bcf6f8e120e7a54e808607bd38376cdbe3f176132c7a41f58d10022368c7a7b84cb4a33f03cb227535a4bb273880b55ee7b520d2e82252ba3b05d9f26afe6a6eb71d0badd90b4459;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14ef574a166be74c92773329048f72fb9ce030ef707c1e74741cee3a0d7315301d7aab865a9ad09b6fe9645117ac5bbf38af5f560ebb18c3fd6d6048e9407fc84e18adae5828aef4f605a55c6ab5c0471fda0cd8a67076c897560d042cb6a76ce629aaac267e39b373d61e832a8689ce69ebceec6d7841d82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d8a80f7184bd7fbca1b0c62cf91eb920389d187f65a83570c3e65c20bc0df7d162dda4055a515f57a83afda189b84d75a05f8c0dd155d19fd8f5ffc556bc82e595daa72e69c6c3f589c1eb5e9a93c3ea841313426928fabc44c594017fd2f8ca1b5d3161a962743a45dd3eac43e513d4ebe40fb95c42a8a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18b660ed7274b9e4701b8a535c8d5ede43479902882e456f79c63df2c2f0ee836f07a246923ee109c6147e893bfb57c31209710a67f052dd61c0536adcd54a93f6eb4b617e271d4f3558aa114aba81213f02b3be7d2d91e577603180cf43a8c35e54940c702bffe1f4623aaf9916cebcd380ecd5c2987b69b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2d764bd931669e20d20754e70b0b03a3d548719564e6f2187a26672fc143ef4dc2e000b599d01c70145fef2be41afff947d453be23944319c5b73a4c3ee8292a37c1fef78d8f8c72d42a49cf3156332d44a1dc29a6e3f88bfc2047251d0ca18d86e1a9fd3ec551958b24b4ba80c44f620b9110cc3efe337;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb261de76e7e191876ead4423a942ea21a291774cd8943a7f898dcafd6995b11b733027d4da9248bcde463eb57d18c0f1624888d9af7bcccb8388f3643f26d22a0e03a49518e901a66cc1b9863db32f4f83ef7429fe3ed6be2f90f6ae24b9992a01ae0190d037b764f54be0abd738a2dfc83264f818aa8ae6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ea1919293dc633bd076aba4382d73fc06d216ae89caf2886eef05807ed052c87da54c34b3e4b4456e67ba2e5eb89a78efd9fbae61aade62c96e7cfbd23230c00d60103e3533717644929ae1a84648fd87301cd1329e31faa4bed891974f99702c58fd95218653f18fd4ad94d7cba41df5046e6a9ba799127;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15f7d7c814b4a4290b76c58a9699bb34ed131752beb0caabb55119f6399a943b83530c95142763d8532c95e9c27195d42575e947d558df84a56cc6660ff7a955f688af2cc325c162862df9501e0bc7d3cb99fc9758f30058cddd175e818efbf50b1c54c967e3bffbe29cad697f0f5e4ed5e6d9f22ce2bb2e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde91202a700a00c4bd75e0893e1f282bd76856a345d1e21e06b019e538f55e380ca85785695fcb16dc63e76da09a327b2a1498cc3c6c2dcc66c0dce9df95bc592d300192b59127a69780c919227cfc1651525810be82ea252c4ee437cb7f4d9df82ee75a58d5e56648a5a137244905e04ea87b1bbaf743ce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a76a77d0e0b45c0a6b9b37ff0f298901841d5cea593135d2e7ce34d20461808bd3e95a5fc083505952208d57f1d892a2d1f2e5019b6ad2030f8420e5b745e12b20be48d2f2b560d25dde34f36fa380bff0bda9066b47a6c2b6cb18a546078128028018c30c8bbde4fa0326ff1577f727ebf31f4323170399;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eabdd3290c4ad48d2eea75fe14031933a2de77de6407573259391e1a9137f613efbfbffedc822bfb31d782e5c794333ae2112fad56e3968ef8014459d41b928d12af0d3b75411f36f22b39037e04a86c12d6571f678ac3c7b017c39147cd0b9200b9c859f7548d539fb2cabcb3c129ac69e97efaea7f2e90;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15cb53c5271346bfe34a6e0b26c6b96225ee909a980af63e48592e512969f70997d130fa5bcc8e2112a62e3be0437b4c5f099992595aebc5a8c14910547015e065c78d1d7145e5828fdef6463673c0e73950d9e6036e898ed7d42dc662fe3abec53567165cb0471376721502ec6282b2c1d94223fa87a17f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1debea7f81d9927ff62de948acd7199c6c2c1cf4f44c9b2976cdc57d2f968236d84ddfdb6a9a430362105765c643259592f0b60e0ea6c7ebbcf55b05dbc2ee3c33b0ad6e7be1931f8566911ef26156126f044c1ea785518b1fe52e8781dea7048061c9f063ffca154cd85cdeead8cd93ef838692de15cf30c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd520f1b63d9da403c5eff4fb0ffb7c1efe1166a929b64a3c099d196e32d4bb95e63db23d4216bba7160020c8ac51027d9e08e97e551fd0e378bc715224584ee0e9ccf6b1306d6895809c3b73ecb569925ff5c95cdb25e691123eeb1612a7aa18bf8195c0df53af365544ab04eab93e8fdc274498cae80f80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3fd373f4c7c5f7096a91ab4439fb814d972a6f40f0c5d0ce1bfb2c65ebb7c0e7f5b45a8296a4aac63a07bc71ad0b870ca65b0752d64319c5e5d8989d6d3e50df208510d88bf677bbfa87be918994933a5ce41299fbc07325580c8d3819da4f313232ab768936fdfae985e7846294f366fec7d32eff4a330;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he1879e887310819cdb13cf7bbeaa568be6566f69920b67f97b18dc8b67777d75cacffaf983376f57d8fb1ea6ab4e1ff2cb7d26cfbfea0b25ca9ea71da973ae5613edcdc62f09ee43b5e1bd714dd355bc9ab1586d580f9ebc1497a8d5eee12b8aeabcff85d03426a347e3ad6dc61719ebb789d0fa573f24a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e1a07d4a5871b442380facae8b9c473c6d2f338a0a4e172bfb63dbf4d24eb3cf8bda62bedac95bf9b763d2626ad1478d8f630a2f05ecdc7588b9eb01d6c6a89c468c7b1e0de04609350b80ee17e2bfc5034808c7732e5d72c38769f2197c4e7577ef2a6d9111e2dccca89352a793d3762dfe3c87670e2d5a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aceaa3d4c635115fc1425fd9f3dee610b49ee89b36f6400bf187cdb71237279b23dd888a5b1c49527f5da401b55b3ee61e5e0899650d9f541cb3f0b62f9e3208851a554fc48cbbd87a34610149ab7cafdc17916942864ee32273c167753f60ec85c645d0d05d5657521a013062250f1c259b5ebaffe1a685;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4696bba0cd801a0398e5d8509a760921171d257c1de1a167e48e7e1bf7662efaa8a3a3e6702dd180563a2bdc3abff32788fc595dc262d801e585ba55edc5daac5fe52080b392a8212c0cb89da5b8e5a3b8e1bcebda86bb094e579967152a234452da4915c1457f6fa2ca209bbdaed2d706a7d3e0c4a7e6f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a7fdb691aaa3ad3eca0321d3260723e0e33613dde2fd4333a38ace52c557840c20f702fb61e540fc0c50139f7ba945f04454fa7f87c5a434d5d70d2a62e9ef425937e0c7ba201018f82017b5d701d5bbef989fe5060bb95f357efa7048e38876519e8531bd6b8723e260ad5880cdf176728184f836a1bdd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4667fd923bba9af6bece5a33804d474bcbdf8fcf471c0563fe6cafa93338ef3f46a4bada2428e27046e643d6eae80095b8cb816433134f0321d65837c83d1c615d049fa541ea8e27a11b3d1a4a9dc66a80c3b6f8e97a56c2b1ea352df0296ff51bdc223446fbb4e2636981fdbf0253379b1ccccb914fb73d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdce39e882c8eceac684ed6daacb3b938b915a1725f18f98487a71403f38def786cc8adb2aaabe3c50d08f6e009b52fbfe4f636706ca553d246344cf1cae97d2fa1b2112bd9f6be1dad006a63bde97b9a57f6aad5fac76510c14a794ef34438c9bdb7e140cd458aef01900ed626707e54a95391d5ff432212;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h120e2203642f0be06a64dbf24d9bfd8bede076a914e2f4d7bf1cedd4f00f80c49c77119b4f84bae8a593028c572fc75bc8d434e6b16a09a6b7c7e9aa18d07fe4995f675d5b62f505812f4fe216cfbcaa8f1d8c511588a04cb11b20f8255f08a6c9c8cdec07d324bd44bd7f588900e00f6a5e6778754b0fd39;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd077797f0a420d508ddd60deb1e2c3460e3686a0dd8246d12f250a9f1841c23cdca023a39a67300d80ac210c38d432e1f3baf349eb38f1c5247a33785a2a17940e9574dabf91f1ca16874f961a877c04688524640cc0d1d4f2080fc28ca63972256b836ee8fff51e4abf0525e9ec5ab2e130be765ffef936;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h108112a1553fd05a672a836da2eef9c342611135f895914b9d99e9969cc842cb386bbc9248557fb533fa445f626f8009a20b9df0cf44e390a989d5fdd3bbe0c27d5fbc4d48759318f0239dbb406b7801d6352a8afdac7c21ff49dd1398dcdd5fa74d7028885dfd7c061f2a1d2b9b353b4fd44f44c86441caa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbbce5e89f415713d2fa83c92c0ce4b327df1d8f9c316703e8b7d5ed586d4732a0950c164ad2c1612f684bc5d6042bd0ac3f02f0858f2965d39bed2105c3146c706fbbe55c45eeb4bb9aae0e508d82177470507c7fac941b8c410a42acd2397a19c340e4434025fe4b11c053628d4ec3c4535a7d214f79436;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h38c24a516b058e8bfe539694b0678a702d419dda0ed4cbab718598644bc28f32d15f9bcc144eb94817d835945beee38327b4476fe695180b3e2ab2c663b2564e4cd22ff7fd57503d0d1e12dc2c772d97952ad8cd26f7cfebb3b6b111ffa1b94db013e2dcaec255f973fc9d046ba58c33c073379e2b713b3c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc84070762fef13f938f4595c7e01235dca91223147001c14345eee3824abdebb036e0385a40255d385b1c50dd9c96cb30d6d6543ee7a7cc3e7d892426c275c60b060f4e39f1fd7a70106a058b837df762d08a6dc3a2f6e1954dd5aed473e6c11ee4142dc63ac43b28fa0bc0da32ad75c637c730fc329b431;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdff2a4fe32f20d6033509d3148769f03137edefbbffeb6052ad09cff1370137c88b4b90244aabce49bdcc8e803f587f62e503cc562678a6f08296fa72a132daa921774894e7e26e3ce641723a42b7d5aa280a6f283277798b6afb4177b4124a047ac926e76ecadc08c5b2336fd21b3094cb1b3ac36e7ec5a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e3a78ec028a7eccd799aef8a8f38c4b23ed1ea844adfa041b9cbf65eac9cc8692971b13f19bb36f3e0e5021caab7dd5ab61e97e01c998af7f169b67119228d2ee7f8026c14fc7d03f24e7edfb21ec196a50aed014b2ee6fba55d21d4a3b7b3636ce857108d447fcb7c238538cf24be4ba99418bfd507215;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4cf63333788a8efb614cf7c287611db49fa64e177e6e44e2cd7fbb5b66f0f5d235a97830df1cdf771a3843a080a275bf3d163c85d2bc4915ed11ff5ee3badb75e951aaa7e9f9adf5268941439567d1b251744474aa69e116cc21398eb8b39dbdf26c5488607b283787db00b749ad2ede2a3fe54dad83feef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1247defc73af42da985acf8ca2ca5036bbae1ae2d2c457001f8cb6acbea8495f42698217e77db052849d8d90600c8b7822c2b343ed44285ff2fa3e1fcd9a940d1e4d9ab484915d4e2895e536cb22af7f5687dfaaae2175d9a0457d50cf91c958c23fb7f6a58e3668ce67cb0d24fae578b7344d050bbc3fc9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12fdb5ee7204d76ed302546f1fdc564fda153061678cea089647991e02eb3509ec13522c4207e7c088338a12ae0fbcaf4b5f6f46ea7c90ba9b1c192e7d11db6b040378b1db74de6179136d13af49ecf7e0cd701c6680e41c682e33a50426b43241869e0b3a6ef0643b09114886bb6d3efd69ccd040cf765f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1010f4a3dce359e96bf1bb2bf7ab9edeeb2f09fb6e68b62f409803aadff7d4f2810cd5a62359091a9a61a2dff27595df52bea621f31c00edd27d253b2e3a5b5db62818aa2c22bb6762a43f486bd93f9ef548760d97f343c4603f8c8756e508d6cb2649ba21d13b64b92f29a78c218c81809cfdf135bc1d4dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d25ce2d39d8805f77d65c0115976fab69f1d24582f09af99363572da5453671ef8c79d4b1c9452ddae0d0ad20e1ca7b85dda6da039541266f6c303aecf68c0bc736a754be80954f4cd38e638d309f0e365aa94440d45fd291262ee47114c091cc7796044c06b9e647c069e2dbfc606340382660da4164af7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cd29a119a4ef1c8d63826fa7dd42c18a2f9754816fa06c892cde80940656fcf7da711b94ce0c1f900a0dd577169e1fd228c9c0684ba69b49880b1c685909b3ec571d754ce3cee0d1f202dae876c17c57401f2ad743ce4c04f8d4ac36d34e9787218e4390e11aaa03595c3b011d61f30ae0274a37641276b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8465fa8436671255fe6a7607bb52fa476cbd7e358344d6073b686d9a6511d93b7897e9f3241100d709c24d25b07b493cfb0d8a4e179a79afa1213c4d6a179c229e1fbdff8322a70152a1f1c7ec9f16e8b711d4481b6bced889e1dd3211cbec9a8ceaf71b380a6d94bc695adb2eada5366861e8d6c94395b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha12eba9eae0b89c4b65e2f055d8c6cc6deab0dfd7e20ee5050098a0813d27e09b7d0a008cf3948819dbb57f56a185a9dfafaa3cbc77ef0c9b85a795ed687e81b6ed7814d223be8e510e76d820b403f13a9d2842a143a1215580d939454f2298e2647e09bdfda5befe3712d4effbaae361c4d6b7b2a3afbce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h160ee942a9939b340ca1615275fa4dd51f587a7e3975fe72ea79a7433b7562b9fde3de4ee61a693f8a0e48c5eb1aa0998111f5d21a1784cd450f8173784e554775601498e50877b18f4d54e3d1320586846c4c5c2cb46ddef0ba8ede2cacddab295a8b3cf173404affa6f235135b173e34cefe7fda475bb0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda5eb0f02d853ff2f1a79f41155204c730d8d7937e0cb1835c0de7482b0a08ccf9321c3a417110c5fa78ffe81429c15b0986e91ac449423c8bfc8aca351f4ef3380af137ec7e29e0527de65610041a207f121872397679b19b4da3ab38fb462e333635037e5ac2df023c277d6b2bdcc3b7dd83b54a0bc416;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1386ed99f9584e54161edb13cb7e8e79ce03e94907e4c87058f905f054a63320f7be2f7abecbf8d298e201c460acb11fb8885634232dbec68f4c5824304f19110f4e34addbc61de3c6b285dd205e48a9327e56a5d1718f12a2600306ce53f194a91dd91b5504720e05fe3dcfe77d5aaca5fa64b9fb706493b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c33db5669d092b8cd23a5df8910c10f0102c9e33a4f9453ec53463e41a158cff365d677bb52df16ebe07b86a1b95c8c249b6548002fedcf7de9fbc7d136ed2b2f7d58e88b4c094a587c0a647eb150225e771bff21a6e1e3ed67f064c838e6d69b085791f8d0bc50c544625c6f7ddd8e20358cd33c34ab81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1694b3c3872ff79ed4a83f467294139d9ccf6401c033b3a6734072c814ad874fd2e1ed96a3ff27b685a899688b4a36e2478f8e1862a892075bd99f53fe0a05dfa15a28d50776f3557cc641a11abd5d37e59868cd19c47b959f6935493e31d27b13db1ef76980b9c9cd0a4a6efe8aaede1511248807330380;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14a00e52dc024396d52d40d75f36238cc09513aab3f0f3c548b5fe077da76bde1f0433aa018e48753ede2c77bf5cecce50404b19bd48108624964a51ffb333bac0785238fd708a44e85ed1c9cdd5962d571fa1fbb826121cf3746eb0cc18f25d18d1eb57a7854e6433d6c7eca4baeb632e474ea48a1fc2ae2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16a89310c4ef099a0bb2502d7c551d069d67a8744fb3c55f77aed7bddaada5dfd273d4927903712141513fcfd1a454521111201293d32d83a0e89685b5d183f0d5a54cb3606ef3a00819fd12ddcc0945d86a777bf8a7e6e80d8df012b40c4f20ca3c36965f313609314afd10d0286198d97ff9bcc1419d4d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h248e342a97519e48fd3c2eb28a3e59413952ce69dd218e3618bb6783eb16912630ace2f191cf1cd7b549085b732fbf076aa77b2be9ce970b1262ca0b335cb1299d10e80b73bd9cab2ccd0f54c250e96ca7f4b48687b847d3e17bebb12157856ab309fe2158a4f2c4231c87975a9fdb26f9479559250369b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf29d6cbc0992f0a33649114dc59504b0e5f4a7504159aa1e0be67a1b5749f92e96e30620484db03d482946259c88775b968b5243539140e5715e48bf74001f01bcbc4531c7e2564c697b1408ed03b571cf6a67f615e1e04fb58f0f2a47140f7782d9b0f9db561e90b6fabb0fc83f2b5eaf5c2a8c10fc425a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h148cc039193c5fc8d7582aff90ad45077cf8dcab4c2fd44c35f069d2d657800e36d22c709daf3401680c6acc5c5f6703a304241d38919363097c414c771564577941bb7af4cf291f5d6eb4573d49d53ee702779295b7de5d8f237d84f395623e9e65b83126f5f64c4148657b761cabd5414d845c996af083a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f882a151c7fc008a37e4ed18f9f8570074f7a22feb1c6a02cfda4dab7902ad840d7dfbce11540ba8504789a0dd47da1904221bfcf97a531cdd2c1549f1183f29af9fc5e55ee21973e69f72c293cc12a775e2586064ecf35d24bc4b260a0fe7d432a27d6bb9e270bdb565b9b0f907add1b162c3ca9e854cc2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16a7a8d9261a69fd6fd7509949667388415e7024c6b006aff04ad5f3d4a6a1880f27367405b5d6818b2cc8d35edd8ede62785cb8740cf828694a0ee46a9fa4112d79cfed82a27c9fb166358978bff9380ceebd953dad80d5632f6cf664a7602cb4c2a52bc4b2100017277b73a782712bc3fe485d5d488e622;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cfd6439390c9518059fac04a7298d2aea861f5119f231003503f98a38e84a79e827721ad5ca8ef52df229277af839781fe1cefaeb0408b0b6b72821f7d6855c8a0ed93676c79d554f03556cd5c0c09cc975cee49e358714b724deab03e4dde024295e34dc15960b0ae4aa170654068ff05ae436f5dc6995;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2231e398539701847949d75027d6935c2b0805991c17ccdc33b07e35518915d5dcb5ab661eb10e6fb4b75c798c7efd59cbe6165f87da0ec791f8abcf7955035b9d0b7a619308e30a114572727f66e95534d84e8b2428987355f203cbe1dd6aa1fe6d7fb5179c71450287e305063bf7d1537b2e977665f6df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147d5799852567a4094f1ee1f6641ef7c468d9c93598b7d5f9926ec5773a1e3c95ded24f1499e7e317049882ec3cf1e8d700c2ea0a71a6d3875cf824069c76665d49b1ce363e519436244d8ba8cd3f8663d0d2cff5b1eca1966ab7a5d61d6b90228c1a9064bc41649fbcb4117e20738992e6a4e0df8ce22d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15803f1ed6205c43f7685581f57c548f67582abff37f8a402201b93d411b6aeb576537641d68979f07b38964387db02e0f62c3ec100251b9481b90a4367a8f94c0b361435b8ace01713e92f47847708931077df9b26839693cd39301cc29b37c92e39ba1d1f9eff69328f07f18257583f0a00022df9184a7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b28add1918f2737945a6e5d6ff5342064fb1c35cb8a86f01705af31df115f5223a44d6460e5e4a8be97f6423b6302527499f7d7a646e652e064aed19facba8882fcaf41f3bf80e71c409dc67cc10027d85c1fa2801ada6d48be5e3d3188809b8ec528a15c63d78cb61f46bbf5179e5b3f505428fb49f911;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he63834699b397e4e0c089b263fb7d3a584bbee5dddd5ff5b22bd8f0f6663b03769b895a9befbd40abc78a94cec2c294b38340ce59182414df6fb194b131c17e9d1b03ff46ae034356561b52e115e8ae7e77b3332f143f537ec1cf32dcf953a8526b61b126515da477c02f3c8e4425c3508363cbd6381ce7a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha6d59ffe5fcfdc338278e5416e9ee12931379e25244c403f094d952bc7162c6f54f33f2ae74491e813a9e93bf82906721a095f2c7153e8e56d64b1fce4c64a02d88ecd4216527f756232ce456fbb4b1989178797dd2ba0ac5d4aa8b2a4e5b0ec8442d446210a60b3dd09fe4740c1e360b7f63b47a56da87a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d95971775290c8f1dad88c22ef13fb1dcca58cafa24f00c5fac1ef7b24406511c2acd71b6b2d19d50750ccf0138eda0056106a9bfe29afc51ebcc33854b674461144f558e0b4811b931c11c7c3afc21a468c33291ad130e3a033569c61877232b26d77329c9c34fa1cf2ba568055a28d31e4e8e766b8f465;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fbc43713ab2e695808139c72c5aa4beec562e50e48ee23122e8348607d6d7b34de4a3a61d15441b89d6132df00fbe0154e75548f3ca6884f425062bffffb936322925fb7f08192b39405b610d4b32209686f1526e36f25370d3a7109896755ac81b7be08250c3edba6a1d79c57e82bde01ca0ca0b8ba0798;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19bc4e21b9adf48ff844c762f65c9fb793867fc4cbeb08ce7f3fd4a1c19103abc2278568c625334121736d4f7bc64d3a38f5fd6b3b0783d1658ce768210a14755573edb28504c8b8d6846d1ab48e3037f5993ca32d409acde7c151ae653ce1931130381e5878c39574bbfd4e86db98c893e960cd368b269a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef9f721f717abd014cbadce23a04ba14f1cf06b137d9eb14d360329ea32a50d98cbe4e6cfca3522862244d6c9344ffc2689b2605f603d12679ea521fc86f63b20b3d055f7ef98cc42eabaa414141b2e7764d1c59273d43339620d6f7b534f457a574fe68cb0143a6cef59ddda2fafaa414238f7a17ff53a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h89abd65ae9888b7105f52aa4c143b897fbffd5c4c9f51f2e6c1773b16039ccdc2d008cea4a60344e85d6131c131b1372c133ebbd7968469b91245572e5502cc83177667c074a0812b729a333e329ae43b553187f9b7b81b1c3c55c9589563b24d3421658487201db2af07298957b440e388d4c4d9f260c7e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ddf39367111b41ac2aaf4c9621d4471dee3302b04c1e8a6430c1a787ae11102a980db5a79e09e50919eb42d13b0729178f71f072562d5d1051f658715758daf9788e782a67a728b4c3e1b8d5d8710fdaf6dce0eddd7ce935988dd3c1ea5df8355916944aa8d77e5d9d44a30c0b288628c4004cfb562ecea3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa25c48ac20c77888eb4453e13ae0a4f8af250ecb674ee291410d7e0d1618e2bf7439409e2698ddc11922803057cae0c4e7c426840c9f823a7f155ab593b51e51456c0e49215417eaf88fc9886587323ff97caf0dc85d8dc2d4dd9c7bcad19c30e5beb567afdaef9ed601880c3442fc6836e9b7b5a5c157b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf06af4c2409a25d39655dde706fa0727769d5140d6aeb505c0a1a5aaf36ac7cd01ff210a073ab6dd6cacd30b298e8ce3aa98de24400acbfe8ce3b38664d33b76b178a69ec8f52c5a0ef40b4acbe8223f8091ce483929a5ce3184fd58f9e732fd705fc2945d7ae88fa91a6d01214ed5f175365ff34ed89114;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bfc2a92dc0f0483b9d3b2c3ef7dec0aa550cce9f51d6221f36019d6bf4311e06f1c13ee2fb171692142312e46dfab30464f157d44d2cc1028c904d761f951b5872db21c2510cb936e6401f84c78e06f0411fc809df318aaecc56ac5a0ba3cf83b6cc217822a851d305f7cf96acd4c7b9d2349f087a2651bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17791c2644ac950a3617f5f26e70989e18d15688226236a7b309222bb347b313c35d072a49ee348146babc37f73e99ff0c31d04e4b53d135f08be0edbb018ebb3f3d71bdf79334f72178fa60e9b1e6ce88e151f255788a83f40211e85ab973a97111fc8d350778aee741bc28b3cf3646b31f6523850e3d7fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5004592936d93a70cbb3016358d5c8810d89b3c688d0f1c43cf82fb2f97e2168c9ccb558ef350457445d6be8220e6990a06e134dbf1220a71348704468b3b03aca4f9d586cc7e787c2cb81ac10f2d5fcbaa68606a82918b02936c2c94bf26f4cb8315074af9a40dcf128143445497147a1608d7d4373999b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b61761206428720a43e138e4cb064aa459a162a243d64ad4d180be9ff245e64a7555c8e73acf60433de21ca760bc290f46b01289f8094a65602745b43ac81715cd5b9977dae9da4f925cb21537f977a1a19553c5f1956e8d7a2cec4a689c1bd0d022c2d32d53a1f23f1c895ecaf4fa216bc2f8472367d6a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h234825e1f66792966d9d26a0b8819c6a9278273ff5cd3df4af21689a6ccf4defb8e3550c401e319f3cf003a87defce38d8d527af3c62e6bf3664fc6bc360dce60da9a07f72f30d80e474e36226fb6201300635ba6a6de2dd97017c9d119a189cfb4b51bca782ae07b5b9968ff242487a9936ac7fc5a256f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h166c10bff4da2151c55f37dda7173e966c50b3e4a35a519041d1fc0cd94fe57790dd052352c51b1cc588f96c76862869c2655dd84f5d829d2cd9ea7b3afba4ade120a01bdfca137280ece96d017e57af416ae3189a638807f2306bbb5f32802ebdd53c64fb8c5e709268703fbd536a94ff8ab4fd599822f86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1659c3ba1c69d1885f2e221f844fc7da3b73de88dde475b037263e1e7f9e900b5ec2b17558227eb44a3d3144e464db7779a6494d1dcbac025d235b5decd3283961c374dbf4ebb2dc72cfcfefa4409bad3b89777bd91653edeaba93498af9a7036e338512c23dd0dcbda4108e2eeda90b45265f226f0a68c99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17fb599752dd8412be8ff5576169568dbdf44efd185a805ad7deb259868aae172186f7a1bb7780e1365e8c1aaf5743091493eea8279347e2af5f5e76ab563d58f4466933a1e5c8de48fa289600b12ae9bc84a8bc983a5c6e3ac56a56b2d893c19445c496eca99b30a8ec4b480ce9f5d3d10ff70710ae5bc1a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ec31c3d577f0633a2046fedff891c0837783db2fc1159b39a97973f6b580447b136b11f9316a70b82f5e7241e968341cb6cf2b5fd7ceb2a8b53777bb20dacca51c6e8e367fa55518117abe094aac97ae75d27d377933a7b563da650d9574d69e30481824bc0991ff7e6001484d615627bb4a082e4d99f273;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16a367ca6b831c9092e75c906ba4e67890eb0de91ad9ce2eb764f46344b76df29f60e91bfc4f8b713d0f8b55ebfe95175df78d4b48cb6c7d8b59b95563ee6f12407d7f69e04d2fea8529fbea94bbfa1f9ba7d636b45845e5a6c7e2e1b6d640046a6e8ee00661b4d5b426a5065c9ac4c174c76345386000d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bbf1b42ede9813396fe0bcc961c942bb8085c895ec45cf4373baac1d4d2e54b150685881ec8406d8a66f6a6486c76fdff4734e592f527ce4331e3f9c24825660c4b5f92f01d6339d666855c1f91043bab1aeb0d4b2db18945c477d224a47d8e8a938c3a7017712a136498b46e17a3409703c72a70622ce1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h662f5438b8751d2c5ae7d845a50fa22523930d09500093736659d7654395f11f5636574cd8a50555ba4de35f5c2e7b810f00b30fe2a0349a1a05822d41a320931dac777b01e856c9018a93b54be7c5d76e392670f1472abf5ef8734bb3078af65458e94401695a45c838ee7f82e1278275c64d7484504432;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4b8fc29994aacce0f7d7866f8a85ac39ca7f6958d9ca8cc7870d475e0b0d5a42a9004dfcd18ed7e35c87c1316ec8b98772eb7a354b2fa5a0ba77fba73953714c366ca7a3a30f3919c7fdfabe90de9605cab9170ffc6525bc54136db2876c0daf16b912554cfd8b5cf75824ade52b3bed4dae6f9633fb502;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f9f9729a3d5e7487e13d95f82ed4f90fa217e045d3746b7fe2998491ee6f3483e961f0792470735bfa8471f73bc8ee5fab0f9489c7b9e07ea9e0c2b629046493b7055b289e769d8cdd8de2839dccb609369b8b28c4bff1ebb867db969221424bce0701f9f95ec3a28a29ef50a7bb57147fc14e450e89d97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1552d76fd5e2bbad2a00c6cfb2fe9e60860ea1e0322a440d0765c59f17229bca1ff7fa8e4866f2dcebd7da7d8abfdb4f3f845ce369611bb066500b854898e47d1ad369493653e3d35fca30dd279a2fc5d791e36cafe17a7e5112f0d5556297f6ec5c013e1895aa6360034bbb69d42af021eb849f951f5f483;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186b7e76719708f185837506dba0b64a4feefb7f23f9c9b77972a7e86b80b2f73cb16050abb24091431e9658dd22726b54743578866b3c78205157f63ca2086a0d2759aa135946354a40db61206c4f0bea5ef57c37225ccb58dea10e6949fee73159e5148f534dc76165cca21b15b2fa55479ec658e8b4a80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f8b04297cc0c19b445ae65903e95afe629212aff361afcc0fb312136460283fe3bd414a6e6250db8313d33689b655a3572ac89b39fa2190f59f6641dc9193d021ad80fb3f0cc035bb1ff24122552b43a51ecb1ae3055e564c216942b6a7aabe34e81a65669f5cd87e72953ee2104aac6076acc5346f7141;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d490cf06170a1f6555cb056318321db2d3b525e0d8b7ccaa9a7758f3c66e0e3b93312ec8931bb662aaebbb47a85152ba001e038d6d0837d762f8bd5b2679f2fa8250200cad1648190790df16acfb6b91f015f36d9943d29e8e9332f01ab2b41a774a1dec779a850373aee9584c343dcc4bf26dd72397fa35;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h140b861b640a0baa868827e2707dda82c76ed6d3a9e3636f5e392f99e4834459e7858eac54d923d7611a9a571e9b75b08c2a3db1bc2ee4b032b0fff96d567d24e4449668e4ef37cf7bc4301a1e03a234fca525704a3d39990aebf9180289da0fe241c3b8a3af226fb42d2184ea002676dab86e4b6451b0561;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b2b2ea1a7bbcccfa60b64b7070d8170c582616c99cc2e4b94125a98deaf693078ef746117ad02f20bfd60ae3d2c3698db432a86d92fe05d033035a1ab0a208432daf47053c55e1495d23c68af75ee55d6f841247b7696ff685cc45b5420af9788d6ade49c8bd796989dc7346a338bb3fb3a995476edd1e85;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc29eb787b7243f2db366e0d766a8f5bcde5c504762e7df57a925acf53cc95c7eef3d2b988079f9c1e0bde1008e1d7b9113d621ca31784f8d47112142d58a25511cc342ff566f9b7147cb3b8f8073766f1682e236326b99c9088c4f1ae81c613fa237ee0dfa409d7544561e630aa69ac3dbc18a6c06e0ee2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d77392a33ca744b0e6f6b77819c3ad0cfcfbe9e7c94300493e8d14621a17ccddb556af57b7b60282cfa80d4fa977c015fead09a50b386adc91140f84515eb3584a14140081f32c09dfc0eb5d57616b7681f0c72a1018b7761fe2d1c7a9d9e5a763bc7618a54d17791b481c841546612864d65d3c9c39b8e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf01dbc059647b3dd915617e7b3e8fb39509a43d7fd002156430b5d83894f830d6272c2a25297ba201327ad46d181276fcc570237832679fa9f3f71f7761682bd7815e1dcb467ab41a92988f06fc0101af4e9191eac3e3e3b80705689d04599b539e484c8909eeb60ba9a28ffc2c23e8e3564a9482325c9de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8bccc20ec4b2ef5d144762f272e45cea50ca3104af1bd87ef373aefbb398cd523951ec565a0e6b2c4b18f8cf5d9ac336c93831f5c0af09b0b94f1e92c619e2d8ce740b04e002df08c1e9a8cacd48f42ec13b9b014ee5a4b3c9c136c2b309bd272c698c1d436fe4fd63d14ba34f81f85a0710f7f24f6021f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d0333f96bd1a4b38045172b0664eaaab76cb56be5726bcbec8ec5746387e8e722769db57aafafbe8feca928c3796ca118063341d8328dead1fdb718a7d634f062cb05af46d8a3fba240839fb96ecc184a9a5689398d590be570011456e21256ae01ee3f9e4fb7a3fe51527cd2310409ccdf964d944c41bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d0ad5fdf66001cb040b285c8bce953ad5c44ed5b9551630dd22aeb22c9248ff2df467c1de8bed9ba8bbe1cb709b1c9815ccf8f673099b090db7876187a49e1a207987545b71d8adbc528a7cf0eae96b6ad76954412877749a3de26f6735535c888cd9f62ee8cf8875f4e29b285b2539ff96db1311ab2cf6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2476159ca272347f771933ad30db33d15c9b8763714a06d965b1fc37eca31c6de51fc29eda744a6dcf9d2cdab6f0382de307a5fc434963c74195d40a692e9c18e3ec2d9c2ab74abbdc628ebf05214a223a59152e9504a0d1533277d3d5e476c929f857a17764a68aa51803a79e06da3cb22384c41756880e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13d599c8587c8d48f7b75a667cd3ea33bf5492422d573ac2525c377474f891dd12a771633dbea93e358068e90aaabfe7ae5f16fda471c5a3ceea5a7f6f35f63390ada48a6fa47933e2c3f18272228466d384a07e507faa202454c996cba1673b6eb257922b3b989c0347a8f06df30b564333d26648e135915;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he1ea420ea376712b81fb99c6effc3b326d1c65d717c77247962d83ccb9890edc5f5e83a3bd30cae5862931ce1f692db1b806e3349570f36b3cbfa6db56cba3b23a8f55eafd92ffa3d452adb6da89dada88b6d4eaeee5a52b73a7c8aed23bebf59afc57f864655243f6f264a9d78abbff8694c6bdc8c2c590;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1162cb1f69c5a5b06c4015ad95144d094fa955904360263d327c85843cc5600d4235992ec452148f82f0480eb5a36ddce6dcab7dd4a2c3b3d4f2b454e5ccdf0c1f866b8d81414e9eb2f4a2f5dc1168e17583a835605becc35b3531d233de67dfb871bdde98f48b214b8720f9263ef068cbb5f824896e4852b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47b540f8e7478b85b4b50119ae3c638aa08d7ad2e3241ee796404ac92098971d18d753ad84dbca4312e1843e113a2f96d9e1d15db2ebe84de9d44100f318e046676c0151c9d1dbdc83e83d98f79e33be359066c3fb8132037b9a2cd0c8d671a3ee55fb17e5c4a63b7803bc50be4bca9188773101453d44a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1965d8e2d81cf1c42cddbe7397be93f863ead293e35a0e3d001f2ba2d191e88c18e8ec655bc824e7dffe38a5a6acaa377ae3a4bdca5294797a892b55f22669f528ce7a00151f451af24f6262cba6fdbad2e7872ce0ff4ef923500337c504615320ec33aeac4c02b9c0faa495c8c09d9da6b75108e69568b22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1162cd407a19f199ee4979b4e919dc27e0897736ece85b7991b87313b20f627d09d4e22ecac1e8a5981e440f92908e31aa4525e97cb8d052ef6309c49c97fda59e48822b69a89c959d30f6337df9c4e9540c92e6df3b2ef6d82e81d3312fb6e0d994b0c0d81dbf0ec8ff722269b813bcf5d4cb993d85db88e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a62e2ec83ee102858408a012123ae284af7fa5887c88b85bfb7df6d93cdf6b9067bd42a9a653c566440e7f056819d191641ac9f9599abc832369af0274a80b36aeaaf757064f2a9897e679c59af4e286e0d2cc2e8763e398fd7ca17f0233cbc6a3d7ae328fea06ce725e681d1f38cf4beab85ef2de084e0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9da5c9815c359105cb92fc928ec182c230923d140deac28e83b21cf83168923f6ee1dd792ea2fbb42c53b4f2482a2df19a0e28beb5507a65055d6f2509ba3f85b0e1caf66a1b2f07bed4a7de3af86467d93b589d9ebac0ebbaffeefae2d2334a1ebdc61f8ba7397498224cb6051b21d09915e092d394603;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e29904e218e5d0256faa07f65ad64c69d82a000ceac3728c4f4c462fa2dc0ba9985a4fe98021211acdb57a724b5bafddc2c47dd3d1fd3a128fdd08441950c3b5498b02e95a8077902b2ade3ef91285b4577f69ef610347d11161eaed07e3c3bf0678438a75079dacb00ed2cdf68ebc8f1e485875acfee59;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f6e105d397fab2d13a91560badf0b990c4855a5d16f5eff8af6144d3d3722d9c0cac134f4388a56d51613c7eaa6e2e3bdf2c0dfd9c82e764f4878eb9fae43f0eeadcb48c6324d99222b812ff13d565263f754611d9d4642b578f54537d96c1f538d844a7deb3239e34fa5fc70ab242a95cec8e5e1850f070;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4dcf0cea487db6efd01875b66d8fff3bffa652d6ec32891aba1006efcaf3cad185301b201ad1632c539ef9b9103d6bbb6c989ddb7e42dc6f7fff2d1dd532f9fbcbc2e4e62750903b7bb8a2462ababf858a88b31aee294cbcd6529b3ab249ca831caf66526f9ccc10d8dbb27dc6ab44a812e0512ab4d7eb0f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193df35c4cdc39536b8e8e3b7f1a12c8ede88cb0a5d950bf64e5d209a1f8eaddeeca17a2955aa4793b5f371f5b994f9474ac1b5f007b9f843beaf4d02fac99af1f5b2f959e15b975125026e6d7b8779ae8cc1abc77cf9703192fd32bffd42d8f2bf61bbc864e4f94395a47699f4cdc8a7d4df4cb0108635b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde6f64ae71d19f84b7f668ca49ca60f20e0c6e498a29ee0f24754fd73b2ecf4b6b5e19b74056e9c1526bd0d36f892b7ac2c2387874129b840d906cfc8b684f4c5c26651bdcffb88f58ffba049b01fd317c5acce2e7512c152490a964e588d9fcf2efc87b04243a75a4bb871ce315a895484ecd6a6217c749;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9621c9c152c60b59af2ac7a7aa7add708da1f86632718f581f54b37a6831427547c1731dbf7945d777a012fff114c7e11ad5494c1d5b04220ec038828fdf865db11741c9c93818e8d15793b084f5d9f3a18ea25c421ed2203ce2ab74729335e64ad70d56e0fc88d3d24d23c0f66b2e4a3052ba453b448bb0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h182440d045e8cb45530be775aeb6b27e34f9c1b3bd0889449ec54248086223cec9f82ed6a116241e85961a04082a237675645634054dddf446b1ca2cb6d20039fb80dda240bd785c645954718f168a8656551a81b86a1f4f231b7fbf2b78fb4812faf924321bd76324c5bd6d6cae30dd7bf47658bc48b3146;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcf3112f399eae902a67a74b66ba33953e1bea486b1b1641ac8088ae64d3c3fee86be0e7f947143c104f056d44978abd35c4b0c1eb79c6748bc606830503cdc89b70706ac2b6e992a474360f6ab108e8a4abe70640bfdb3f808ad6b0d38edfe5a775b2ef3a1ff0de9a1abe0855e11a0124bd6a35d29a914c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h36cba66f3c13b3af134cde0225ee7aa11f1c3c565112ee5c4cfabe3155433c36af4d04b1ab910bf6674b591955457ba9813120e936d0f3a3f79561df2a89424529ddd9c3ac4983a1fe59ceba9d2f02bb106d14c07a67279ceb6ca091cb2149e6f5cfbb0e980cd5c1bcab0499971ce98fbf178172082c490a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1588c2fbd84dbed90a77cd57548ee79f3722e076d6eb444c09caf19e3fe483774e6fab2efbddc354e160ee77986814fc52cfac5c19a5f2791b99e6a00ca53681261a332d418c6bfc8ad056146f07673ece73ee986d95dc50ffef8239d0d9f6b8739e6334d57578a7ffc174888e54ebd21137513b98bf4f32f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118c60d41c71bfd9bd743c099a77c54252d790e5f819be016a0c2e3409160e9e39dc7803369aa36fd79ff85668fc9d2ccb9da87607c4d2e06e7fa1bbdbc201bc7a84ccf79b51e96502ed0f9c674079bd5c7efe842bcaed273428abe2d926cdbb5d2a30e63d98221f6e3674245f4b69f0d9b51d56715b8ec7e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1581f5e427d1983b14a06a9636b592dc8532fd2764841bcfd107eb7c473a5f41b8b90e2d61301554717d41b940ca5e244478c671bcf9d5f9953871bd866dc710230036292ca08cf00b2d746c0a9c903a66de5ae27b919431d1860e536a1220200aa9a57b75c6c65be39c75844c82620e1d4c9ad73a95a67e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c8756002e61688dd3854a78afca43decd4b00be94533eab3cd328395337f376097d03742da635a2a22a30d7910f22903bc47c8aa900c949f6f62ddc696c1ffdc37432976438c0808d7bb69818facf72d2244e111f2157cfdeb2eeadfd361a614ca0fa216c4b3cdbe112095c2b356882e4cddde6f7ad7f59;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f38692a418849bacc6604bccc662a1133734c0beed9d1f63765bd45c8205d2d8197127c17f4016687d20dfa44516fb967b4a1a503bd679227b36730cd67434d4d169d1db276d1f5675450239c4106adcb9ad4828e414415776c42aa19d00130a85499c323013dab29ed55a6f4308c701193c32f073e38d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1bab237efad8cb08542ba0db6178f756372ef164e90ab92467f2856578b7c913cbf9458a3434f2913e16b485440bb8404ce29be25a3cbcf64dd5d6d54942d27bb6e30b6b61e9b5d3846f24b43d0b9c45ae6ad1eb47bdee0df516e854050e26eb4489af28538fc1d343ccc84f723f573f72d7e2d549f9244;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb4a2c09623ff56f02a6062ce434e8451f74bf40e4a2727313affaf1dc8830505fc5c838991b74113d3450488ba1fcd57abb8155d9d3b768aa139c2b4d6e71046652ff6015ea28f231f5e44f189b81bd39d4c4830c40afb6307df1b5f15d213b8c8b714c89bd370ec466abceac670ace1bd20f95cd3329f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117815a710afe35e731596bdb85855d78fb2efa440c2398fc4c296deeb02fc9989fac459e3ec86693a86160bec7b7ea217eb99fc99f3acaacb34eb7d1007b84cf8c3a76c31bb21f1dbd9ada714bda2c427ceff0a80db8b64bc34324eee775c490214e04c39a30c6869294923dc151142a2c04c5af6097781c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h89f98ab4131f2098c3f60c93644bc0fc6791e59cde42b692263153985b9223db3c2da393e1b8614076191e6b42baa3272e81367db2db594602c6b5efa23d6bbd45a85b56bea21778f8894029f29e6d7a5b6eb58cb0c0a6d20de5520f85c175c16f91f402e8eb7325294d025f21566eac1c008febc2ffb201;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb86635823ea0406bf41f38f355b0389bf3bed0c8c2640548350bcdc2bd75d8705de404a818c85dee5105fe954c73fcd662048b12a02029d6584b0a9de5514f08442c290931e914612fbf7289f330bbdcf8e87b7818caebc76db0f217cb20deb140f74b2f9d36a50cfa97bc2883ee52080ee1acd985603628;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37777e8d5f9012549b170e3618687a202cd90e23874505632a4432411e8614e9502c32d8e67596793fab96996ba1c2225de1a4ad6d125d0df9ac8d7430445e49acb505089d4cb3b25a0fcafbc0b3258acf0a3ea500d4a954b9ffe52634b5ece2f0097ae38430e8e4a30b0a19077143c58eb3e832232c300a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b7f20f215b7f348a4e66975147b2314539b787047370ebef04eacb5e60dccb013d55ad3a95690578727e28ba22788cb479f12fd7a1bb5ecea92a45332fb2b260f788c7d80be683a68e1248e9b84bf4d40b44929351859aab82f4b99555083b496638127dbe76d8f056a418e7e2e9f37c2a1ea2c5a14b7c99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192aeb22aa13bf7fa248de23e035d205e0d9f873c2e83c0cdef02252e9882775162cdffd4d09389b5009c2c66f88c42206f251a8de2684b6b8b4d097a157421d5db002dbb499694d07b770035c4dfb41a4867673c0544c96a33ffd9dc3c7b868eb92e6789c1c6785b80879c910ca99badac61c2c580ebb891;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15d4741263b664dda77175f14bc22ae1774c891939383670bec86e8f9176cffa5fee6460bf9bd401bab9bf359115bf45af37928c9c5ae6486a6ab7894558cc4d11dc5c99a4511a56ff4e8e885ca1069e0cb7a0158d685e051bd115294fc6fcbfc120eb04fdfd0ebc75e1a0c7d2223d47a78cb04505d38a6d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19cb306425e907e17a4495e983c44108920b9ca7bb8b53eb00dec2fca69d73a4a4248a7631e3d7a1a1c335592c660b86359a14d6ddd2f4be42c02d8e52bde5ac0418df47ca6a4ca497206182b5aa15d9bd49e7431e124f854a462f4e60ade759826c869cf992d5b83ad2270c8af8531b1028619c9132c853;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he7ec37bc8f0d19c9c7907e09d4cd4ac201429952f1d83846fb10d623ac92c340ce018faee5b13dc10a31f22121f180fcf08efcdd3a7c102c80795eb4efbb42f6bc0a2efa5110f6c119c5320aa6359282641746364db3689f6625b10544ae75dc1411918643c4284f8d879be12b921c213693487de8241458;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h130e5e890144f15e99bbff2e7225eafbc63ecf6d8616a21bda66b3d9d9e93aae1a1836a7615b65bf41c4df018f06ed99be8de2cb4fb020ecbc051899f35b46a3d78d43068c617f43bdf85710941c3ad2dc5cc8316c8dcb0724a21dbd1b98099f1fc114a23947b932668ae89d68d761d0fe6dc64cde0fb9337;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb6f4acb892c1622f543ff32bccafc44fd8bcc169bb381cdd262d84a1d0f9cd74f4ae6c9496c847916e3738ff7af89fe3970dc082753cc6a7c379fc1ddd29e2253982dc3054cb32499866c249e43360fc8ab715e8d4d50a1ed8bdc1f1aa8dd9133c5204406d08cdcb603d286683d0b1580912da0419f945f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb1dc221fc781b57c5a52d1e44d6de83aa5497c8a07e936768f63c5939e7c3682117cb600cb26c96b77c396ac0dc0e10aa44606376bd8ac6c02a9b53b0482f243ef41a7dae09e3314775b7c9759d8ff308d19263a00ef08cd359781ed20a661354248f956cb598e89293787be797b364f27c81d236f6a696;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfe39f712e380bb0522364ca13ce1dd2fd87a80cdd91bff25e68002addf51dbc0c66da2e3ebf194f57017aba54d160b52fcba5e6af81db9cf235526f31e1955955141b448ea2a385c1963c7fe901d07f7c857744aa5f73c9b9c1333f6420abbff461c4daa7a6bab8506ab129bf9f3e139e7d3f6ad3baa4f15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h43bdb115f87612aeb529861dac323515406a11c0ca193b6e071d5d9552e9ced3b6bfce202063bbb5445573ab9d5d6e890444f4a82a98b04a7f4fa99884618c6b1bd84d2c8165f28d5d87f70b32e5ba182dd9f9c0fe78816e9e5c3a24ed642c1f5f84787289a612d241b7b5802a6877d2fb6c769a2134ce47;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h588415ebf8e2a33dad806875a271f5039b363ba3ed6518d39f3d5ee8af8fbe14fc614f4055cb65b398b9f7d5afe7838d324008b1e84e9b0c90c2f07ff72a842ad526308d9fecbd2b4eaf920c1d289d57e669cb05beb49d7c0fbbbd391b0e1610e981872c1d46236284ba01785ce8729c7610f7ab8b35da55;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa349db86b0fc8364d80d0ab079a4cae7cd204a9b2bcb9b340cc8e3084323c04c7506eb81c33a4b62c057f9c43cd48d0ec6b1f5af7dc7731b6f670f2307525e0ff5cd184113c1e764b71e71eb7cba689d8e7a2a6e17b29940cd23dc4ba244775c3c43babfe696e015e45ba4e1adfb2be21b5b22397a9836c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf393c896f04c28b9226566715cfbd7b10c5ff41f6dcf44b963b81de5d5cbcd940e4e62b7b976f8ea5e2b1788b6d66a58045387573bb386fa78782c98743fe909326b60897edff26afaddfdec19513c067cbe040b1ee9c16ed5632b91652d625e57a57d378bd2856b165dc391ead6432ecacc4f7b642d6dc6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1086eadafba778a7eaf665dc4f3d3c70e48d9cd4292c29e54fd22d288cc8c02a7e3a866907b1238686cbd1b69c3e46ee3715135605b271960fd1256068fe1da11fdda25edd9a664c456432d2c8bfa679588e43e81cdf853e883e20647bd2bb153b47ea383472e3d7e53b4c07929f5973ff95fcba7c07448a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15fc2360d5489f3461471f808c81e5bbd9a0392704c282ffa0370726b9469cb9cf12c91a3f6c108666a0f9baa1c3c50c1beae406cceb6dccbf8e6a4e9a8f8fc5b22368920d5a4288c88c98bac709b2e561176a935a4b436f82e6fb0b85855393636edc15ba7c5bd9a5f880384df2443a2ce36a2e407ad60be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1562bcaf7068aea5e11c60c01b932a1efb74819a38cf0303d20ce13ce43be74e109c17bab62a7700af9f21a6c1c6a5babbc27d31fa0b1af77e4f45d2dd1aa27c2ff1082a0bc36e6ad04f4d9b60e127daf8710a18095f646b1d9a3a7f774c02ace161d2aab631749859d8bb1e69094a669e0dd8f93fcafb53;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h717b4073f7932562d87749d0e0f57ba947080827367bab7dd55d686a5c02d9495c6508cb1254b71ed6239772609712b4d0f64ed4f78d9e2e88a3808a79cf813b87a7923aa5a19773d48e36e10861dd6ca4297f0d154ffaf2046f82dfe3cad275393ce49fca23e8cdbc34a52a3265e57bd749c799cdcc59e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc7d88b8a9b3ffb99adf8018a8d5267f19e1c0ab5aee45957d3c44b1933ea8a5acf7e8881fb83d258ddb07788eed6b86587a9fd6189b7fa698fb4b51b38b0d47a714176912ef31fa53169ed51989bd79f2bce36188d92028dc4f75912a57454ac579f92556d255e8e60365f80d300e7f5bfcbd8dab494ae3c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15e5cf96643189ae5802edef0133a2099dcb07675ed85b4713a56c3f59c16d3178d7014ecac3f0968cf7f2c71a06640c0b7adfa7760359ffaf299d8a0e919640dec76d78fcc5d844c5875f8567f546c5ac0f7416258c9fddf98a5a44b3eb093a3112b68f6b137ff23bb6f989763074e2ea89cebfc37ff14ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ef945d7ebc671341ef859e507d0ed0f2d3fac6bd1f6d946a517d5adc3b26cbd55f092c4bc1aa9c67e923edb4bc0e268e9786c8b258a841ea321019e9a95c53b3e4078ffb906138b16abc0560df99641a958d4035179b4f74b6c8cca334f19be07ca72c596897bb0133ced0d3996771b1ecf9ac8a578546d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1080838d85bfa35b43e1acaa2873da6ce49500b293ebf02fcb327c667bb76df75b3f960cc003bb6441f5fdb69c9ecd19c1f62737027f88a5af5fd7d6e8dde750e98c51369494a2f3b0fad2ebaa7fc59dbc5ffde9db8343d8fa14e0146fbd5cabf3b213455dd5353e3b785e80a4b241256ded3f21e9a074bce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hafa8bb10b2f2ec6e463a65c8e5e1577059d1954af68cb8433fd2f8850b76de8dfc413a1fb74458bb0f8c87a76ff3e5c338806cf9b10067d99fe3c5f677930500c0e035b6daaba96a8b1958849b512421784e9f0f64da092ea668cf48833f92301113abc4a754979aea7b7c286847d5a7375a68e5336443bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bda93adbdfc8a9a71ce25bc189911814249030c88ab46de84fb1d751d4d3887f89ee48785328721489f1c8eba134b027ac824eb2592b44a7093ad2d70383cb9f0eda63dd9fddcf5289be697ec163d24ff05e807f76e172a6d3ab7d8fb2eee58a5ba74ab33263d66c9faa03dc0e3f279c2ef3e81108f176b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h773962553e6f32a35fc14f868348f0025049ec515c76b72c6c19abcb4df5ce562da736cb31974459a6edbb3d0ab3be3814289148441408b1e3440cac7a5ac1c22d222cef9517400876725a10b3bf8e1c68c339ee29b5af218eba305081bca7809f66752f7aeb6d344251dbb79319a2bfecc9a6eb03fd6e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5c7464b7e85ce729642d7f1027b70bea4fb6b3c255e7df2c33a56d7efa01662b955beff2b7430c291f901085a6e80d45c24e39678a494f71a899abb93d1ffe9bf47a99e50ff8f6cd3faa26a83e61347e6ec66e6c7dc0f3db65039230dc193d4e53f76e713029799be65b4d87b36e9c24561abb33f70d5d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h154ce5559d0625758c6639e92d47840ec9c02ddf0fde0b889552d78e582807d6579029a3d18a548d73159ca0dbfd308c3dcca784a8b6b1f803a3f15511971d525f03f2a01d6995ffe1e5e8f6d68aa146d609429c870c99078666ae58b9efc5d4d4774dec7d936c307896600e0bc362e3d08af864db0db0dc4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ae6083f99d9c0f389759c69e02c1e976fe9ff2b9104785814b758d8de833b7c0a19df72969a7e808db370eb97f3b7ad2fd077a9f20d4f34849ddfd6cfb05f695322bda49aec7698094a213e7674b08c83a3b17dd34325fa61663aa902e0905fa7418863ae390f51e3b7bccdc482a90f0afcc2bd3cc9d45a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1766c4edefb2f732a102f905d3b537f40615ec3a95de9e33e4607638ec82a748b7453640d450942a8bea9f743eedb35b785bd98cd9ed5f123b2f2bece1b1c17c78fb874c4d5a3e4e3b9a4b8388cfc2c5a5313bda69223e093be9ba98e2ac398076080db40e3e601bbeed3b426adfd838cf0a6879c68ab6ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc2b6b83069d70e97e87718674710f4a245587a2e162eb676e09a3e56d9a370f3bc349d4381863834ac5ed0340ca76dda9d9b755778ebd441c78b3c337a97c69d47ce37475c4b15d856d8ed4ecc9b6a8eb00714d65bf5a3bba39775ceeea50b46de5f4e199e809d2822ad2a0030be2f1d1c9b1a3e34f135ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a6768f632a1719fd27bbbc2a7efa5a1c5825d569c0c74839feb9bab1d04e1b7a5dd08eaf1c77826e628504b3506a9870066f16faadc74ad1bd8600d5125cfae6b87c4dcf2da481da058c36cd72df3cc93161e23a53a5622cfb203c035f4b0ab35c7f8fe3e49c2c464bf8b1795d9d94326fd7b06821626411;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf59de7e2f39ac9060e1ebf2891f0f2d1f45c0ed44e580a95182215ad1ce5db27c50347bcf302d371c8d98618959a5440edd2b025a6c8f5d783b89f24a2a3bec3d79a463aa3c456e902646c8b3ae0fd7c224f7b5e3f47c746b7758700962c3550deca6ad5d5c82a25577812778848afe439725bfa2a8189a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb59b6462de110913975f1aefd9f1e2a707fa0191e76c05536c30a35a1d75c16b22bdf929293aa51958b0f6eabcf1d9b4848d6793ebc3e50671b020a0eafa28247057555031c95f52ab88642183705784ef316c12178ced300fcd57d0d9161841356cbcc183a95f86adb018c050c9f9b574ed1ab3efe68ebf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2288c6c2e4dd442ef9407043ed63e7087b693eec527806568d02b5c8abd3e77c2dfafda4e2b946ed66c5d9eb2da524e7266b4b96449aab4b6196c18e3147175ee8ef57a1f439b22b9a94a6cf9ddf3e90c26214afc5174b4606595e4ccae33b78fad451caa61bf042a3c484af2ce18f2eb35142378b316952;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12abcbff627614765e56ccc99f7536ab2104e16c9617269b836e4c2806e089185446f5b4ab9462462a4209a745289a2ca84ce7a05fd8d1f059b35cd690aef5becc915a953a175129a595e67c9e2754691dfb458020539f06d62694bfdf7364c7c59e588f1dc525df41404bf5e3d61cbd8e183555f9fdb612f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a042140258ecc8a59015abcf5b0c46904468eb302f181dc325ef48811e9bf59fccd8c98ea0093ffff429c156f4bc5701fb9b186e8bbccd5bb529f9f4c12f197162bd1a7a5954968921336501ae99e84a1eae485b4e6beec31e37e37bc6d59a4b34a9fa88cc5a53a3e0ea334757e7c1717342f750d5d22bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bdc50e614de465293ffb76637c9b4aa16be57764a831f415a5fc63e4c7fb5c6d7bee5da7040b88d2a18731fd316f36d042e47c3129c7dc136c09076c3a62cdb54d465dc4f79d41ad9bef77f5dd85592b07cb56bb6509251e15e25f879f427ecb2a7396017f804211e1906ec5dfa86988c9f7d488cadfe47a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h67b6df00985c06659fc5cd7de08ba6d0792a6316cde9b6d4de4c18498d97faec3a68d47a8c607a89fd2bf05554b3d89fe0ad68bca3e9c9f1465dd15b991dce5ae1f32279d03c7e704e7c53b1d12cc92d34605bb8ea38ed48e9906a6a79dd355c0cde13648a054297b2241c1848e857bd16646b2e039fe529;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34763fb271d54f42bd7e4769570edc99432cab28a219a30c011a77b9f1cf802167d5360bb95b100d0fc7580c41fd2bc281884fc8f7105a85cbae1f937a7dd65b25779b282ddb09f6edfb83e16ade0a2f549ce9dda257235ab0d49498943ff0664223b494d212a4e3ab68c63aced89b5bf0a3b9063c4641bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d4812d287594bacceb3a0bc78da1206d24986da517796fb883c267d9ed8fc7649a528060db1c15076c99ffa95288c315047a2d7a394cf31b453e390494286e49c6eb9ed317304d2d4c207f990e42c93c7b7db5fa0fef72abbb3c97f7e10bfabf8edd1684427f2cc06b6843e31272e52acbb0cb3806fdf012;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1688ba7ad185f92c47f4da4d85c79fec870f60d699d89f45b6a3229571f080544d3248951d6b22f53280e91285c5c55beb171413c8c77dec9a7750e924fcbe52ad56aa74541d11723aa5b6f29fb6dbe4f56d69867ba89cc78bb95a92e6aef357d9defd82aa146c58323455e522dbf46720c34b938449338cd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h97c9df16ccf61d35c416d2014957a1ee0dab5912f24a72c17edc5bef4a9e7790228901bb210821980fdd74e5f2821999d3336e7066958d1098d3f47759e7e2195d5d58769091c3cc0c425c7213a75a681e5b10881f48618fb2d2f9e9cc058903515d21d58672c44d112f7e74e3ef932057ab310120df6211;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d65e72fe1933bd65697ba73f8c3f27114b983f3701d8cee6d4880959347a8ae576389d42fe1098f0fca1ee113b16916105c5e382a6969fb92e195df74d8b5704bbede7fd80a84ddfc63f232aeb8ad567c8dbb2d4b8f99fae9accdc64c0731cc4b126eb20fb844c8b8c5e0c1474c97a9c34f7a45f5178baed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c977de1ad7e562ab2bd37d8b7725aebc0b311e74ee8711be7bde3e347c0d1327a562ba81c68f8b184891703c815450b7fb716b3ea02a312bac85a0993b381342a6553c6cc20d5ae77004623f470f25c02f42c41adc588c8165889bbe8885bcd26d861e810bdc06779289a6751830d72461d9c5fa8b51d0e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18a400a31aee9282649a5bc9e78a9222e48f311a6a96d49dcaa06197d7b997073af2321cb5b41c9edf03040a31c1b7c06a2c61fd8aa10e9487f729ca6087d45b1950ca15f37e3d1d649e189ed3acec65504a1496322b6072c849e7439c7e3fa2fce534847847f8ec5098309e6e273d2ee91f6ff185105bfd6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4762085aa704b3b227b6a138589738f8e5b8cec28af509463261399e49614ec0fde8c17350d3134d190b71a09a2e84e986d3b97795d05f582a4f924f3b7f0150e901c3992a2453035d800a3511df2e302260d0225dea8caa6df5d5a60982a494655fdd45b9f73709f1bcf57ae4bf5bae051dd6abca698fd3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ccf10dcce9ff850fc1941c33ad2e8a81ad62f0026292eb438ca3ae27c7639e6c5e255018f9393f9d5f28008b730edce571616ba3890a859c5046f123a43885bcd999ce0c4c6dbad212e8676115dac1bc217ef81839fc89fd5b435a3af430eee8d6c11e26fcf8f535b14f9d0fcf368c2be9e19287b0db9e2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d62dbc900f99808a7f4f817da7aa11467686641050cda85819cea362a771aa76a159cbed81c0d77e88c6cb031e80fec9db10bcce7899a2dfb985506d1c653fd79386d4dab65d275bebcdb918db5ff45cf9a82e9fc3e0bc9fb752310c9d83b9114626f76f006116ba86b9c051bcd4dca88858f44d0c67b961;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1357e6523ee519eba7efa5ee9f4bbedf1f513f1ad0926d607ba5271a3a30f22b4ad627f0e0d9bc91c8e68e84e198b7fdeb3b04b79f91fbf6ca99f1b41169060c7b3089d48a4baed3986de06d972d8b5e3b89126f378aa9b14b9cac915e915a29eb4e0339978fa5106df994af020ae600edc99edd99ef82858;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfd7488a9c336d1bc0fa4f4e6fda1df6d90bff400fe2c3a75587dd187ed57adc887db831d663a7142f5215cdbad66a9e056b08ef49714a325157b477cd47396db4ade6cdfd90bce3979ff73e7ccd0ea608c34ad7b24f1ed5825e7f836011f2762715e134d1303e27fe52713a2db1937683689e0e2125162da;
        #1
        $finish();
    end
endmodule
