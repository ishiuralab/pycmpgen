module testbench();
    reg [22:0] src0;
    reg [22:0] src1;
    reg [22:0] src2;
    reg [22:0] src3;
    reg [22:0] src4;
    reg [22:0] src5;
    reg [22:0] src6;
    reg [22:0] src7;
    reg [22:0] src8;
    reg [22:0] src9;
    reg [22:0] src10;
    reg [22:0] src11;
    reg [22:0] src12;
    reg [22:0] src13;
    reg [22:0] src14;
    reg [22:0] src15;
    reg [22:0] src16;
    reg [22:0] src17;
    reg [22:0] src18;
    reg [22:0] src19;
    reg [22:0] src20;
    reg [22:0] src21;
    reg [22:0] src22;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [27:0] srcsum;
    wire [27:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a7e28f3d4ebc1f5ca644f689ba7dd246a33967d8858c263849046f0031fd244625d693f7c0559428388814db309de9ed3662e7d65d9a5e689dfe05a871be7890dc14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h44d7af1b1305c246a7d7b63a07e219b64f1aeaeb0307191260f7014e93ce6b3be7a3261a3a307343906a08aba3d5957a71b4b0c2884abe368f73f0ab89dbad827d13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0b4ed1930f5e698696307db208c65447ca33adbf290c2620db880c49ce8b0ddc85deffb7162e167ff8d2be2e71ae12093029595cb1721de3fe67b5e20a684479b31;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b1857dc66bda76ae9f1704260a765a79b8715a6b25c1e40b1497f9f77ed2b32afd4d607e32e832c75e3738768f7e27c41afe90697a0156234c289fb8cf5cf1bd1dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2f72987a4b92abe99febb2d3d54a29ee78a74a0aa9084c139e12f5fd48bda5d796a407da387e677c0218c8fd0cfb2e509857941304975a3f7b4e391e685007c0c09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf799cc829480bdc33f90183de951b51b299f12b8cfc0e66fc3cdc942145b952c50f01ae7488f2cb162f33b9f78e0da9a1919baa96d66604feebd5403f714c6bf2046;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h664d04840937b56f7c40409c824ff1f355bdb82a1ae45180f35d61d5b8b13ce1faa20aa6ec52c1b98d05f0e1aa60e60f0383c4c9aed1676d3397a2581ba418ff4531;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bd0b1153bc334831de785f2c6feffa2820f2991cdfdcc6c9079a58bfc83f2deb6dadb2644bfac34119ac2facd6e1170648c1e6efc5ac47f907b308f9eff56d8818d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16163a6c392bb986496cc0543c1b9f0e6608edfc08686ae27ceda102fd74fa782f9a975dce414a2a5688c83dea38bdc6659e79b459e69fdd8f2ead4302a4b9d8f5f4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dd5d5227b49e5f499125eb9e1b74888fbfb2a1ff008863b42c4a32fad68663ebf9471153c1fc475a0782f5403848e15c2e05468695cae5aeace3fbb4b6c26b690b8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd4d31ccb419cded8ad553687116ccdeb5b99cd4936ffd860393ca30263da948d3dc36134796ad6d29238b5913f66d77670b2d0dfbff78449853dc509f2761ec31cb8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a331dd1698919d72db88e63c5116940523fc325bd626e160ed52f089a35512f70d62d4a30105c1d672d495bf1546b1d2556a0a91cb2a0445d9769c62d6d875ccd0c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1174e2384a8e85b7bffbdcaf3c7f5cc452f47f872ab8223b93b3f4dd7c6ad4929a3cd4beb5c7198412720e0a9d3e0cb6fc26dd6525d1e666270e4c35ab213d2721dac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac38169a85c2a0ecf8307f1f2bedad1acaf894de2ee65324bb75e44756717e0c3f3324b0530b1099ae7372046a9a138a9236b56c66b93c96e4245ae0b7bf8dadd91f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6513fff11bbfe9e9f6d8293a7a7c8deea5d43cbbacb7371e0d0c71df5f1551ece48053c866dafcb1946736de1175e531f3b0c624d119a1b07bab63d72b9c37ac1cd7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f81d13e44903357c1f19281908965a4d8c932eaffaf55b009769692ced93d1d1545f30e14deacf2d6ebce07ad26665770625533edd6e3935631c51e2e884cc24a847;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5088d62bbbe5d36453bdea40c8094b2ecbbc125a91841c8058ca0c547d3c87dc370f254042110ca43fccdc0922a0ae7a18f37675d823152de3e127b61af87b89c62d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0a918e7a4bb8756161850b66de7b4b3e35b85307f5aa8273489d60dc671417b8ab891dcdfb9f00eb238736ad755596980ee33c288c9df0274db7481430f02d338b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h181552f3480f158f0cae58535ae2a5b2251098a64b0c6d1b6e76941a35357414360852d5ca040a6f1c69506cdfdc13af24e04c28f2d93069ae5799b78909d493d8c82;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc58b40caa432947b183d7a40876c11abab4208ce2dff5983f5eec43eee1464045e39b54c35d0bead7cdbc7a432ed41b179fec9f749cf8c08050d296132f0e12d799;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfd5519698ae0732759f86f4c6a89eb9c612ccdfaaf0990c95eeedd2def79fb8c505bf34ac16e0695850f61f6af6aa35fff48abf65977d2242095319774f219299580;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a1bb0268d1d70519fc55271decc62a21392fec63c8824559d2353671f101fd1afb3a5b2e4e5d093361c0304237b322cfae3e7c2c0922a47b237f3864b15fed11542e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d073938b64d9c674a5f92f394a66462839944d0c615f07cdb61b495842ad637997885ee718a28f98ff46e6067cbe909ac0f16d71cacac29c88799d336f667bd745db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1520454c016847618c81f630be915c6b8016d7785ffce6614eaf627ef5657b1675e7c806643a792fb4caa95a4360af88821ce93f7a4662a493367e69f469d676316c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e65f09c7f68517cbaad18c54c76caf75c4ea5225b1c07d0049af8339f6322b638fd4ad67bb74962d01e0e2b97141ba996fb46d48c08fb799c5bf1c9bfb680f418676;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60f9cbe813949eb8eedd6b8c2d7ca5cb556bb554de86023d9441374408d320b7941cb8f314784a1847eca70faf068877da991823b444a3ecc882d4423295fa76f5e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab1df7c7b57431f80229e44e4e2bcaeb0fee9ddd27d6ebfcc9e0c31827a32f51a38d208ead091a1a655cf33e984c93d970e9beb8c865732a5ea38d26029a91e8bbe4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6293023a702442e7aa6b8ce985eb3214348a670bc70394c5af4d6888b14f77080c724680a03fa836227b97c555b192e47427a9d49269e90cca1f5a4bdad1532ec3b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c1050d92bb273db3c7eeb0a264149d46a88ea5b4913075e1b0cc0068645c906006282c0a3181f994ab3407fcdb76d008ac8b9df2e87539192a7bb954258d859c017d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12bf08e19fbbc6b7700a97f4933264a459f559b654ba8aec956a53bc5b69030f558859dd439f7ce7cf16e1fc6cabb4234c61ce2880ddc8681a2c7b77a2a7f770dcf35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b57a3f28a7d2b17ee40bbfce4f891a5c6fe9a11a6e8e05780705b92e1ba410c4308cee67711b0302bd2ca168ee03e57f41e16fc1696a050fa5a726641e7dc24a35b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ee2cbc6804239dc9bb079a7af065d771263affeb0db9485af2b53195f4c487cadf71c8a155c32c7c67fa0abb248409f99130bf73747dfb8795ee102f1ad2cd77dc8f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf42a4fe64ff0d4dd1fe1d8fa4b9196e91fdc5125474a68bc58ffbbdb01e1cd40796a8e9ae06d091fb42f35dcf2876d46fe35f9c4c323864272f022f341f40a31854d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h418e1cc6720d3132fd17c0bdc28cec43a9712e5d6f01e15b53edc121a61ef28d47cfa16e5c6eb4e011941761d5b0bea5a3c91d08ef965b2048b0cb1d140ed0ff9602;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c1cb841bc57a37ab5df2ae3735bf4e8943fc5e6614c67268406abc891b573e00a109e4203349eed8393305991de2de3e8cb76ba72eda2349dc44a3769a8e8afcfc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ffeb51e9aa1c589efb1ed0f717633dfd939079947dea326c0c1aacc985878648216126f021245b7f9ce6dc4c231745610e0d902c7bf9022e166b8724d945ee332f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a52e4959d8a2b1250923c2b009ffb81c1259fd00002e28012f7789ad4fb2c7a57997f530ee4143c7adb09e74c03420832bd5f8c5d511541ed28258631c70267c706f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d2454cea72950aef163204e0defe01feb6aaea293db8fb9e0bccf33bc7500d37e9396f1bbb841c9fc575666a2c21efa3d6c89f8456f2f5951c8237f5172fa767e530;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1edb9469c63168b7a954e8dc2ead36ef1dc3f138598b839bb34ebb3225862ab1a6cc740be68e9320be1ba19931dfd07d64610ba6105c262663f58cf966f86cf6f0f22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3cb37b542c7d7386cf38e457513896225122730be3c0618eabe97d9d93fa477713c6c8e12a4f6a52a7d0e7bce7f34cdb2144d106409d4b27bee2dd1324d734aeebbb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66f013ecc9e37334d59d4c61c69c47394eae1a6c48e9e1e2c6f4d4c5e3aa2dc6d4b8e20d7fefabd8bdc9be565c97a7d2a7fcd2700e2655ea59bccc4f80035398d4f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb1ae8dcd4e585543ecc0a6eb87443977664bfdf2c8282eb2e8a0eed07fe532ec899465bc9c2730818ffaa9010dc44d5a3c7f7a8d42c2fac6c6c7757da58397690f2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfdcd730a77126bb540c01a159735bcec25423111a8e0ac0cac5a258e1ba4e0bbe5d708fba639a9e73922d1be08f706d1c76a67a69f2e6af4c38077b01ca55c06e8d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cee5ebefb25346b782544eb867fa6fc0d3d96fe982b9e78de32935ce4e6fb5d852800685092844097d71d14785ec92763d8b9a6700a0af13525b649497c13b046472;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d70a685531b3eca075aaff69534488b46e2b6746d41c6785a89651dd98f3074cd6d852f3249b4af5a136ee3da839571206ba694db9cdcedffc3bf3475711d10215f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h58dc64eabe35d0d954661c8100a9399de97d075bf5ef11cc7fc3d56f6f9ee5be173f75ff4f0f721c255332b0b612d6ed642f16db3f10e2b16b46f425818877d3b9e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7df16f0673a1ae28cc038eb74908cdca10a55aa21d936e8620693a280e8ee153ecaeb0eb908e2be94e75f3ae95ff4c094685a47d65fc2c0baab0353b219eb576ef7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha2af5bf6f218e275ef75655c8c6e28c4a0088962e867cca116fc2e57b4517ecdb7842a20130e0132684e56e3ed8d37cf46452b05310d745d191e77f2bda0b44e3c12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13de133a25c7a8ac9a7846dbadb61c19dc280ed8a525ab6687bd12c8c74483b22d4c8f2f426454dac3868258547e3c779cc5602996dc48ff5e003d1d3cd6c14f550a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he535e6cfc146f64884cbda820d0d3208626633e1a2212184f2599c6c88e3b7d38a82544e81385981b351e145b6584e61dcc945f91591eb146640dc1a6a302ed8b2b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac4172cc12c1dbdbac9096b59963a92f085d3ba5e974df1bc799a292956919501bf8c406c3174dbb73d1c442f0b74655f6f08bfedf6e9129e965101030159ba8ad7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h468693e9968bab838236de7396618010e86298d2a037c6a37128b7f022f72793e05bdd39fe7ad6cbe4705c94ca58a9850f11ecf0899c908f2ff6ece818262decbd0a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18e18527b6da413912d893f1c5d01baf3b1c7fd0a5f2af64fa5902f2c393b010597967c08d982b126ec908814751b12afe32c6fd83360f8840eb802da6bff06d73849;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1401d7adb45e14f866b05b7cefc06f78ea4efa6a096d9cd746be9ad088f7e5978eb358bb8b1597647aac01954037fbad18f8c2b336d31c3c17f3c605a20e5d559ca80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1248718ed96228a4a8c22b374ca7f266753b23285252ea20e7e081a82f5418e18c36ba48e3328c4240adf96e123ea46a3a9d8b05ddfa844db6bbc76737bdc9d9ad0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f1ccb0b3562b24086ab5807abb7d0f312c766d80abae6aae61a8408debb6f2efc62971e83d5f7c3e1d11089f4e2e43f91e7c0ea436848235bd6894c9b3cbc6b14f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5730ae0f6faf887bc68a3ae87f7bc10dbf1bba54306d3619513f667ae54ec91a4a756bab3bf30a8559db2d371782eea2e774fce4b272679fac5765adef70503307d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d6b02fad5b59ed7e90099c0073632ded014e5570e052b91bbe84ea6cf1237a3ce83ae813b40e06eddef2d95fc5d14795ca6dff91a5b4b5493f64708296b61779f5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9788bea8bf3ddc4a6e83603731eda71c74634e32d7fdbf58ccdc8ac3a678c3c45f25c57e913c3f3aad5102f17beffa612bf53cd93faf32c0903eb575259a0f697070;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bd643ae4305a09b733b67e8841a5b98038a906411f25903c99e086a9e658db95e5637810bbad771d85d2caec994f4e9d28a8b180ed7e827aaa2582c2f48b7734bb1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133f0295fcd1c93ca7e8ae59c1105ed3dcd96c3d6d1ee712625bdabc5a10966854251e2c2b40f068bf5c56e7521cbada90cd54e1fc6041eaae84690b2c4505b669c1d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19f67408cd8a2e3ea68133542be95472789a4b92169db45126edd36de6da4553e16d4667293bad07fcb5a90e1dad5a2672e6cbfc418da817a74c3c3d31071144f5bcc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1142450b204f8a5776944c4a18605de32e55715ca97ac364a45292d2a51edbd1be3903f411ba9a4f34357be7a4777b516cb636512310ae296d4c000a0a189dd565f1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3190743b96d72f71f80dc97539d90d7b0d517f6643caaf834713b62c7ce136bd3eb9132ed2f4f99ad01fc12bbf2c1520ae9ce58f25a6ccb683f1d8e801317c2cdac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105b7381d3c54fd2376b1ab2c159d0bae9930b1a87592434eb953b336018a29283dd948136a39ee25510a4ca725bbdfe6bb56f6e1ad47717e9e4d1de4db34824915c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bef7722bdb78746236d4bcc1daaec73678d366fe18eb2684666b853440843ba6680e831bcc8d4e5ebbb7a4387793b493b2b72f451c5a29c054780647196e6189b191;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a2df4ad25234917bc3be272704e5961e9e6f5ebd8ce21ae871cff373b72fc66b9fb5e4469becfe14633736cede5e0c8bc4268e5aa7bc46095414db856488a000323;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbdb101aed5b4e07e618b00085fe4509ebcd8748291a3e99683975d0ed2034b75a40decba9bcecf35d55759601f6f2520b83cc8ce51e85b4c6efab6c72a5d0e2b8e52;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b00d3ab549189faa07da977f93e2f638c78251c51458b0f4f5f677bb30bb02eeca8624b8f4606acefc22a0d87e91b9d565ee64cf669396c9b738e15d3b082ed13773;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he162de43b50bd9eada33ee856ebd8fce2598c2057b38cdf6f0634aad6d1c61f1f885db149769a0094c4bfbc8a340fe401de72e5030261f279c76fc59808e36167e93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1712645bf7a89f8224765413d9239cb68ee0b986ff8025401e6b8554b5c2d3ce8d77a864f695025dedc975a02c8ad513fb71793fb60b6282bd6fbd80c46d65f72035c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc8bb638cf548486466e3ee7076a2215ca3a55105fa143d4b9f69e54b352b72b2b0af31529a536a0951031e9b22a1c976a45baa9c9deb7eb77b893371f5d28fc31199;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab97493e18343b53f00a7cd4db164ff857e53c1482c6478c87d04683b1f05deb22e19d7f62a62dc5f8c4db3e43fb37e04e1c490911b698efda89c7441db6fba458c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dfa570f2b34d45ce06c44d6cfaf33bb8270927f2301920c117850c6d0f299fc6ad4ada4ec18b3cd3324c01f5e3ca74c7ea8f21785724971ec4385ad94cb432ecb40e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h47e79db991d2786a7c7a7e227dab5699f0c06d27dec02b704409f12569730676442f799b03b7afe4a2a03324bfd1af4db928a557b095bd40b698a4021ccd755b8463;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha9b27008f7850158cdd5822306fd4c58453951d96d184dc97ef50fef612b71921e10595f854167f3d7eaa105984a98b2ed481fb4d978692ec12bb463f36826f6be32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h22c83e81fc65a7246e63b563cb93016e2634097da9c7c6122c9254d4285ab55638d989a506210b7c7c446794c0c68c420a6b122a7abc6f309e3d2121965fc185ef8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d36fa8b1796774b1362e24c491cc27f263b9f391fc7ef182cfa68ebde809fd8774808da772038569b0053acce9859dc730bb4be73f781e41d04dcb319f2f3ab0e52;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef22e30d59e84a883b8782613dee3257b2cdab75ec0cb0720846e618e8314d7fe9b2a8331c42abc1b1a5979ed3f29375f2daf4fb827f9f0f43b1d2fdcbc9305e938d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d98dd702b82d4a493fd2b566f9bc0b64b7eb765c1d3b2edf79804ad88d55a9719a7e88a9c746cd16ca98f2a2436c8058e9b0b6c3bad874bfbd989a6672838222417c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7657104ba8deda1379f1837a152393512b7cff051b1c53a375f9e226de80170a40b700ddd4439d59171a13c60d64891923d8fd33f3eb1bbd317e3b360171cd2face;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h178e018c10236152d3c56093ed94d81ae82b4910026fd5beb4b21383b1dca422eaefad95bb311d241e2da14d36f7d97fa770eb093bc205770e05ce5d6b4e2eb77abdb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aaf3625ea458f34594a4328191407e1fbcaffab22f8cf3f2c48646acc88f991131095e6cc728e11694ee2d9e99dbca37b24830cdb61a867ef094093dc8f0b24dae4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd5098a20bca887dddbecfbf798735087055be4e6214531ba9f9539d5602a16e98d160e8db7c071ad71819f9136d627943e76cd051cfa4b55e482710c1696d5211ebb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161bb59c65012c8e866cdb501ce74611304d18af7c017b8518d6df093a21e378f6ed16b9ae898a3fd7e8f4f3ae68216a7850b73c852b46891585b08d12d32ea8a9cbb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c60502496c77fb946c2a9f5e1e28f340feb2266628cf67054635d3b5ae8e6f2d053f84fb2a557edfb90e55cdad0e9be6056edf13cbcad663f03f35ce4431f18785ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h65f011b89e6e571a08e76f8607f6bbcb0f62eb5406a603f155f0b4b275c6637031e452d072f9fae164d3b367b5afb686567827c92f7a920ad2afed9ca7021a885867;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3043f1e6d78a2a13e545a999b974de967765769026d68fd319601b7f39a0db9d539db253c9cf0a1e128189f0a327f87c1bfdb0434a1acc45a7b4b0394a3caf61d7a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d4af95e3fa7c2e8592e4b585bba903ecf785d43436898802a0475fc9f4a64031e89e72aca77d428e93b844471ce31bbd2db3d28f967a8b9f0800d5aa68d8d8129ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1412dc30bd7982a49eb622314fd21e9ab3eaa8f94f9090a7cbbe106030bebd9f671d144c7ac6735e7b0c66cb3572969f87191e443c5301aa959feb4b4c84e65eebf4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb549dc6bdc00038c7925772bb13dfd497ad3e027bd2c07c766b1959ef1de9e7f9b777577cf4d34bf9843f146ee831d36767db128a2053f5300fb149074e698d38cb9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heeb3db34488bdc1b373e3f1e07f514a890810cbc0e481fcb2c1daac5a0c751a86825441fd26f202432d93be0c1cf8f7247f583ff2afd79cb20237a843902809422ab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4b972b341c1a65087e17b466045ee045318d38e72023efc45eaeacb34c00c3d76903bfec507a0cdd5ade23cd41aa5a2f0165a6c9f06eedede5d715fd6742275ad160;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h642cff4abf223f2e600e334ab704cd9992c9ec443ad42e883dd8e06b070ab0a405f7eff5f0a18e6afb6fea51b615ed227c983883fbae32406a62c0c2099c686fbea8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb9b030dfabc7aec69e952170e2c1e94a7f65c545a486a12850e7bf87b49cba3f93bbe37fd16b28d5a83894dbf2e6095feecb3cdacbf090b5ed0501c0316afb643488;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h78bc6c9dc209bb6c31bd4da1938b0bb64affb71ce48cdf79f2df876f995de70100d58897a930a052daa4dedb5640eeee965218d725fb0c9732669e033bc31f5e1b6c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb146114d2248eb9d372ff38a0d4be9e3e34c04effc1d31de44bb59421b6276d51d56cd659b232a0a2121d5dd81b43a29caf3607e5c02ddb64af2958dbd762759b78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5045a5613cb762d4a74bea55a6755d46d0bea5b80e3a246057e42ef59691bc4a30e3000e23efef11acbc45de2517dffda7717740306842988f89388562e03ce0b565;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6339e9238f66aafde46304d1c5dca03dcf8b78cf319d74019a8962db3f03aefec2431afd8a670f55d1ff931789c108751132990139e5876eb0b159ee980b8dfb06e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1835848eb59c8ee13d134c1de6267d3355d6e4639a440b2cb9a72690151044d29c53a574556b24cd1d675b48a283c2b69a66164d3497b569aa177ce7f530a58c1d7ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d990dcbee9faccca4269b19274789f93dcde8a6a6a2b2b9946fd6a8f59bf73d42653a336f6696e798262b40dd99cdfe40a310621edd44e65a0cb7f4c8ba850867ee4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h155f4ddaa09870817d4619047c243464111c1e0c0dddd79465dc1ef8ba4140c3ddef04d61267305738df16851e79d9134d22c663da8f59d17600c1dafbfc4b12ec2ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74a9ce303e12d17e0c9af7d58530c37f12e81f25b6cf73a8d59dd4d6d5b14ad04e95eeca7e747a5013eb94492ae18dae521c9e0508202bb26ea590a2ea38bd9595c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6e562b6fda96b2c674c592834566ac778c63276977f87b6858862bfc4a858ccd87b6c3831aadccda6d89775f922786e45741253e5f89ef2c351ee42a927e27d1c093;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f1f327bce7cf33aa957f3ff199db83c9c5b33992cc4a5ea4b0b3f0f60fb3536a2c13ef5e4153f068c7dde23e8b3d048901eb32719322ad0983deb8ec81b36a3e077;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb00274addac2a31114ec9a2fb407ba31af9e9738212da58c255c8c7ce6f51b76a9918e71fa5a8adfc0f55c06261f1765607feb972b9172d09ac3e78160e0fb87ff45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc35cef2f2437240981b719846e020e06b3b4ff70d7377e881be6d69f03f29a32f8b840681f7f8f4b1dc2856335c621d787018be0b1438b94d1b66088c363ee1a1b88;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9143555540069d7bb83849b665520bbc570e22cb333d759d1a189168f121e2e4d60fad1f94c1a44b6532f65b91a889a897cb80d3ee3a9da14184bb8fb2a09b77a559;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14061f82a7df6dc5d77c9b74fae709dff46a7a5511865b58cd9d6d3ef49bf2cb8f7002b81ac005488d8b883f9aa7ca19752a2d74dfcac14ccaefb6c6b2e12773b7347;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb7b983f644dfa4205f09385cc3acee823e02c8f85233ab03d1618a8895f9da614c53b07f0831076f7d0cbb0b88ad1d077443f83d5f39d71fd4bd0ff11dc1fa18b0be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37f9c7a50e118218881449e8705a4c5cae0f248d8b167fb63f4c06082098a4dad256331a384bd706593171d99b5f09119bfe650a928fd009682cf85fbaadf73e81ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3d0a8d56e18ec5d2dbff8ecf06073a9ff087f233b8acd28d15f838152ed738c373cf1e28a75c106869934ea114a4f85c8b76808a35dcff136387350e4d5fdd604b99;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15822bd428dc8a94d00858f447ffb3e60be7152fff57abe0b08bffdbed018f1d709a83a9097ad63392891a7f6eaf7a5875f7fc11ae556fc2f353172eec2b91d089d98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9f0f848aa91c1b963d5e8b6ba9a726fa268b7291a6f3d391427bdedbb74ee0a886d8b0ec98f1f982566c62e3e3cc24d79cfa74871545b53cc6c92b1848723cd48a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12920c03650dea145bf4d85831206dc3f6eeb1dc7391204d86287112850efa5eada87589643e34a53d2704adabf076dea3f5a62b4ac3ecd4a6f612f95357eddbc1654;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7ee287d646f6d9c1a58414b5ebb7858e4f579d0aa2f69fd91a98e531dbd657b7464fe6ca061f4680741ce8277d64791c6b9040b8502c2e338168cd76933f4dc5ef8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha5864940891c3a02e8c52688b40a495d3cd2e0fbeacf1f8c52af9b455ca279865836c02f124e96a0db26e6e732d6e343649e540b322dfdc4b070fe27bc91a981b301;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e80a0010760c67268385202c9672f623a6832848451194578c938ed1a0c1d762574a29ec62000c112d5c39aedd57347cd9a8babc32a7d68f99ba98766c7371bf575;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1084bdefb0f70e36746017023a0487de06e5966b7623611d8d232f91cb2c500bbf567fbcc6af338336ab591ced50fb0f2494ffc222ee70aab302447c9d22b74620ef2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7b2acb1e41f9cecaff65ec1067df08cdfb3c6ff990a6586aaa594f9c15a7c0a90984f6a859bf1a0a1653427e0cd06310625e61bb7915b6993bbabd59d0d94f3a921c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h30fd70873098e5e1b2c54d0ad387215dcced66a0fd1c6f9fa4324e2b6574bd7f3ba29257626282f5e361a7a25cf035737ead3308e0fd61ba9c5b7b87ecbe81ec8510;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37a435dc782fc8e0662c491170b2bc1273af39660c8ee219190bd39f5d22a2b3c7b54a5937a8a68d0313477e8f160465c78f32521b65ed7a330fda5cc927c4cd1d64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9411ab6de21d9c731d10111c33ed1eb58ead594fc6deaf7c81e2f0cf77a102bcad5de38bfc7cd7016b1ff267b01b3cd4acceaa7fcef8ed5137496d3f6cccb2e7f4d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8eaf038b3030c5f0e67e4cb500f6a5734e8d067a276f0c5e1c92a50fbb3fc5a771e06df80428b9bdb0d453f36a28f6383236a2e85ae0b16a07f2ccf303e5d62720ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a24c5f521c7e7d6044a4314a23b4c9a52f8bb61753ee6df565400ff496991a33dd6c00ca6452fb555e23cd5a95e87a5dfeab041c830331b5add6aa056929da78f66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16072d05f1df8970db5dfe8f7451cd0b0e4a7a055f92d1b520a96a56ca7107b886330d7a3b4794b269590bc63c9330a1d85d00237cca3963f37d1a92c1e7b4060390d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc0c53c52204f21a63fea451d129d2109ec7007b2b5bc4d5f3d04022004322a404300f0ae8f790f39c38f027e5e23869fa33325037dc8a2455895e00723679e6adfa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd440ea810fece6a2fb36be27c63bdf926d6b5c04f48a730afaae49f9e96ea7514f9a6f8238f3986164e373b4b4b90e287f2f2485475542fb51e947d02d1a09a30706;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf47b9d1123026272dd8070300bf9a02793816c547713c75f7ee147270fa6a16769cba9602e8c55d4d59d777a7c7872030d820a5823d003d7aa3fd93a4900e0d316f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf5198848eb9a23849e9ee6b44a8537a5be08a0659fef418f0220f352a1b498e46b30f771e376807b2a0eb07d47f777eaae2d9e3549488888fba3e669e0ec36635faa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150bf99c964475ae523c9e02f8044aecb770352cbb0b1c7073f7ac8b9710fe0052cff919536e03547121c5d94f995fa41ddded968c4ac9b3f6347707bdc579882fa55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c1b148c3ea9ee638a505a343c9662496f01b3b2586b9b7270c2b890426eb1919db80a83535e7eb3a8389059dd330371e809b6e5814f54574b5370bd6aad082014e72;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d2d93400628860012184c0f2639d11632e156a3951f575a471e936f52f788fb13c953deeb03c5472d782c640ba92818b9f57c54025f70b87ef63accd699d5bfc231;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd76d1c6376b3acffafae9a86c43c90bbb85a6345a84a9e84ed40f7685680da63ebeb07ef1b80d27ee9d7e0c881a0418b0ed0afbf89779e031a24f6dff343290def0a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h100d63848f34485aade5ca2a542ed34b719968d91614d57d6e84f2d43c792cc16b3cdddf13c8c7fb1d4e19c67b4bf7743b0e1bed823e19e561dbe76341f5c751cc0a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7851633ee7c7d89b2bf050fc07af2de4a4f696be5e4d2b62dff3a08bd71ac2c75fe2c2b68b236843b369a73342cebee756b85dbd9f4ec3da2ccb3b7137bd2dadda50;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18db3ee94c1dba65fdad39db04d4b99c813cc026f0adc40e02794ea424ea674c8e0c804036ec946901409ee32ae05c1906817096c47b70e77d3a5a3d74cd67c796203;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb2d94f9a3f0e60f16e3ed9e04363837f60b618fb1cf54be26d2d01a3f11b79835deea05ece7551998b8ea7646fb07a1a9e06f76a233cd6f6902224904fe1f3da857;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a58aed09f2ff2ecce9133314c3349e730e5a3e864afded5fc614211cbbce414fae9ece928e3b397fb4d1c45b75031c4600bd822d1aeea64afa7d8a56aa625a49f0a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14af75a8ea38c3876d02db0ad72346c3c8e8002aa212133c74135678d49bab87dc71174ab819a18b56131f0a6a27534349f1e75535b746cdb614d4b60c743841bb908;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9d29d72a2d4c3e20a0531338cb323cd0054538ef68fd8e6e6b90809670c1085b64fa20a716509da56e47f32229d94d667e090170f3a6c0add51ba7a5932e0052172;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1749ccab7d1802c4f6b84a5c213f8c34bf5a65735ba77e8d037bfc9144755bc5d7d41d9aaec60bff14f9d6136c3b63c0d106ceca148e097da79398f65a209d1bcd126;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h176265dd8044f29ee5dfd164726e491464897ad871d022b916111e419bd67ac8ecc941b1d24b6f12b39dbe1adea9692f178cab75ad0f49428563ccb7069265af4bddc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161995715fa97e64443d89e478005883af183c312c97ea68d7d0f3b52a129eb97f7308c518750df45ba1daae25222d3b7c333b3b795622245abd545512c0dce0ffd2f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h82e87db644a4d2c1d3650c0a2bd6291aa67d5640da10fe3a1d826640e602373b42f0ba814297176742881a1b12405c8a75cfa7b8acbd9b47787adce747f875583798;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1972d991fc606f68856f8d20652cdb787f3342736575279d9b965cccdcbd3fe3ca4f09ab8b3e0c5ae39bafe38617e869abd4210078a5a80438424c4fbd29095e2b1da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34de0a1d4bc343bfcc463263f3312838cf4472e1d568daedb4c65ee06199838287aca5c5ccd380564d8f57f45036b8bc8d3216168cc46916760c529ccb39328c75ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a9aa48697c50bdf878e042717b39fe3ab09c4c72d3034e3aa5b9d76291325224559855fbb0b218f0e9906b81a4c2e39acb69d38e885e7ef2be221e8deb825aa06fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h336409ab9b5733392723ab2c607485df05bee318befdbb20bb0ac5e02697079a89bb803a163c254db435aacf274e20c26d3eb0d0e93edbf3f5f10a6ee2d1ad696a4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194896abc9bb05e83c9300280d94da9646790180627bbcaade2f21b266e67989d0f4eb9948ba5f701cbef36e8f77cc0648602dbc7e7d956c16443889808d821d2501c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1baa57f849cdd78ac33d970f5877814b50f56ad1c8c1eeae5ee4f6b73201ccde4131ec2043647eb55d894f3b174873aaefcd117b83332320ecdcc8f92e266bf091e7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he159237328bd10a9e2d86ca523500410620bfeb9b2f927f1e343512a68f6a959949b94a2ad6e299db60f8688510516b681e0065a737d7840b2e460113eba549c559a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d7bcc9b1c03cf8cb069f8e51a8dd35a916e6dac4945c2cbb8b2d71394588e7ccdba7605d088c04c742daa04d4b41081d9f8a6e28c6f18e2a5702438e636d85da9cbd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe207c87a9efe3840aa9c96bfcb2cff4ce43bac12d9c9d3b9487fce01f25ff43a839f18e3e1a138fd0fce58d37072fd2560e8caf7ffeffb4501d6062335125e3a5ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165cf6a3cc1a52c723b4d88aa97c6558524adc7c5873d6ed2f5c74df9306ac17e904a05776bd8eb3670de6813d2c63b51b29b5882da7cf76a9e67b42843a3b688c72d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f6e3a255505c2ebf7db458a9dfa8e7d53ac01f2f9fae851e30afc02384748126dc82a495f5043740ac8d0b1eda1cd91b903e276933fbf6c6315bc0a10b1b2957def;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14245d9c3f7d7d7db6bee2398a08fd1cc1632bde76c5e12266471a37fa34ef6a58028b3d52551a8e86278380a960642e3ae184b794b2a88da43b992179db6944a33cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf4ab46d5723c17a748500621a051ce8ff701f309ad805209a6803b278ccdfe2dd81aed4d286218177c51e26653fae67ec2f57b9dadc5210b2cd43825e65da8c735a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6748d168b2fd8d54ffbaf0ec89c160e0c388e633f6645a84a05a35f86913eabdc59f944d154ed8e44a0bd61cf148ec7cd1eb1ac0c4d595f3cc38bde90a8e92adf73c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15ab968f188de5003c3cf75a4d4f98ee9797a3ad59d435f62d3bc35e6c0d9b5e9552f35412c0513ea491d6e73073949347322ff6678b6619f118825e5661c3af82b45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4d8c09a60ebc5ffcd895611517c63b40f3403b9784b4467a2acc1efdc40a3c2764a893b3c826b6faddb85c9223df00b34a053271b6f6ebfdf0448d4878a36760c25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a99239e8e7f852c66d3cf8433333be72b740d37edfa18971596107303d1b3085a75ae0cf223ff2ae77eda0f8c9b39cb0729a0d309eff66ce2bbba45ce3dbb320fe9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h172f9d88e2828e302c33f388d38063bcd921a9cdf7518ba72b8f2270d6f3fcd0fc68aa75f4bdaeff034ad1fd649faf63baa36aaf57e1bc253fe1e7d522b7e85c100f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f52b872d3bd629798b3ca23419bf1d533dc42627f70a62af603ace323cd0c86c0cdb866fa76df8de4f40bcae456daefb8648383db243d5faa66dba8eff6b2bed62c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf9e4f426bac95dec80240c87aabb15f1abba550bccaf2f80c0cd7164defcea59867fccff6b57cc50ea3122643f80bf634e90001850e7de6c58f2dc0e3a66c8dd9df7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14f152a87ec6e742fe9e0501442f3c7c0a5ba1f21dd766dc734479f04c170f2bf2cbfc993a0d7c020429e62a4fe6292e5d6da869c29812f8882fd4d030a05d3d3faab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc76d40238bc4c56bc601079a10c366299929c98dad5c10998ed9581befbc3aaa6466d5330b571930f77f7259d5cff9d6f00c78587bcde96f0b5e9c33bcf33c971a67;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h329ab539122479681c2f4a8c4d408497f4b4ed8b6b7961b4427b0b6fd30658ab02426d891b3152ba432fc3e1131fd4dbe74d91ad88a016db54c774af07d8e5a126b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h84b897ac11f5df2936e19e3a83bafc93142dc012430dc859caa82dd5c8d24d625ffe89ea65f66c7aa7758a291791582a7905379cb090393c954239a7e6580a5d7540;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h717e7a0a8a7c3eeb249e2d1c9a01e3fcc6b2ae5966f061633b8a36c683bd5b1ddc1810dff5349eabd4c189c7fbddf7110938c5588d7c138579565b3ae1c330de57a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h70d7a02a65566deeac0f5905b3e49959be4c44aae780cf3af82f88ddc6ad46dbc99b7aa3ce230276aaf8ef8dbd549a1494cd881b683a84c339c9d92cc149170ff052;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h646d36bf17ed53c9ecfaf3d16ce91954f29381be3e81f657bf37ba67d6e3e92d9f3c4058ffecb5bfdf9f3e65acc36e98eb7bdb0b0c0a367d158c056881bb7e1abff1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19978d9c754aa782c598947dc401e580ac9db2c91511fb2578c0c9cff3ebe40148a0c49c5e5fa036134fafbb173108f422adb38f825aff2c2faaa5c92833ba3de7cf8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9737e269515e441a84d6870e73e16a03ecb0304777fc67d65aa7eee8c836934506287711cc4c6be75b0491a925690535d5b2b2cdb90ba5c6703059f44ec6dcadf1c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he8eef857a6ae5210bab10b4d5a543f2c3b190f33b6b68ec2001addeb71dc8033815c6ee3b4b7bcd923a5141a42ed941fe064a7666deb7c8cb98c4d0761b5c9f38735;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfaf2d50201683dc897d4f71a75d0e4c4165f460c831e6ce9d8c027f9c8bcff2696809968b1c531186c61fb520a708ff80b1f3211379f895bc1137f7445ad4ed16cdf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h72fdea335c3d8604c04155a47e2584885127587176cf9045bd191e71d27adf3a58800506d03eeae61bb93df66bc4c5f8eea9bad68b574b22e37c67dae0b3a26f233e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c4b5a7cab77f4ed621b2f1e2cfb0ff718868089727de58561cf6656df6e3d0f4794633a024583d103a844ba76d47759394be9db41d370043b0e298af43ecc5c31b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h174e1bf98b0ccef83aa045dfbe35d3ce2b014fbb56ca47d708de38fcb8170c5dfaa4627fae07d3ff6b259a0172cc5bf988de7c500616553cf5ed2bf3a4883eae4d599;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f89c1bee30f31e02d0bfbd5b591e2689a0c37b33c5269df47a7c787d0f2b913fe9118427a5dad935d56250547bbdfff1b928a4d9fe206acab19f2e38ca8603f37c63;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha986e0c3e56ee0378c1e1954ce3ff29c170173f2133d8d81df4d54f0c292bd217f9cbcb3e506ed15b91fa821b07c14f1ba2204669c5fc180097a09c9ee7db8057621;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ba1e8e9512e840738db46b9f4a99a9fd55994619820e6edee47bdc9b431840acc3ff8eee08a0950612112f40a2dbbfc68535683a959190c82614b536b5c73b7cebd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b0e39ebca2b4d900265f6e87e512e64dac9ed19b011a532139aa1cfda94c24dd8e6abf7d0c897143c285c4b2d75c99b4b200072c12a53c6391abd2c9b45436a76848;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h778568c3504cf93669e57a7d33373e2928dc10c4488d48ad0c63f857f17b946bc365bf7d4ba08502d8c1725eafbb80921577569590a16045029aa670b5da8c3d5a82;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b0c8f961dd9cf78df2c01127626f176740961414e6122ff600268928a6100e5fa98d3fffdc72d2b4ad685af82560790479a7604e3961f19c77ec0e9e38ba8bddd77d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eb2b0c96ba29a81171c05f11fdeda5c09c7336183a09542c1783909a96a42f00a35466c2bd4f2cf36bf01acd2805d05053e7b6730da415c5ae45bdfaf19c9663be45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc21ff7713f8f9c2264309f523906b533ebe618499381e7905b361aec271bc0d9864112025c141f5197657f96b02b377a36209ac961d062a56a8704ce139ff750272e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10907a73bb562cf8ee1ad29368322bae861e0449e18aed5950890971886b06d5fa2694eeb3528e16c1fcff249ac4b143c23b5608a12f9d5467643c9ff55544edbd2d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h998697f94d0a6554e3d52b3843e017a29d1d48e93bd5db93832966dd76b0c5a6243524a98cc358c6e8dea924ba14059775a2b798e57ceca4a0b57c319673de5b8d09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h109a2f34b34e2b346c30bbd30e837b4b5aa9b1f5bea890be3eb6e204b2b23c36a62d9bb8d67623d92499007e1d5fcd60dca5752bf48074f7516df355d42269bdbcc32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1194f18c51ecc3348aeb526d79dcceb3062e91ba67d1b10dd45ffad4e2b0d47e99045e79b2d81dc0697bc2a4b67b4e03dbd0c0d4b9a4bcd68afb78da12a365c161537;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5a9e2e4f3bb8c39f349a93885d5c4afb7da7e965ca71f561ad171f716f0cf41b6a36c51762e9cd88e35c0fab0e1696b7cb769a505624bdfd6e89e6363907fcef4f56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf20b8c62f5d49bddf8570a6d3637acb64f3f8b0f617924766ad21ea1a3003999f4dcf98242eb7c7ba13bd854f8d8e15e3e59338040329191a95619d1cebf9631aa29;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca0df44acaca20b399d8a544af24c18d11bde35feea72a75cfad4fa6e80e62e86d8f3142c3a9bc131032f41dde4e65fcd213976433d1ce7bbb0f2d036bba08af1705;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1caff04b91cb9291cf306d9c5a03b03e5472d2d488638eec045f19499ffa88b8409e76cf46680df7ac3769d2b6e1af8d8ca66426ab8505eb1fc1764dc60398a2ba2ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aba83c1a72f62bd24c7cc011c28320c637ae28da4b5ca8987c3703a6b3d030b28927e530707c1c4c6c655ece80d43bfe11a4bd1aa8e20d9ad32c713fa8b2d34f0289;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6140c96628112d6395f5b37b617ea1a34e118257f3fbfb4d8c0fc8746eb6d4b2057bd92e303d85e765b33719ec5acd740e67fa17691906b241e62543d77d2cde982;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80ecb47ec7e082e84f4c69c2b96690ea1343192c1cd2b566602cfc7f2b28c798d9fc57a47e49701511a4bade750caba46b54a06948173b03c5c4d696eafc6453306b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89d1d1aee13009ec2b3ac8cc922d99be401f1aef693061667291d586bb953ab26f15154898f23d09f310ef6e10bd8f8f9692f2df4dca17e67970573a95dbff484d27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c5d5db51ac85ff39a152558a8c416816b8369ccc3b4c9717b70726a35efc4b1b5d3d6c036c33ae60855a13331541a124bbf0c0e2cf31f2cf9daead627a47733fbc8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd61c19b43db62ab69a9a2f9bc98eb46422df65a72b048cc225b06ceca2c7a8d74d5a5ee5544b9da2248d200ab0e422edf202c71ab2c0ef5dfe7dd0c57ba6748b78d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13b918b3bdbd3477423a8fb5ad028b42e6e527dc6098c51aed664914e666315cced4b14fb8b2195ad860cc89c7686431150f646d4a73df6c712c3c457361f6baa15aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15db091a464aea883dc97420252fc70407c85a5afe2ed407319c506d9e4badd3947596a095ca88bb89c065eb3d32a20e629ebf728721e2dbbb5e99efae002e6e28394;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90a24ce232f74dfc2d315fa6d5e97edaa790af0232bb719de99e3a9c1e53fc1542238a4f700035724b33d559b13ca3819555b36b03196c9453af5c76b93cf4d3028d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9dde4b965ed85845fc73a10f2fb3c310825fe98fd36f37f2bf44b710c45f9bc7a9a4b116b334b1bf22396112ffd1040f2ddee22a28afded014be35374f1dc514b8c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h141d7b6950c1814a67f88da3923647f9399de9385e42212599c6121a8b1d8acc58b5aa29075e557d05d40c6566f2532cf1241e8e2f946655dcb0b1cd9aab91efc9c40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1676e54936bf581c3197c3a661f40e9db4782a214e022d31fab4e899537bcb1789d98e1ccb62a848691e22182179b906a6eeb5f77f191219b77bee0b09355abf727d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14bf2dc96d0815fc9dd0458457ab5ba095177d1bfdc8b3488009543da412809f155a9fb3704b01a807acdbed72bb6350cb54e5328f53e3f2ca8ce32660cf8e5b87c41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f3a57d0be0b38f57eac7a62d108898314e5a75ffbad26f9389e7a92e883d089e9d48b515b318a726b8ed7273048c5612cef22119a3ee2a4297ef52d3b63c7c6cb4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a2ce3ba2bf5c663777ee5a50f60b2cec1a4be836baa4fb38af354711c4b2e6955d5a2d4c5e488f5e8fad3b46b672b075f152deaf882da86b8593c600a7ff0de78536;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5bc89ce409cec3a620d0c3890c9b4b603bcb17d691c46b459027ece02500d3ece10486666c0876672b81d79e77e5371b2d0f881d86b2995ee0e15da5b308ce6fcf0b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c11dee1a92bd143c6809da9ef2da3bf22dfcaddd8bb2a2f582a8c09bb3fce22c6a66c549371548ce7b073447089e27b509fe37fd97c2566f9e4f5f71f0c0f93c5f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc56d4f8ed346f2e3dfebac72c5dc761ed6e246771c6091f821a146a5d3541b9cfcc697d820180c86c0eb4c4ac1af3dd093adecb811aa5b29496c009bd4079b0192d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d833d516128fe638d1ab5a12f79036abccbc4da345dc31db693e5154aeeb490954f7972e28c6d98861c0ef504073b75597d59b3e202eff02f5e37009746ead99c3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2f0a35fc4c593c5e5721a973f91b894d457e3e45b30a4a11522b831407a3ac972b931e86c50a3f5debcb83b12857fee02fd53e18f3811446d2fc65ac5a3d3b59e1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7aa19357068f18885419863e768d75dc1ae9a0eea27214b7e8bc63a94bcf89d959908cee49fd301db9425ab48908eb6c370cdaf511e304b417c7d1742629737ebd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e751b2b0e471d3bed214c81f24625cf6d3bc32ccfc59dedf1aad9d90ba9d382d72560d310cc1a213d1d578297eb62dfcb4fadb7df30edfdd871e7d75553caca87e5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a8c78ff269eef1fc8b7dddcc8346034f7fb150e60582f89ecefa2b92e0bb2aa99428dacd31bdc612b9ae2aa93b77425af32ba8722dbec4ddd2011ed0c5b2220502c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13cf8baeb18c32ad4a88a2dc77fecaa399271a0c60a77a0bf4d4e38116dcbdfdc3379521b1fbc342c804173c6f5e3b8e323573abb173a40e42b38d279a98fed19fcde;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19ea219c561654bff7e53b86ca0cfc7a0e49ae63f693a8bed99e4667a4821a8689454471e3aa6482612ecf2973ddc800285bfaa85504d832c8996bb876ae201c338c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h23799c0b102ad90a4d0c5645ee0cddeaf353029c41ed3ca298412245e0ab21e970244af36218e89f3ab31d263712e86eead2e17529e8050be5510b896af23b97055e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19e5b59ea940a5876a6c0c4a06b1aab6dda67a33466f1f0efe83ba61a1c0aec07320ef0e97c1d086b089d21c0899d4bd64f3fc33ede75cd2fc62a0b41b3d62ecafd2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h29bd9f3bb082f68a860187e661408e544be990d29449359d9ee92f85bc60af2da7e170293d72fc6ea29af55cc5f5e58efd03ae5fe4d8421752673dd4a918e8365819;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3bde947515ed5c50015dd788f6f5f511d69c717e4640d4e93e2a1aecb8358c2810fd1621fe3fd719be67d26906dc2a1ccc5667a24b5ba2500a7a0f743672f425136;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h55a10d0ff9256e03cb122b97ac66a26ebe467a560dbce6207209eb8df769c11de0fa26176c25a7d16be43de5e92a3e3a067609825cb9347948c0f043759845d9853a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1187aa26d81a8d71120c2f84aeee103f0ad1036dc2fedc45a0367ab6831d49cdb32302e53c1f85fe6b942fbf7f3b29ea76d0faf814450d7505976322dbb71ff1f2537;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f72170f4739d45682c173a1e88f3e4192498242c566ff7b1db7aed081e71310a344b9afe425a830c8a0a228395a28eacb5935b398cde0cadcba135e3946363862422;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa240c6e6f9080ea72f819c30855d2be60d061001fa986174c5ba88328a27e6b25665590308fd198ab35690a07a4c6e431af3339402d134c0bb109f889b5b728a7da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f65ff1260074070366a27995f941a7ea86cdd27ed25ed0c1eb2a7d3b952823dc6a56afc1830aa654e9f6a5442a6702587c0628334bebf50015f10401924a8f90afd7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d3c5f63e859b414d39e0602bf042e64662d8c0346000a2fe0b0719c0bf897d9ad165bf7b5f00a3ba47766d911eb809ba6eac00190ee724a136996b240ae98185464;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e9f7e4a43852a66dc807be9e0b8f9d0890a16ecce215c399f809cea8ecff631cbbaf2a20478870268543c46ce48f53b760bcd4efc84e1476750d633cc06dd6489af8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h35375be4e27767a9c7139bfc746ce5e272900bca8d29d705ddb708d13888e55c1917764b9961e5ade23d2f23634a11341666c425ae2a4002b61d7c3d01870f70912c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c2718df8a1dd40afd78e62a053a624303411f930c75fd37378e66d33e7c5a49023ec7dcd03c2ae4c1e844b68c54a810a9bf8b24f60d990eb485765f7d9fd3a67b2de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha33dbceaa85de811912bc304794692c2b6e34eabe4ce7d11cc8c8ba2bba4512e55d8f5fe311eea36d7223521a8eb4c9fce179b482cf4669344060a7dd0a2d9d1a9b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha8c9218d6c5fad8a505b1293360c2282bfb9b37b0775f6eb2bb5aea5d338570ee0ae18b24893a55f649063769796091ca2a2357fa103f68e183a185142adfcd5dd42;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b96f23f90d595f18603b67bca2d39bf0002576b085fca2501aff626bd153fb7ca1445cdef8792afec9db497d22ab7075adc53f1f8e423fd53a8c281fae39cc0dd8c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15677028df92a769e8125af30bd35c9f61b9992659d6ab70e9e38a0ef1cd7ac5b5debb0f6598ed248103b95eec387405f4c14662dde25e14faaff607e7d784a03880e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2ca8a6f6a4b46a9932ea164f591627fb4ef80cdeb0612becb5626ef4391085ba537a55994144859bf3be86769f953c078fbe1ec16708aa653da14846e494994421c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3724d99202453c2e5e4b55081aa3c87bbaf0e7938013523cf9f40220296da4583eabe4c34c2ec47598e93bc006c8b52492c229ed54c5289672c6c6bab839b58787d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h50167633c4a56d9e45a82c274859ac2955f9f6ca100e063efd17db13b4124afb4d5d3c08499b56e1a72f9e408f36042b16b6078988c48294d3269b2942d76bc947a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9c8a6f33758bc9abaa1cb2c3942cf03eb09ca23379647e15a6295d78e30a09d31ef38065caedac447c325a3a7d601d78877921da99a5acb01e0ee8bf28809ed4dc7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f72bea1797d07b380356bf2992713dd6462a7612c2cea3954ae7764e51af58677d598469e88249e1be485f3059a47827fbea6434520dd2c0bab04c89b64ef96584d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb3e3b2220c6850179ccb67d05ac81731f815160e8fa84f7dc2044194c0e5b5744218da6bf5b0c3eb0bf943865d2622df7dd3ef4f4fa5fd02b7f7d3e7e5667533d33;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1447c5d9812f1f187ee8026e9ca87f0a8152ebf7a85c4a607cfe56b9b1449974b417ed76dd4594737605a02831da232fd63e6c5103bf3685146bdce2ec1c11e369f98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e607103c428f6d2678f3b6de318ba7f24e0b8aff0a9cd10bf1ab2be216185b57f2c1a4aa288485d1e17a7582bdd80d96a75b3f3ff8490d38c7f8b620a07262adf2db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19726f64ee0b58cd3f683c665857147f82a507c3d424f2041562489e791d22c19269b30e044f5ad5b52f5029149fd8e4b1e523815a00cf2d4852e25cf41ec67bddaf8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a26bc576049f4ea3bc5ca2b735f3dda80d5bce6fc066c9b5ad1c659227c698660d32317caeaec8ba4ff6387cf4976b2b0b9319d91b31553304e755e961a205aee301;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bc76b311d82b8ed6f5b3e624d6d1dfd815fa99c984b93ae3e0a81cb70d26e019dd913b18debd32cf6e293933d0a1d23c53332b3892eba4d272a0b635770f5cc4fee9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a47354a6916de7dd764e13fa7b1b3a4c4be6315dca201a166bacfd0886c825e2e248b6e90eac6e8bcb08ee01d150787e71c6cff9e5bc3d711f74762e8025cd6aa87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9c413056fd255a1429613aa964ffa60e0a945647e80d9f7893fd3384c9027996cd74b720d226bf84f643642814f2ee5be50357b9123fd65d889a22acdf752614977;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96e8b8704da5d851d1ede00c856366e7bebb0c8ce8cbdc75b3150cc8338e22b00f84bcd205fb7824f97443531f4b0f7ba61f31935ff3c740a552a894d3bca08b3854;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h158801d886d6f609a0676323ce803d397d30d3e6c1d3f28fcfcda6306aff4ed5d5891662e0ff14ae026127b39ba729245a002039d7326bc0732567bb3a329fd1bbcaf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd74d878c4ad243b0f86b3609ca7d84ca2562736922c432c5b69e603f878f436f9b196edac9276d08ef880d08882312bb7a543b94418e381a9f5e43822ee3ab501f0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1abb6d0bb0dd8ffbdbe095096d61c2f1e04cac1529c147e93558e347a2266e09a62299c7977d7f6af361f6c656dfbbf2b25e73cc3a4657bb566d83f08830c6aa0d8d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a5e1860fc81e709d771f70323818ed82140f996bbc7162709e7e970d3cccafdec23e4d7441ca019d91157003e9be02f37a7686f602a04f18e056a2579a83ef4120a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0d839bc9c217468b7b31c82432d1650a7d346be9a4de511e2759258c6cdfd4da5afa119ea55ab4beb2a2a37008f8750f9a08104b75a66e57263ede8cc4b7dbb75f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12e69a02b1fd67ef9810f069d6c314a4a7012a7f65c66903269d560329e736e6326b216539ac1a88f119e24735ab641060476410c0b13fc4f2940103c1819c8362c0b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10617094a21840a5138bb3d44f0f9fe0e216ac190507c066fce23e64978c37783db9327b9dfb1836ab7ee8e2608fb54fe6236bd25fb1c9be4a29b77d3a299744a35d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18fbb8a3cca53159ea2a531394b82f4f354f6ac0bdea98bff115f6758238c2cddf174a40087a55c5cbfda9d0da15f3c4e613dc767c5512aa5eb7b677864bfdfff977b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129cf24c0a269132822f854a282a3cdba6772dd91e7290951cad57de1ced3666f7a447ecfbbf56ec72d7645bb88f6179e20340e98c61afbc6ec736889330389dd0541;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13aff92d505d48874db35008d854031216712594c9b1549a5eec36791e15e3105336094b4248d06a1081cbd59b5255e103ce339a504ee2224754f2b001bc3d04067e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1278c1a121990c0e9970cf4e7cfa23436925599d0738c734e3dfe344503ae7db1fccd722ddfa9c6564e88affa1502e95eae23285f8abb1483b81e32006e0299b1d01a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha8308d9b6b0c05da2b43995ba345e8267047e7001bcfaf0116266159ec76886942c381c3478cee3f787c8e087a579c4e1134d2804feaf96487af04b18880e0d7b44f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14357f9c43093b2bd9b1b09e2e5923105c9b3774f030e2f93d1d552b0ac16b3e55066cd71681e07859bc1175ad5b1f12e1f840cd08283d42394a59af5d17fbf607e22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hff24ddbf015cf00d235a0633c956fbee284a05f174f45febd772e35069379b548475f6230aca22a76475f8a6427ea9b5ee3c2466d5d33292f9f10ad4ab23a55d3478;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5517fb06f9cf6b1fa4caded535e75d20482a8e1fd3559c7d93d0d4882bd67190caecf1a4b9ca0e9b9f64632b5d682d9fa336287065b572a12b03d5b8045df46a5559;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1519dadb78c48bdcc5f582ef2908e25ef3ab2a4a68f2b897fd8096304554d9777a92b5b598b0bbd88fc500928bd9f207a4975cc914ec842ae1c76194cc20e17f728bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d2eaae4b0d9297874170ab74cce42208fe67fa687123c540f24c37dbffc47c1163a7a5ae840dc0b01ebed859a0ad7c0ae25eea021b9dc049021ec1aec426442a098;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3740912ed17cfd1a360a8891ba1c04e47f60fd246285e079e1cfb146e3b6f01b95b05a1b6b87be1d913ff886d02938ae3a9c486e7f20a0c8c0159f7fb05e5905526;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1679ba985a521a9829120d92258e6ab41f94a569654a3b44cedaa660817aad5dd2a3161f07e1c5bbf80157791efaebd4136ff79e49c933bb2a2922f87cab4c5eff411;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ec2dc5313920ef8868aaa5bc10c8f2c130ac9e5d9693aa05a9a47e5c63863ace01879e6550620024d712ba1a5cc593e2e2e1f36e8d4120e7ca6b36a778e964f47ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7bc84b0350ea3c43d90df046c26bf78e9e6cdd3c6ae827e0eaab8b755c2f3f5c537f8388932c1b60693993ead8354a2a1f64c52133bb6a2278d65f3b89663e15283;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hef6eb2d4fa5047b19bcd25fcbd541ea7b98764193fabd361514f52b1f5ed6f9651d002fd7ca483ba8d3de64f2dbc44b87a945a6b448d90b2280c43fcc4e5f1cc290a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h142916ce07551d2324c534d28f5bad1c060225beeb559497d608aa4d69b8da9e0c56440c03fd5bfaa81d585337b09e692c4ec6bd488f311c7eed5403e82edd0cc4902;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1803d98236e098f0be6130bdb2d5742e17a92f6adc4b3ccf5c1e639fdcdfbf83a6458e6a5ff53b1ebf83c1500af6b675d07546e3382b54412382f73d2e04ae2f73847;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h188ea85ff472c2d86a9e766aa868c305657cd7080779e72886d4a718719119e7519ed0a1c09a20d16d86f5298d1cffc3f544f1cb5c931a07777d53d50ca24988338cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea319797a968f99ca281f42dc41ba744b30d43b4688dce202619a54c2eba7b0e5272e0cb0c5e061e578f8ba0775dcf65c6e9524317642f6404d9042138e5a62b88ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3bf3ada0fd4e20bff9a243d63f43b7241082d4da66b3089e3a49de47f722a164b9316cd53148e805e5ca0a5e392ed5e85f0ff17514d50f26b61ca3452793562d10ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1959deb30394d16410104a3545133faca3423681f62d554989d876a4de548a6b6712256a073ccf7e3ff07b1070d89d8e17280e6062987613f7ac90a02381c3655c068;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h72e48b434fb21ae171c40a1fab51db3b7e37d977832ca5afed6c05bccd6c851ca2c159011d5dc3ea3bb3288ec420f3e42e2fb36606452064bc9273b5079ec139d472;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118891a22b68f0be4877eccc75be4deefda44693e7d55363aa019fbd2385a678317e6c727e3af201b172b4d1265a4acd9d218d00de2043d6d3acfc295b6cea8ac794e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfff523d8ea969cf8e6a7918682d956105c557d25397836377ba174ec9595ea5b86edad51b6b5137ac675eb344c04355a8c8c4a7a2d40a01e985ff9013901261fb6d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h58b17fd06fa436fc9ad2881c99c2dcc6b1d293793e9f5d192801b640dd06c6df20ff09e1407796088ae286035d3ecaa9240b70f63364a346e5aa837655d276e5b87a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19015a7ab36a9cd4856ab61e13784ccaa5f80ad8c975be93cfd2955b679023fca102724be31dbeeeb86327d89c0dec3bfbe17f92fdb0b9f519640b7fded891a30482b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12e0c538ce68d89bc252239bf5b91c94d50304f4db8a13ac8467c00d4eed1dd0cda60ec20e2b276b6554d2f72187afc45c594c1c3d0fdab97596f95c7b8379abe5df8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f505f368fc580c1472aa907391bb6d56aec41017810de8bb912d145ed7be3f7e20bcb70d8beb621c83094e590baaccd2169a614ac1fef537541af8a5bff93d5498ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f2dfbecfb51bdbb7c3d4c9bcc34c271583f2746db807dd8db717c4e4b235e606ac82db9acb8fb3f70f4b3a6e38e77831facc869c6496600ba55a92b4b3f395092c24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165d5584dc2f576e21f3cda6561c4642acec0f72a3c0b577e87b5fc3e0dad7080508fa619c1a830b5239dc4a476ca85e8161c20bb11eecd6bbd44565885253d323b5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd665e9ecba65a08de94bd939fb9a5986617cc3358bd5b8de87e3e60faa26276dbc1741ddc468e2d9e27f0325fa20ab3ce53910730fdd6ba796d18cd65fb1ed18f81;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1695c2d66a8abb93486ad2fd7df4505b519215a9fe905069e050c76de238feaedf767ddb1cbe26ab46bfa4fed6c6511685154e2616e8260218b9612b247bbb1d57fc3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c491127848f25d72f3c749ba165312d5f22c38e61bceaf0ae83456e6dee19e41a1c9d25460e54905855222916d0f7999b032fb80c79fc38ffc7d519ee120bd22ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a8fbd1d4125fa0d74d552397b46d6210d06dbe875be6485b2278fe737b28315a244ab3a6d00e476f3c39d2763c12b727440c1de4140c0ae50048cd86ea5fee3a611b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18215d133b014a9a8fda155b8835c978f52b7080c503e8ef5b0b12ba4f9ee94e1d5dbfe3b5267ad995edb0201d9c0dffb6fd9e3e3f35e2d5053fc6aec3b804f0fcaf0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ebf2e58309b90befcab79afebc2f62c99feccbee9322bea1da627cc4a08cd620c39b74d4e18e3b63274812ed104c6d8b959768529de80ad59d14431a116ebc0c0ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d114bc244cd0cf0783482526c732a5cf33408188870ffa13b7e6d180c9f24ffba62124872be9de0946ad9f9878ae60e5df1ee007d763ba8a8c7ca2fd974ee0177d51;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4bf442559cca64f3267d589a3d6a72d65023890a2ea02ca82451d7216d4aeacc9757c587166fdbe5b4e3d194c5d999419902256995e2b0606c20d0a364cef3f00685;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4546a147dd8f18e240947a73e16201697262f2883d456ce7618595758e76727ffb36955ba03a11df99dc377d84b1bf44b1199d82f43bc075a587aa195bb903827168;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a691a39bb3be1e88b550dcd5ed2e6e859ed03fa7b8fc542d5b40cfe9849d9ed961f92e19c01e486d559540619c164c0bd9b7611d19dfdb0fda1dc2e267dfb83146a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1470ab286e894b3036767ccfc0980edbb0bba562b60b4f8f5f9ecd0e7305bad4d113ca1105d46bc3d3dea02392912523c48dd58659d7298310d0c96159bbf9e266039;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc42aef49282d8abc0ab2409598b7c99093e113bdef5f107a5c77d768094b054283cc67ca78ed415d9b2ff49fc102a71250ffffd7e9cfb655eb7a1fe1e046f86d1cbd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a02ab7751c181f4564ebd18f6fc85f867ebec17ed598800c9a58bb6bbc01fb63a7acfa9ee6ca9fa13f526b0453760e666c59d528af62e92a82cee8af75abbc0bf7ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h58166df2be15e530a586cb9f3f7d101a92b1eaa799dc8c900584fdf8cab59851ed209601aefba055e3444b74b7b60a06935e9c881419dc9c966d35c526e86f57d597;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14de099aa603e73cb8ed255736e4077931be97a7cb4e77b167a7705807bf0219c7184b702701f932fb968104c74f6c7bd5311300f337175a645be5b55e9a3cd3d5884;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he863773f47d1ec2e7dc808ceb785ef96fb1bbe4384e6e4f064d45ea421aa3d0940a4652781b176c1c6ef623df413fc662668d87e17027506dab6e401900c8213bc88;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h82bc08224919a8ef6970b78c59b77e17d4ca9872a1ec44c587852b56c48089b94977c8a54111c4c68407c30fef2c524712ba9d262d42c7b027d40300dd2adde0d322;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa98eb7cb8b7816b3acf08088392567daf2887d8f51234c22591f9bd0ec93755a11236e5132c43afdcf96c0cdc1190c65231e5987e8133fad52748abd7a575b7689;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9acf29d82cafde8655e58c91d958d42e8dd1f5f2fb794c7e54a42477a76094ad0e5cf584f484299d7c9a39016601b1da4dbc1e3e19efa19093dacb7a450acec5682a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha0ed852cd05635fca4d8227b959ff6129e64e0316d0d5f706aabbbbdcbf86510832b9b7d4adf170d252b069e43c978b17226cb619ce83538631d7ebe4d0dfe872df8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4b2f88f2863a8b22f68b0bb88c14104ac536335bdbfe7549b45932a22098619276eb65677828bc51248ab0c8a8014c8e1c7b34a335456569bd713a351d43c0e6d448;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b81a04bdda1568955da3ca87239dcf8e7664a37863a7466e4150887321a1c944d6195bbeabfa63c7c959bff53dd053e73fadb505a406bcc1da111ba8686b80b407d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d3163cb86e227932ac00340b66d0c6cee9bda3e7d8e450f020524b4102894900d9f203b51ae5cc59d3731557590dd8c5f6c7fbead5c55a30d061695ee57444984293;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h26f96d559d57aefefb1827976e789113a3975f92addbd2f6e0257dd899725cd9bf8a934c7928df00c0dbdd975011ff8eac66fad6be31df6e5c386b7e3a22b455d56a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a043f96d8cf16b2953576fb52ccfd4ca8ee0079581f7600fad9036bc4a3b3df82f79ad9d09a742afdf5eac64c70ee97d94c5e7112b6f6b18da10c338f5773a85f4f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h145ba2d2d4a45220b7fc52e87f324efb055baa90e0c6e4daab31c5efc2f795ee496ae3f23e9f35fd69aec84ecfb047ec5ae1d79c37cdf062f40e0577d97ae6238903a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e6b755925a5e2ca259631f1bc58b85d3018ad260fb7bd6acea22bbecd107bcdc9571df448d5752ebdef0ec784e0e3ecb8748b3249596bd81c35b35557febb56661f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10fc23515aea90cb4afee96a634feff836145d1fb0588f41a9c8694cd9231fab190d1cb5c762f77d199d02d1e31121267b093faa3ff13594be58ebf89c2fdcf1ce0d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91acce06c2c0666478f9d1e834574eb40f8b549e224fe1febd0cdaee68039724fe47d83288cd233a0029cc275b6778d2f140b5b2e9140cf091bdd73424f5ae3943d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190d4ae8a751659bc6bbf545aed06e5e458b652aa56b03e7fa28fce137926ae8c439a8a64ee42f8dbc6f06d25940758e941523239bcc4273e7ce696c72095d542ff95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10037bb1a76a36698023bcfd503650fc3c7276a1f1bf3ec3e291a0d9372481eddf800824fcf2f9e6f0c0d9ce49abc7d80ee6343154692d2f7f646016a13e07da7202b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c868109fd27e5f598dbea8a0582d2dbd622b2cd8d4919e1b3e00171c78fdd24fe46561813b12084be036240cd9b65a8bc3773386d0b137638fb0a3f6388cb4ef8b5b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14d61ab6474b27a092ab7ef51c6ff694fcf4b3ed81bd904ba132c147926fe74c8bf922ebc8576bda4f23571b8192ca9d3db77e036fc1e69a0c169176605839c3e9f0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbad383b56a838787a691ad744a40df6cb567ec9a2796045adcdd4aeb0b3d473c0d778cb4ca1299fcd45605e138c3be1df4c083cf618aeda39df03626e32dda3b1641;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b08985d840069cbab049f798373f94030a227b97f4b6ff01fb427882567baee51437c74c51efbef0e193a5f7eb07c76d33721db505e0419a34cf2c095278cfdb118d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbaf481d67a38ac76e4950c1a87bb725f9612154d6a0c89db9ed458fe1eaf6c67e60646531938ac21f13f6835785e6793ddd6f15df79501491fcf479847ec04b31a96;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3476f36071a31f887c6af8068045e1b85d73a0d8732beaa3550ac7c976260a4d8541633dfc8ce8d6801d3635ca3655fd5d0f237804e28f4160328d6dab77bf89c3b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12641f082c2cf2190afc813c0c549f9c39290c70ae107af484b2d02258539b64f6e775be728eb2cd9f70c235da844546a50aced2f10abae7ceb04e5cd924ab6eade1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6686ef8b64caeeeb23b028b4dcfce0f68b772cd7ed7e7e6627d1c5ba8a074d0937a9a413035203bbaab11f9599d85b97648b249293d5b3ca4104c0d7c36e3b47f63e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1326f79e4a9d2bdf85629eb0f821462b91d34fb827da3ea078d64e35147456e44f9272eb32507cb25bdb901a3a87e19676bae47a70c2dd5b0599c707aac087c56e77f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34e2bb744d580bc26229c4238f8eeab4a91be7acd5a4be48c83ff9cf034889d0c28bfd0d43b827cfd100e880b62947efe0cfeb3b9585804f6b697b2b4ef24a0f9531;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d466cddcfdc9f427a7f16c8881cb2304ebc08028ac08e3a1d2725f91ddeef72f047176193f7538d5d0f7123bd918f5d5e129d9abf318538f01099cc0138c89bb43e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96bc5274c6ae11827cb750a2cc69f1572376fc0ac1be6a2d88097dcf934a8df3fa50f9a13bbd4d027c860fe768f52e8fb0e45785028915450a8fefaf14e51cd8f40d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcde5807aee916d464d7a01f8b68d311095d2561a143b5dc6cf6854ff8e700504ea6050413b58357353c07440d23cc64648d564ae993d0c2d4b30fa98f6b5daf0f3be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h134ce69aabb20dbd8f0078dc3f99f9a87650f0f455a561155d461d38af45a639a050b192ac8abccecb3d52a644aa7654993d1387d459cafab7d9c48c3c0111f3b7ce7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190b4f6a60004e4cf1a3a24dc30bfb04433b2df8e5808e7c2ea21722d4bef25d1adbaf7105697d9ca815b3c597456b4b8539ced16193dc5c430308cc62238d4125788;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h177da21002d15a74fdd566ac0ab2ba32e463ff95f1b389d951f5ace949fe3ee2c14b54e1087e8481ba73aadea950df4459313049cb7ea38269c999d9723c271ceec75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he96ca42eb6393290c17475ad9a53635a95f86186a8201f8a53205f2a1978edfa6e596f52533182a41bfc72f71bd4781fbf4fe09247400ed7f58a0c3c72bab873cf17;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16bda55385728dd9282dff010ecf8518562a0b506174c96ed3ad0bbf933b3a4cbf3d8df61d5dd0282c370c46eba92d4c7845ca8add89e326301513625b45c5e0507f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e4949e5e1c1a52fe06a134c6cf0236449294aea6e3b86c88e435c005ffa40cab3f23916050c7e7964ef40e810cc8b2a2b805987c8a868fe915c298adec505385629d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f72cb4e771e248f1d32dcaf0de58dd7ce9e39098e5bfc8dd6c14ae92b2b0b1b063fe2b6817bafc16b83ffc9a05d43727bb712fdb26985a57975aa3b4fe506c35dfd0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he82e91189dbb99aac28c959384b9af5eb77b88f6b820313a580077e769defbc00254d269ddd4fa52ecb89f874351b0385d1ae290c9916cfa99de68202f3923aec900;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1376d995fbaf231c7cedfb5461f5d0d0c87f000c45f17d707f7ad983bff36504d60eb513ad46b10826419f1530be4070e1ff6f691ebac459766ebaf414c6c1ef9a88e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a22718b5c7434e2b0e75eb77d6fa12fd64efa3560c4d1499758802354a0e0a66859c20a0e6bc7a6a35105c2c77e6287230950abec15725b2f61a46644722f1a96d49;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4583338e00129d748c129e8d2dfd889c1a76219a53a60e4374bb0448ad9aab35508c6d67de5a6624fe9fb5299f6ff68b7ac0155012bd76b32c1fa35b58a64f7d7722;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfd612546336bcd90367c440f190e958e927a84f6c3335df4917b1be312a52998a01c800061f3c4c6aa274b7569d209b12b1d2328d9bbdd240c674c7f28093c75ca9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a506ad3c96cb127f3853bf757d823bc253e9a87c97dabf9802cfcab78b950df3696155e3782f02c4d2be0ff5dc2c7ffecad42f5e6b382dfea9c2e533483d52895c34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbdbeb2b5f16d6cea95dc4971e2827e23dd998564e11f7df64ca27241731de0adc3740e0e6ba8c2f428939ffe0fcf4e1b370df9060512e97bd8ce90561df29c9b453c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f5b93212c9c95ce23003f6a6a76c182fff4d05a4716d60157d9d4c20c056fcad19010a51cdc791c2e6f2046d19341a516a243b3736d935b528734cecc96d18ed8a55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h62d070fea0837ebd42c34fdedffb617bd9e8a070d46d51116ecc7de61d23df5e9c62d2b0790dff3a858a9440b7f512e77c3ab3d724bcf0176cadb9f4d0c1aaa94d99;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf74ec4f22d77231ab00a9fe888704136d41c431a1e38773fe15991ac7928fa4ff3c77c76584be5eb7605ef3a6a0bb84c2d48eb471607cdbcdc5a63d6e8b17cf959a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d40d1bd4ea45ec6ed544725a32d72bd4433a0d35c8b261ecaa70df5dc607b164f032191a08464f50ac6c6d44538b5708c3abebc71a89c09a41c3472d7078377b91e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb02e573450852aae2c915fc1db4740765eb42c9fd8d0d1c8dacd31bc1c167aca0da90ab550815c4c3f4168f6bfc2df87f73582dad6086a66db3ce9afccd8dacc74f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h759477bcfa3b7b1a15279e5106bdd56ddc844599a2dd4ba51edbc7508b1ffd4aeb88892f5190a4ade2545bc50f91035f35f6eaed46ef5ac00589f2edbfc39639d61c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18714445be5958962e8179253b2a66d6a00f854bcedb1bac765951fc8f55f1036ffbe7573527f2ad3c1e431b76aae11bab7cc73337ad850ad3edf769cddc42964f51;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1899fe8ded0323c60ea3e11627acab76967b5a7e10e5c11ed10f8986599886bb6d622759b8744e4a63899d07352c3d0568141575bdaaf48a2ac9372e70fbec11fdc53;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1457c125ec0565ba674b9786d8d1f96114ba5b75e3498c8e0055bfb02c123ddab21f4262552a7ca7645702ebc9d34ec078e62e2ade9979311d5739aa74307c19e2c32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1edc9ef4be51c900acff1473c7870f86e4758bc639e0473a79ae58f4b23d03992970c652e424c833d4f44d31c88d163236f5f5299c5d6bfcce0500dde761d9f718dd7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc793711a94cb965e5c352a4602c3715f79436f804d8a898c421a7b0a0aa8e21dad672ab1eca8e71edb12e2ab1ff90dfefec4f8a68169534df56a425079b70938547e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66e38448b983d5320a92ff9a43334a28072b6f9f991fce796e0eacf1839f684397938fa1253e78925fa9ad93281c60375ffe60987d961bb0fc3c3b40d31d04c65951;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hff7c5ff0535c32a94698302e42300b087203db6f2a7365ffcc73e1784e10adc793bcb7203455b7eab08f7ce594bb7e31095b3187b0038f0a569b7541fb852a4dffc3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha85ff6bedb3813c89a289ebf4719d3c6bd5c828e96dd7c6f927f87b08e926b4d9f21f3ca9a57196c703e688ea67c98fd00e77c9696db7064e7a999176c347734f8eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a28e977e5ce85158b58846059a191addc8878155975e0841bd48c28cdf4650292d8c950cb15826ea34bd1c80304a48c084ef4319ae49af61d85b87f5e5c7006b00e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18805fd9cc482e62639b5a4123a51ffe1ea5488d1f8e3a2f192a83dee66b62d04f156d91e16f839f8ac7a0a2d663ad2c9a86cf475b5918b895eefd0601d1731e6bcc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf12aaf3f795759d8b8f7da930e360d9bc5eb7b5257ef0134028ac1543adf8380e28fe6a6fd671144fa7a74bacb5e95769bd39a37e68a57bf0842bdb31012fd55fdf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1be94fa8e5a5f16feba1e210e84c04621dd69588d5745362e8bb347be8bfbfd6857bd9f62fde71ecb2fdeaca5472e86a6251867bcf714f120c66d61a8acdc426bd77a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c64dcc28bb3c374c898631a16dc3a57e6090693b7a219e9f1d58ca634f6ac619be61691f9a51902d4215b08baae10581d499beefca7c394a1131d0b29666814e233;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5a801b7067db6fdef8b57648e14cafd3754af37469cb02a0f91bb3d135a3299fc921620416a40b48d9b952f3ef6bcde970f08aaa09bd861c50a24893d0bebcc20747;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198b997534161b9e351cf16ad88315e2281b86e81fe482e348bdbe2acb6b7daa6a11fe47106ddc16eeb1a0e9efca2004a535426ca2e713bdeb50f1e2ec1fd4d254a15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc023709f5a59509e0605c546e9577073207a593fa559d2bf77e5b688b13c27cc005d20b3efcf752ada4552e8dadc58a046b0aece6baffabc00b3735ebbb681333f4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aeec856823751c17e7d1c70c62ac794d45ffdf13bcbb1c70bddbe2bcfc2130fa1d55fd5decb950346813ba04ee54f887afd5261795f632a2203fae24d9ad5aa56ac3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17dfb45aace7bff14985e59b228539a02d1d2cd16e50747a7a02f23c08327c00a4a4a3896cb107969e9d933e7b2dddddfaf2d9731e5ecd7af753c3e5f358654c97532;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf7504f6b206bae945461abebd09a459766bdf300e82d437ad41c7c0fd062be503111c1f89e48dc71a6567a426a312019c50f57ddfad45a81c803293614f1e2936954;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c16977c8670802561e8f8a181f6af889308738281f9aee7663feac56be8c646398dc8cd91a8a13997c48c77d4c1ffdfbd71d11b6f5396f2a4107526e4347371eaa70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b298584b9740b604e013b57800a5c5640640b3423bc5ef8fd7baa1e90ab08063871937d6576f3bc88232e4d18a01549033f2c4a6bd5290749c6876a7e0e0dd1bcdc6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heecc4ad473c74af120914b8a6e45e606ba0292b3154cd4137653c950f734fe4b80d4306be87b423694735e39404ddbddd8f7f90dcfe8fee683e2f0ac00dbb9e1d855;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb7f519cf94b1ffffe1381fc58b67d050cabf14e4fbaf47023ca9bfaa261539241746ed3bedbef7f564e4d42e8ea1c6adb9ceb1a740e1d8ea3eb2d41d1f466774a9f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad9f81b57492e13ae14d2079b10b4fc420f30c31da4aeffb9296211c63a9b23b0cea2492a05f60e71eeaab33ccb9a8df63ea2b23633a8a562babc942c3804ee590ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he307a9a9d9710cc300d9784e79fc2f82955596a225449d45ddd02a95cbb27462cd5edc965ec468534cac9fef9c8ee45a026b1ddfe348d03a1b7a5d9a918e53f94887;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165ab0fd0b0427191a8919a884057cd194146105cffa8f6d1d063b908d1ad7f26ef0065e47982dac641ab6e21aeb6e353a30b0ad85d2938e05a71489fed68e663aad6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb201f6d909ad37464a058ad7a6e66dc16ffc8594385f59b8bdac4f5c2fe2aadc9bbdfe13db6909ddfdf5fd766a3921d695caa0a941854edc242273cbf80fb35fa114;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ddab6667882b16ad381860b95e6ced6e6bd34d549d65a6f256fd74d4d630dcf4448d9559a360810dc43b17f31cb304ce0739e60ada93d1334824786406192087091;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bd7a90b71e749ebc1378bcbd8226a18d933b90c847c13f6bffa7299c6b8371bc212cfb4112899644f17f463626efb41675620441de3741f95a3c4805d71a05587269;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a6d2413778a47bfefb3c8a34232ebb72816c133ca78a833a71cf08518a14684734616f8d19c7440efadac7f0c7de05946e513c3ea4c5a61ec3ec13cd06ecb4362b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he893b8506cb8c320457980c60e0683fd01f0038f6e0acabdbc8d8a73b1beec4ae508dbe34c0aebfb95c162b16c9d5905d8ec9803b1f720c850d1f9377b4b415b9f36;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2d138661d4dd508527bd6a04285fb2c5190163be857b1e3b6adbb98bd7eb8af9b77a9473dc9be691a0d85f2d20f4ab7d0b68505adaadf9121b2fc6a78204b981e91c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53bdb5c86e220cb18d58171134a30339ff359bd1e40d7839f9a1385a2702c5c5cb9c76baaa73680384d8c999cb28b8170c091de9956a3a6732aa3f2cec9823525112;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed6734a39a9388b187ac5cf8e10c0f5ceb232e136238361bf1c582e3b8ecfd4205dbb7c060ae79ae107e48580907ce4631aebe61a55bb86146eab25cd806613f11c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h41fa41ba66c6c7d8c8397ceee70a9e065b5468c29c546ee2bace31c4de45defd5b797331f585535ca2c28f70fd7d2f222f70ec018c582ee90257acccd911fecba414;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h436120aadac79fd4b381f85adcaf05b008bcc4102379fda844d003cc4ad8a7224673eb976c438d6b6fbf6614b6c2bd510f2aa8d483b6dc482a6f9177edbaf3be21b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13acedfa332a4c51300273fd9132d329ad352507285639bd841c3261cd4556217b388ccb062879cc5577d3a3021bd4bed7641c84611ecf617bd643238cb1752eb9473;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h173ed44cb57a269ba2e200249d516e66b4ab6c20b0a80cc540b2287bf165224031be4a1f8f0681e29d3f889d7919323ec4fe1de67b40e22233449d7e51fa0e42715dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1023ffbf7f2737aaeb5807da7c785c6a69bfc632c034ef9b7eb6e65b8970aeb7984f41bf15d41fec91b1ba2e14c838e59d611be257e4375cd9e1ffc2c148165004d51;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h30d3676ee45e6fe189581e3e1ceafc5fe65ab1b2104432b71b4dbe48ab7dfd6737e4bf346da126fe1ec18181e136ccc85cc0d45296841ca45932749769dda24283ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h20b004ca9808570472fc2c523451acbac24099b262af5d069676542241e3f7a7441071a2b8615048e7511569b4e835a3d6f82ad5badcca75cc0100b00359267a8b4f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h109a7cd463a82745e23911a2bc8526c9213e0e05bdec4e930329cd875faca93b8305efa15456f5e3ffaf4d9591ed6df06971d2ae94102eb27ae3ce15f0ca224b69d07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h626469ed4498bea4d955dec2ff65a2ee07201119cf525e5cc0baec6fa9dacf064110696b1c39dbaa758971bc6bcf3ef65b5a945d07bbd2773fd7215a9f6013d7bc27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138554d7133fc336e3192d8e8969cf0d9e91a51bb4a0939eb98abf2efa636ce76032aa6910ce7102885c2c27b87b1b859861a49faa8c055433158acc6dddc0f189857;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h100dc2950818c94d0a1f2fbf92f3c7c26f1425a8e202c6249c1f1b507ca20107c223e0cf24e850554f55a21933b75ab87d169ab69bb8c4104098f614e040341981fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118534c686cd0db064092eb1d28652ae422f840613541f7be78d4d8876ae7b1e8fcf417c182fb37548ba33c112fe7acaef167a6329212967aefe130d5bc011c8ef619;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdda1466d20c33d65d83b8a39ff11ef3c828c1aec80d886f7db97def5239299d3742e6103003bc07f170d43739609fca87f10cb43d58ce43b68d030118e2ce22461ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a063accf6b89108db0e5488c8bb959c312a9494ead0231f856bd1b8bdb7513ffc006eb7f3c6b0c09b96b624b070e33d60c70f759ff74d0698395ce315338d6378ef9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17b2f7073e0edef9ff5270011ea046156c6bf906388388c831b5df46da17ab679703ebfc54e2e7a163d1199725728d2c018027570c5c94db210f8500af7f0e6609542;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19983138297240f9b4d3d1109aa882f4ef64ac0b1468766f8776c767b7baf235ea9ffd775704554e75eb63c067abcc5f7247ea59a3c64725f7bae5dd6aaad3e00f1fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h112e1821b168d895cead32a63b59a1d64e244d2a3aa0a5db570d509ce92bb934fa9d6d4387d3827960f0daba6dc13f273fa3caee57e619fadac9a3888fb9cc8e7e80c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14fbfca5e73bef7cb69ababd1029e99179e06ff16bb445d9551bb065c22450ae74c424b9973ae5b2e0f8c8bac55d8c05147752c835160fcd3b721034262240a11fdb4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1066fd24539a6d54db8761f585c3d2d022af00f2ec7a4153871c46a5a7628cedb4befebf94170d0729ba1055ce4ad36f2b19c95c63aef0278a9de1f0e9281e791584a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1664c981769975f06003efc7ea07c718b6fd1e3c5878d0bd096e8265f18ce4ab8cc28950cd7bb054c01ddde74b07f88fdbcffbc8136b56358d0d26b35dd1d35ce057c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h985ed2c3ce36f373c6c8f803af682b670856d35e1b1558319a0f1f2b3368a0b9703ce5e51dd979cf8680ef18059bd80140d321164a39512b4e11893451c74fb9145e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14bd80de1fb94994f1e8cf3fea15768e7763aa06458c9eab31e2dbaebf3e667e0a5a299666654888a4757420a5cba0c4ebbb3b9234857666b83d8731cae5a1e863b3a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h116070c24fd8b98aaa603ec683ed366f26a11b7b5001654cf48709c24f5992eb18b7a8da55d15eed4c45f249705bf2c30ed0cbfc2aa67bb17512b9eb71628a9125568;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5583b24fd51d1afd464d0061511ba66b1cb8ec8a160cab136cb467af7c294f337a89a6c63fb7e7028e5f4a47596549c90dff0d75b2035369b91dd282004740b9408d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5be06759825c1dc701df1512bb86864b3f1170680223e97ba841a0943bc83800e3df782262f42c99b0d83972cd4ef3b143162d63ef0c5b097ab0ade39dbe7f3c2ace;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h122deb0b1ce9ea8560626bb8a20922194ff585be96e0dcb61d9278b92d72976e3d4d47dc21dd0f328687797aba526f0caadd4222d1d0c07d3999c498b4d66768465e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd34e7d2fbe8e38e7653a38f724301d598bd8e5e451f5b277821c2c26af939c0aff98a46e03ffeba1734060a4a02767fa343c3956d640af1d9760554e18d0928f67d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c26e3321925ae62637b37466759391b4fed811cf5409d20d269f1a990c7eea63a5efa57c5425279f8efcbb217d5c3e86727d0d5cff5ed84a8014a8e519612e0c67de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h629f6d5760aa857799c4f6e8ce70930cdb7a92241c0ea0d250f33b38cf0e4ebae166d05059566dcfa764711e71daa5828763e3cec964d3c30d149f9ca66db293ca62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e5536c730f5a5a09f09f95a015ab8e1f7dacf68bbf06fe14e8d720fdd1ec036db2ec7ac26fab618f38b5d6ad2a227ba07b7e3a02114a25dd45795c62c7f08fed85f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10879057ab0d7a0df88a35d244e0132a0f3247d6c015c96393fea62d8b00d1e3ccc30cf56797493555817ea870bc2a123503fb2ee9107b9140d45be400b2cdc92d4a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h30a233b1ad4fdae9e2dcaf1300b84029288f8f7855e1f6d40e171499cc4f2124eeb08a1b278ab761afdcf9e610ecb3c1e8dfce700d2c2d957113d461ae60acb4e377;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e7007e15e3f893afa03e92d9e9c918cf65fdb68b59145c89970dfe5a996f43fe5b7aa0a34eba45f2dbb245526618984459ef895d087c21880163b981bb2456ada6a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb273905409aee07a91a77c5e8c95e4ba19f29caf181e5a26796400fcd6c13bf854b45ac4c7addcdedb44dc5b61214c712420a5619a8f2dc31882865bff303a11013;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48e26f5242f46399c0398d5c9eba92801fa0b0c7213a4f52a0894d581dbd1dfc70be9af5dfa00f7f27d6c81068290b4896d52e597dc8f5ed277a966003ff662ba7cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had64aaa51652ecbfafa4986de31891e188455761a7fad2a66c29e26181db67aabe6258361b3238ea041d35b34ec61a3f6a8a781b199b42a7a0dae62ab56674ba4e00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2bdbe62eb64852e61988c8d4478ec7e80b0d749b0eb115507a9484c6b1b16fa6eeaecfb652de3a8d4e93d5f94fabd52d03b69ce1e30c3ac0bac932076022503244bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1980afa82f8eaeb650cc24aafa1cd16ab346604571887c6e46b2ba09dd5de78fb32772e3372cc3c85326280dbdb7f6f203006c9646e21bd3338c7c6b55e14fdbb00ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1488ce69becbe78ac522ca19239cddc882b43ee80c0dfb1726a80ccff3948d276cd4d1a25a21d416669a4e4d98af148d48776544c2abd3f1e8f1ef35866d2faef1944;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19e85d6822ec4d2907cc3766164dce5bd0970032a21337391b6d32965cbe59a28f491be886aceb6a74d3efabd7655521797dd8f4d87fb2019e1653ebab7e3f3e4ca04;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66135fcd2784670fadc2b731a654125fd2ed03fc438a929cc8a53a3918ea8b93b2f077b8557f8c230e1443337ede7c13e233d664abc11f625de96fdd9028ac138acf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h447eb0e986fab23ed44616a13de493a469f83bc6bfb8de0f7a26dcf61f710ae4d9ceeac5ff34c40e132e05e7aa119fb4396a7dff4a3fd0c62dd32dc0d8658655cf0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha1ba0845d8bbd19f3f998acfbf6c8ac2c4b864eea3609ca336dda609001dc69796b9b5e38cf2567c0e072bae95374912d8e474b4c4b7f706d9e1035332ae9bd5b24e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e536d84fc22c29b3dfbd72577d2b6a7b966de004bcb4d1f06d40fdddac3686751a0f38ea519d48715bfc56ee4a56f785527226fed851a1198a111d09aeb5b0f83e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he089991d5022473ca8a57fc8204abd8e1f9e0570c4e656ae152776f895da26e7523e6b55803d123def7a28ce19511da7cecc4126d279619ebc3e2fc06b7af455166a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8dbf029824c50101f2cb4ca93918059b8b6601d826067a92ad42d834f8dfb2601b064a7ca9c857700b8330bf495dd9c21cf5070e676e8e6f669be81d08b5a644907c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a21517579aac74fb1b66e9337b5abafff94aff201b2121b1133f865b041c2e3fe2e4c1c5e933018cc4100365ee0873221ed08efccc3c2d515230709bf97c7d7228f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h56db40dd4dbdfe8824bb79ebd92156ca204b853a4c32887dc6eff7337cde4aac7464aa2caad273c74942dc1ea1a4a5d2b0f88df7571f6d7ff91be3196802b8f8be62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f4aa42c7ff0daae6523c5b32161097ac5648355fcf1d8530b0af17958b576883e85ddfd8486ac86d94f272897ec34ceb14af67d38f20768ed70a5bf9d284a5823e7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfb499243a2bf76ebd88f1afa2c0942f7a14ef95596c271a2bf6faf907263951996e5c8626832381556c7221691f736581d9a5ec317ee52c874cc0a2d5f197f5a433;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf120cf239855256cd122a45e2f1ae1c5739d76607100901aad9631e835df3c333320cd67084645d2631ab8f95a05f37bbbbdff3d02af8aeb86db1ede2c876d41849b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f5555b7098bab65af3ec495f1032993bcd330619683e53c861ead7ad2b73b7e0702651fca2ec50f3edf43d25bf244a33f70fbfbf9c38920c4d879a679cdcbf4be52b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hff9e6992e8611d7a6b0e060bb68e8333c965ff0703e3c25f4bbc81f75d72038bb83d1c4184785ca7ca40567815afb6926da427f7a81251802e8a57753a9c77db06ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha4b1cf70f39b815ffa89ef2211ab9efd61a25124f1fae3c556f47a07b90d9a17d061d30358802b815d46a76ccbd52c746acbee15ff1138ef96c4670bdd2423f24eb2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b14020a4070158664ed80d86c89135e7d5e411ce74b6078380845772c53c638e10449e2a0445d5c6128f8c692151709896fba67d7b2fe0d8bfa1d1530739adceddcf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h51c2769fd2b86aebb93f08852aeb3842b1d79e47ba4ab5e06799f3df406220209ae9e50fdb2c8f202acf84fcb68c3238769b70605025c0ea9eded3b8bf531e7269fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha7640f53bc4f8ce92545c73b6cad28b4139becdb9e1c9a8a559a079e6b73e87c54fbf188951383119118b8e7c183ec3c68c242945ab8aed238070ecbbfcc55c15028;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc3bff5633ea55f285e917e6a3333076eef881bc6a3485034219088fd5380b17efacafaee27aa99d0ec3674e0da0b88361339e097881c1ef3df9b4545d3adfc32ff8c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c94590a653633f4edd1bbec0e2f368add11f015df25eb30aa6ff1af29c6d8288b16e78f53d9303bca312fdd65cbd30143788f41e1e631ab5b98cfa4cbd6a0dc19f0a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19e1a6a694aa01b7850ee415578908a6eed60bae546ae9ffd92c5874ef3993c6e8a3cd1c39b0277a83a1dc633c2d0b16a749e0debbe142e2049faeddac755e7ce0616;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h181d5ff944bbc8fcbd067f5289320791e7c103c941fbfef15857859ab04a3a272ac51070100b9c7118a89500a9899c4039bfaf0641ec147910f65e531ae663379ed90;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12976073869c02faed63a4182d681449a92a4cb65e530cbcfb49fcbf2a97c9b88ce14ae55bdf65ea6c42eee10b4c673e172bf5787aa23163f36ab7667c67f8749e9d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9b2d6ecd2d3be821f30e0721a95dc26bd93fc8c05a55576ca1cb680b1fa60f397c0f50a46cabea738774c3f777aa8098cbc530393b0e826e044eedc185d3ca0ca1e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b72ef071a1ac3c9a0fcc3e195659393c794579500fcb920eb92f078c637a06ca3f48669f72a5961a91f291764482d4cd0b9d52c84166693efa14434c2db1525244de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had357411f243568a66b3e012e14735ec57e53f68822798e84714df976b4497d2736ff9102ed66834d220334e893f1458df848d9a7fe140684d6482c648696359d496;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13e16a1c4b2f2f21076a79b3514fcbbec9bc76887009639e2c94ac5bd8aa6c44f2ef3d3639117e62bd63358ac4655ae7f001622d2894b7320dcbdf317e5baaf1a311;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14125a221fec0051bb997002b6341350de534502eb45dc2288b699aa407b57293e03420482f9f9a8254d54933a7b1a38771caf308c2946bea55028ad23e062f2dd10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aaafa6e6d492f6853598df3d7a266d49ea91fe31f0bc49d92d537ebb4e1b5f007170eb8d614b5079e48e26edb2c43eb69ecac3731f48677f534b4e0a2c21ea5066cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e9d97472f071f0599c7d63fd220768cfb34008f741435a66df6307f44c7d9900b93b9ee45dd2ca2f41c323fa1f659b39d9f6be6c9b9f032df6f77a34b88cdb9ff09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f1b365f03e30277f271d2a527db055ba0eacc11ca6fa46ba5aa5b21b23cac46991a6657d26370791b1f71b427eb10dbeedbd092597b64f2f5d9a1a8ac53285d6e138;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd882c1f958e1c91571b35aada4e3f3d5100d94fc9f47f0d72ac01d8b550e0b170316390ff33ae2086b65a9e773edcbb548989ff150aaa2db0ba23c99b5a9a2269f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133758c46745a99b97d8a494b2376196e5e8b3f76974ce709c7517fc7351f499d84b04201a3cdf36690a8092625d69e66762d3e8e090f542e46ce4429a6a42579f201;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149dd7779b6a3c2b435f20979633549941a4de9e6545970e301195923b76869f42b1c113de9da121878663246f5326d313d0a0cc1b08f25ea0c3c404b064f21c456e7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b02e76644d0b1f38e42ee297e838cdee1198ba9cacee1999c1316221511506b3deefd9ee79e3c2d515dc0d51065a88806dc8cc512f64345f3b7b89f3384ba8f5a96b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb522476eef847bfb0d0a3a0017c1c84a2a42363eb63eb1b6a54dc1dfb17c6f838c8dff2002c2d2dd6dcfaa7e73148e5e6f62a445ba4900c60d0d294e2e0b5e35b4e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h95558918e155379bbe5dc874db1960963741cd7460acb6d8ae7e34717a64e7199852f4b82fa2df98f784371c516e2e8f9b4b92213de4aa4a1268c2522bffb95870c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19b3e96b823707617077669d527c24ad72e779a741f6e8a3688954c4e8dee0e9568d747446840890c9b8ef87c84d39e5c778b28c4c8f1ab6c9d904d65623c3ec53bc6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h384fcc54caf7195954921aef1d8cfa466b11bc18798914441f98b008d249179d992c2066cbf125a8580f09a1e74676a3f409d02e7959596be017a13234425aab0035;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1218be4fa484a39fadd6dc27c2443708711702f1bd2661040c138ef5bb98a3d71263835aad10c02a4c2ddc372e0a371cc1193f9a332fb2725ddc2afdcdcda31fd7f29;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h179242e876fe5a8f5ddae6fbe2f0e5420aa7c496b6400492029fbf44a1bd344abef3296992887f91db392366903ee54bfb5bba6d8408fdefe9b81904421b9756a543b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d629690b11a86a2c76ca7af4ef7a96041b29166fd50a08f549b4f902d4cca3743d5e01e20687252ec31e69c6c392c0661afada12cd5304fff3e47560c4bd22a9677;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2bf81d4f5683b122b4dd18508c62e8ffbef77cfeedda8280deea9e041994d7dc88f021f36d60c33fb5faf96f5a67cf6816ef899338e38a8d99dea3b4c64e994f1c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ff897be6bc1c479e56c820b23a402cf5b8a34c56e437f14dab9733ebfa031793240659efe2f514ad8a0ddb89e1f29def6bb0ad6920c861d0bde5b8dcd8059a5d976;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97065141c99b254428f6b38b7cb4b6982840a047a81addf7fd4da46b1df40fa62af6d54a0f58f07bbd567a4a19174038e6da95a3bc7412a746100fa582176a0c27bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48ee09817f21b4e8cb5d1f0f8cc4a1040865ecd63fcd4832f37d926246874731f92b0498a6af2439dd783d54664e3aa15f63d3f3864aca8e9030caab04c41a1a970f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha1ff518f418b88a804c50303d5844484002377cd3284a929d8506d27afc37786fce64c2eb5ea194a5e5baa48fe5269ad0d0dc6d799b627754f7f3cde54a96488b64e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1216fbb8ec3ed9c532c93f4b44fca3375e5f77b3f60773a371a1c1d3556cbb939d295a19ca2b190f568d54ca086c7b0022e046462ea0cf882cad0e75ad1b200429718;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71d4658af0e977b089d56dee02fee038004348fc8a94e7a26380272269f2f6aba3b1a73561ab014d40a7e5d1d236bb884757ec23ed7b4889074b23d7e10ce746c91b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12764c0d5abc5edd0e8da29ebe1d23c45cea084f049cbe6f9f25c61fc080d5b07b8fe2142ca8c00515eed1d5ef5813c5a4dc7ccdaf6dc1902c3b4ab521e98b185c922;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h76ea49bf91ea3c974a698ea860db351cad8dc20a16d83de1ef0c2ff8623097f73071ab1720be37fc209a5fd9cb00c9e03ec7403071d63d35bc1b1d0b026ee60c0011;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h173ec28e6c9086389ccd663dd75aad1ba4ddfff1b0790b57ddec6ade854cc751f93f40257476fd9745f4ed323d7a13bd114bd5d92596e4bd7517ef6874ed45ab3ab8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h148d55aee4741b736e653ebf10d072ce88b42b13c040aa0997c2a948bfa279200598cc9f58f674806d74df17c98703551b6a7ed8773510016e0915ffcd1d999007da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ee1914f0068718aee222a56239eef18be98d690cb5743cb207dfa065936099d8bc64ece5859add1f9fe0f3876d4ec5083aff5e8dc35551c02b736cc7a0a6b22c838d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19dc9bdcf4913cc3156bf7904a535a482007e11b585775119bec36dc8c0c461333f300f8f9cff4d475e4064d9fd060e378411a20ef2775983c18979323652f1a35fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ce785267fb7e61a1674412d66496f98ca7960da960785c8878314a2bba50ba84b879c66aed1adf4fea55200cce90407218e77eabfa5865700324fbc3cc4d453fa73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h32b60fb7b826caa7cb569e27fad9b996624a186acdae50214f7f24251ddbcd8f6ef5ac652a477b0eb140f020dd6d22e0846d6d4773a966370c374c4163c094f758bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79f8229f2b91d2612b19808ad955be552b6076503eef32e13dd71c52dd01ed4ec6713abd304305ddb8f5497dc5cb71074d2c1c73e47c765a9c67ea6e76dda43cb502;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h163cf57f3533ce4a3d58c422502e213371363b2fb0fa0399458fbd6b83fc2f2817e2a32113e2bae38613ac92e5e94d4d3e9f71e83e5fef5d5966400c3421129d3b3be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h421e425634c522f5e7c2b9655455903efc0f81dd975ad7a63f23290023b8ba65326533ace651d952e401b023fa7ed71316561eb0721a1378953af65d0704af550b77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3a79a92ceee11b2f655e04ffd8ba739f01dc876433127462a1eba1e01af05171db6c90341c42c52b0871579669f33716647f87c2d0935bdeee664c5ae7e20186e5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89651f0e8f5a3a5848a9f7dc43cba19555951c01fbc74d036aa9b39ed72603791d1aa1e7423d9a57aae81673cad87607d886cc6296874044b19b3a8dc7056cb68c3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8c1ad43d72fbe598049a05b0bcf401db0f188098a01ffeb24decc4d0b9ca4b8178f68d13dd1ae175a74493f6c95dafa501676db17a351ce88435199828f9b793f41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16eac2f9d4e4949b6c1d45061e11c03f6f25416e86535de7ec1555d4bced24808df5523667ef5b63654d23cc5621ef120600e5f20a71b37a0443d63949a9cf441b73c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h25ddf71e6e48b047107f426c232cea6b655ca72211c14c3e24aaa0339d7a86284fec8f7d4d4f6b3d7afc506dd1f09d9b5f9d4fbd995e694b99a0d670769207f5159f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc691a9603f55ff42e2c02a7b2e528b87ca87bcc1e34966f87245aad6808849d83f330e95c173f1115acf127f829b8635b63ae6edc04548c20b4bedbb35428712f352;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd15fa2ce04d7fed3712aa64a0a2db606ca65b9fa6f6960d7e1d37a29a0ca79c0f8fa85c3a7e033ddc6d897509ce1aec33755c1c9dea6da533381d7d70c200e30b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ed7ac93b2350df9c4fbf75d2d28ed050b711929527461abda4056eea1e33ae01f4751e7122be631864493857856394d26cfc7810b476bb8ff1ab90457eb2fba85bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb9a9a581d47bc0110d7fcdd9cb23fb451844fd81875e7d96e2ba605fb256b5b1bbb9793705bbdbd8f2ed053b7a7f46296dd868a0054ea17d1d772303a52a42bfccc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14869ef16c006e36accdd65bde01a2c41ea5f9f6d365276a63b963492af065571be6141bd626b6db4c47f1fc7c7089172319bc36eed6e98fa27ac94a6b7cafece9792;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18851a865fa6f6cf3ebc42c3016fbfb6853e386082beea426f1a890f3bd437fd0274533792e9a67b8dab9d268d52197b9237f69344078d3817538290c075871c6ab8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c151b3121f78143431d144257f07624ae22a2a2d90d6816dadf370d0f4ccd12349c1231fe9bca6c5c13fd13f79aeddea833d2d746572c42fe80d4b39e65656170eba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1280877ea7c6e1e4d4439e8a68209a29a69256863793028515cbca5d424ec658e4732dec521da5626e4ec86f171ee96ec26db67bc5525ce8a7eabb433fc91b7d76727;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc452538f89d0306999bb6a90f854263b0a3b93d88e631c6cad5aabaf5c86dfaf9a08b43361d91092b0b39285efb736981b1af8fcd903483e672cbc5b72e293405b2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19679f75f2714c76e49537b2d2cbde9f58f312d229cfe6325c9f7fce106d9a67f4a1c4b3a78e4ad0d5fd381a796c06142ce9f90564acb1c0b2bbb04f48b30f7bfa3f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h107a0458404f65ca4be3392f7b7b9af472294de8274e50e96367dad3112e4b9443f54a9f0b8483ee80d4943516b0a6d6fb026208dc72275515d99b9fec4f21886d595;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h30cfb3f8df50ed8f6a8744e832852573a0b743ddc6309c837929a7f21fbfbc3c827f46038af9991732ad67ac93b7231400508eec6ccfb66a0b874048bfea27d8e24c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8bbe5462acacc447e327a6dc7498f4592548aa9c3c48e1de7bec9724364d7d5c6b558b020219175b5fe260b80c0397eddd9fb7f1ded5062c091380680a1d25278157;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11bf294a3993ee0f8e77f5eb3c25ced8acd938705a01f425af2414b8c2bb95fd554990a32c5bf902d23dd53ecb5a413a7fc015d0773946f39ceb7fe561c0da7c485c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab1afe114527c1689efa6895cd78116e7837d1e8f42a427587f85d86248084ba68687a81ca812ba3af9f6f3adb8a658a716786cb86e763d7705bcde4f667afcfeaf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h85bfec3e9db2310a508b5f451fc74c54b32b4bd7a6adb3b4c4d588dfceb98afa3b98ada6cab944b43ee5bbcc60a6bc6be0cb4cdf1d5c643b86d32671afb3f973854b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13e1e303f1eff3dd930b8d9e1d49fce1f35517b0463aacc0b3fffb1535b33f9eb41e29e4f8ce3755e8234560042eccc50162d3ac14ddd8cc526cc95a435f652139924;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc541f726ae5cbc2ea10cc7a3dd3e3565f76fd5e3d4eaecc4d8d2aa41283b8d269c24211a59fb8c97adeb2f71d0de5203bc052229b5f8c75591922d334ccd05ae016;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a184248bd45c3a40450d2f9121cafb4c4d75186787f9a939f8db1a73e36e54e126e08c110e009cf20f03c75e04e971dfb5144266667dc08b9597ef4b92af1decbddc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139dd489ac6cdb33b71aefc44771eb8227f69dbfe10897cb887f85fc9cbfd032093bef65b9e94887a0a545538c6e02e46aaad5f73c1032838d24b8474cef713909bb3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a95f673f921dbe96708c4ecca0ab66aadb0db1da7418de34908f10432c9a8317ea3b33ed555821a0da8cd19fee381c7ecdeeaa51e5f120dfcad48775f016f297f23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h22bc020a93ec29769001fd87d96ca7e7a844fffe5256a1db2046bf288969ee41d386eb25dc10c0fd1f305f65c0de0eccd58c7b5a13596e03ee8348be9709381431e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1978ced9cc26aeccb673076ced28ae6c5f7638b4adca72196584bd467ec394a93f524caf83e025e03d9636b5ff1a0cdbd6bb46d0877a25d98c15a0a3052c9675feb42;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1093ccf7332680283d6a752e6b4cb630d8fa5af35fae715e6cf3f76942a1c2c332c5c856eea11c96a09c0275cb8eaf13f11d90c306afbb9b4631d355dd4dc0d62969f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1015bdd46ebb2be473a276c047946222ee063b5d212f7d40adc61956a906576e65a85070fc2e38c27b13bd3fc5c19e337389305f77e8a214da2f293fd469286ae6b83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd031c001eb8c08ba924dd43a4b767528ea193ea5cdf4ef3f07c138ee5e68c2b2d215a8c14c09d5975438f9c6393ed9bee68b13b5d8a60589a713989c489b160e450;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15fb59f1d484ec399e4cea339c3c2e4d805f5b34300ee53197c25de4110dd368c7dbc973fd6084cd4afa7913e97f9b4e400ef2c5a2b87a2fac4373468015374058316;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53e9829b6609251d679e6ff8749fa5b805123e96fda6bfdb43a2c18558f41f277dc0ef651ff9b091afd982eff56b2802eb2003869d5bd9bca1514ba997b40d8e3957;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e30d16fd848439afea4c8c5b58365f6c7c5470d8d441abe9384f49ceaccd1180f420553b6c53df529caba665e2ff9ac6998ba7c893c74d39b874d9c54493f681d078;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1586aac9555088b4140b30db69138dcc4b48834efcc16fa8d4715f78d21b70375a562737a04cd60b4620796408267112343001d47263a96337072f93aef72764fada4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8007a7002a7934322b9b50e4802cdf5ef31f2415905b267f892e12d3c34f52e8914b709106cc20ee594f5225cbc33872211a2206787093be7bbe6f0ad0e898c622e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a301219b5921185cf44b6857e2bbad4c7602a26f4dd51d67bcb8165035689eee485ed7b00a4a93014e436f10ba05c6138b95282128dbf95df7e75b4f10e6c4ba28f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e69d778d4a0ee315846c6eb85a17bb203c1dc49df084dcd1d9d1789006a11bdd08c4e1cce4bbe0a93f578b9cd6961c409bdfc52f7fa2a136151e27c315a25812d688;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a699610c6bddbb2e1d96718a9b45d4bde0c607504ba918c0ef8936be0d83db3d2373ada90e1d46e32a38c67c2e6628cb15f42b73420d4224927317f9f061dd0df4b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha2502cb969a63114710ca7aa3b0efe0b482748db1b117d0ee79bb5d552003c9bb1b5c4df6180729f2446771b5f596c8e374d5c94f18c7ee5218a54a4af07e7b0967f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h40091ffdce3fd016b03bf9d96a11228851883a77e98dc37552f89d14087bcd33ed97a2ce81fb49e131975adad48faaa01af23329acdab172b08ce1453250ca2d119e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h126a776fd0fc4e97cbae807f4d01d70d256bff939590af148ea7351d5df73282caef6cd6a32dc97df62ff7986a5281c8a7fb6074310836656d966e898fdb4ac7c1d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc13b71bff87908720144066ae726c9989f086d1062fde6eca10445c84e10b1bed0f9bbcf0118d040ab42ed6ca9756631cc6a9b5d415d4583baa53a631016ee8568c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h151ffcb391ad49e11c3e19ee2698fe6c74ca1aadb53df18261294776bfb4d89853e5dcb927f74d15d31f0fd02a61b92860aa7b2058aa6454544d3047257811662c09e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a231045b2a832703ae29d6388b0717cae1c4fecb74795e73dbfc80cf80c843f18cc71a3fbd46524d0556607e3600c69019d7de90fdec2c3dbc28f57a67780cb1e3a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he072186eabefb2ccffd202b8e38d1c14cddd9e44ea7a32c5f9b66bbd69f4c9cd20f95b7d349dccf5a1fde8da0bb0157f4f5e3202fcf176710e792f1adad5b72cbb32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8fe3e5dee781ce3b790fb365038024ea28dbc7ec73fc04759d12b5c48522f911d00101c54d940c63ee714de94bd36efc775f107b096cdc0f2b8078f1d88078c9c706;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h436666ea0b2bcf35832ebf261960d311c00e65b672b1da6bfe04f678cb0073f97ae30851bf35ae51dcd046d2bab6e906bf4fd37ef5b25f69d0ab6095aea1b806ab6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb0598e43e68f868605d5707a7916c48a7d241bc2a919ceb8ebdba770ed13df5a4853a88927abd02875501a87a25ba869ee2e60646a2231267355275c59c8e6ddf61f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2843dfaa0cc246ca9ca0362e0c9f0b7ff262b116192faf156a65d99f2a9ed8227b00c02f2aeb474aaef0847bd8b27323d4ece68d90bf4bbf1d06f20dc60f230471d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c4d0d5bcc7d362ea255e352e4d04e0afd72d7b2598c75b6bd8a4f32bc4de95d10e84472fe5d11272453a8fdf97f093a471e8f11643990d563696fefa4e8d44fe3bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h85bec1eec5f13dc1b65f79ff1fbba8d7ae63a44c32a44b4c17efb6b9211e6c6a38fdac1be722f82e257a15afb21833fb7f86c74c704578ea02d47d638d40ca66603d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2e04b5c67e2ebf825bae805499ea1f6d338082acfb6fbe8802e527926ff11394bd5858c5b987587c82915de37157607761548db6609e80120613f2dd9069cb12b69b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5497d435c70ed4260b7c1c8668bb2ca8a00374dd2e3cd512f4a25cd857f624452dd9c459f2dcff25aeea8edd8a9199878d964e81d4712ceeeecae2934b308a189436;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h134e63f646e70d40fa1347c46fbf0fc95123fd7969613e9fe8a7ca3a9d7ea7fb1c9d8cd9138a4106dda4c7972d8dfc8c4ff493208e27cab2b7c2ec3252637e840bae4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h134c3cdc70ef6dd2ecd675cb64735ae12c484c624ed1e2c8efca7aca928df3d958431cec888368475ac7b7de29f2eeee4a1548c96844c027e073e77dea87ffad9f573;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1555e4c9fe20fa8a299142d397331045822c48256ed0d634503349efea86411452b7dbea3f519217d0191f51d6ebfb66b8e7c5a9dbc0c44f58243bff4acb565c72368;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d909fc612f6e1d0e67a72fd1188a5412b9ef26351a2cfde24fc9971209b5e0d8a5580993734e61ddc90e0c038c7e8ebce1a44dc7e105ded3856e6d08f90df9d57a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f893ea0682fb10a68dc9d75a486e8cdfa6cc02a3e3af0563baa6d7d53c2d5537ea1302ea131001cd811421ba51bb0e5f085705dd3b150817350a553dd441efc2b816;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103e22e81b74bb7ceef5ac77ef8f945da0426afea8b955d6a34114ac39248d2dc62decb296ca019a897a82c94e9b91129b256030688f38bad1125c6c1e4c72c0bec05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c49e95750df202946163553da4599f21859a0ced0269fad4dec8bb68f6a2ad0b08fb4cdd1be7ce046bda0a007204cc708027df07c813f48b8ed9660611157d69f48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f2ff5c395a062c0edb421150da7c343ee04adccfb4a57614c727dfbe700eca32d32cf4e9daf6bb0bc599a7e29ea8873622df5cce6e869a5b9759b14d678b18cc4b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e0eeec08e2b0b5ad31a10ed399fbc07de7429089c0bae90de6bea59097889ded7faac0fccf3d287f789411d4e30fe4d7c10731136320a2b1c098c36dc3fe65c80108;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd849a1ebe7d6c9755f9ee9b6d9001798bfa626f4149174c6da31271dc0715b8e66991a9de3cbc71fcc46fcd9f9da7c29fa6aeea1a797cdd401050532f3607f3a69b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a637214a28583c462a35c0861db39dd5fa561f7fe1f2ef3d1f6a1d9e6ffa49fe21ea0e5ef0f2dfe7506d08af8e7c21df3dccbe147eeda47902292d5934009f67d627;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd121f108e323840424ff7181e2310debbdfd39db36ee19cbc1be5c927d74f4182dcb3afbdbec461ae1e222f3c44f3b45c5e6dde4f083bfec1558234b52f108fb63ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d6940a16d06466c43cd6c29878c46cb85417f8e9c675e2f7944251e2d0a9fa591869569e18b1aacef839b54def410571b7228693a3f049057e35c64322cb86dc1c50;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11fa4dea1b45713ca4b6dcab9f33c88649cd01e77ff34c0e2e51a57b11a6c119547e216f2e66e604962ec5e93c7a445d89382a2a514e9faf98564f60647c89caf9f91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14f2227a540de02fcc6503d48d5e020e617f024d8ebc052e0360fe8885f1b467bd398a43b29823d5918e7873e03e624eea77e868f919d87295bb3466d35bd15a4a2e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc32f63fdedbfbef88481c04a1d1ba7ab6c889c32cdbde26a0df4b4a38dd8399494313d6dc7239161e5082b6bf44b24046e10f6d85ca93d8dde3ed8f858282968b45a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101032ba5812e25b1f317b8efaa1d6ed3aceaddd1beb8d77a870011dfec5ce47fde116e5f4f7f6ac9f0025f074a003fd8c88160813e85c1341cc2673bb815d65e7968;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1963bdd16a4138f3f7ba072411fccbc5f3553a591aea35a01c3d8f4a7c753bf7fa764f43a8a3b830395e3ce7ea8339c5ca2b4fa086e1c9b9384e96f939f0f39924b9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2d4bd867d918844f06e2ac9e81ccf08161ec562859493ba902ae69cad10ad6d5ac7fa08503a0d26239173264f188400e46b0742522623ee4e30b254508e65fcaf73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e5ba2f7bb22444012d7675c9a58d26e11cc57f91c4dd9d64c8c3b0c3e25f719e1fa3884e6daa811755acfc5efb911d442621f04a6e83e99f57fc3f1583c7f6fcfd22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa05db606eb05f356113424f0148ce654c48fc35b30863e3cbed66c412c58ab92bf61f4357847be4a47f34c680bdccf9b521e9f19576167f7e6dae94434ca4aba08b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9ce3abf3de1d57c797066b29398b95b5372c56c3935d72d277732781dee39c3f70820c8aad969007f3ddbc492254c7ea9c23424827528c5bad9e4f4de458bf6b528;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fed8de7bc46007eb503bf19153d0b57abc6112b52d5c1ec1038eebcaa167b3f43df9842e7a171119cb7af5f4d11287706881a43bd7b6cb33861365d9b7e0c7e7aacd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e3a6ced2c772e3f85c1767654f780216fb11291c407436cfc9fdadcde7b168e0f9f70bdcd39846f3a8f8734973dd8eaa125c94858907d4a509813b14e4ecd81edb53;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13ef6ac883fd7c0f217373e72322904ca43e81976d44c2ac861a6ec89c2844e8f9e7399f4abaa82728eaa29116a3b26ac3360568962278e384b641743a939a06b5d98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89914cf20ba3155533d318ad7f4c254dc813cbba4f286665057bdfb5d48f5c1a45533087f1c543a4c38c29b42e15c49f76c32d8e402105e8dcb05e073994a4c38ed9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf36a2c2c911fd0896db69d96213f9b6eeff20e29e04ad5155866c199f4ac7b83a02dc5ddc45d12d30d51a889545dfc4cedacfa47450de4903ab084e9fb4e4f6d8ae0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h701285e88eff86a6895a66f774fef18604105b98b2973781a5101daeea2f3ad30636e295bb2021191893fc77c813a3da7addbd899f3141dc8937780201d80b77e79b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h952642b79f19bc4f514c318fe403168393157d97e2c62c7f27d065bac6cfac61bf4d57099495d2d74120dbe9a1378fee44c68064b392c410fa24b60743b89bfe628c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b97624cf69448e8e654ad5023c97949557a76b7dc56dd3496f6d78757eedec24a81ad383c64345911517ce9a537e5367d4ef400db22cdd134896018383fad00b6b05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d5965c9a64b62a48d5741a4321119e98c702dbd55115bc9bf322e4cac158234f93435ed0af0964b6bcd87653396ad03a57c1dadd968de8342563c1c82511782c641;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4ceed05646889f4d93ef915d2486b4f9a4f74fd5037e733680beff4f40549348c85c534c1421fab0d72a83f7d3ecba566d466d5b8e4257598171ff5294b94937e43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1190ac549f08d449c9ddd8d75b1b4eb676b204b5304ddd9bd14a0639c8eb46d5e5ffdf4d098c1c200082f657a9376e24dbb1ee8bae8efad60dbfc81c3e1c2dbec9df7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66ea02c39968a9358bfd5049f4a9ba2377f5e6d7762b59013df9f83fdf0ce50268c9d4da820fb65d356e4e6e504af6668a71e11de8615c477b753a45f031ad40aa76;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd535dd0a2529346526a036cfb5b15db30cb942189fdf2710fabb217d5b9684cb16289ea6ea15ed371275541ecf22df403f2293c989073ebb10d2927086d5bb9dac15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1568d42f445c6817c2a279c5b866e6e1d753f60d534b02bf90639ef9c178b78cee57c438d5e3b8c4f8971e75c5e78cfdf0bd1d8dbb55e024b7f54ddb0c003d76b83b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187e97fbd673142c2118f4b0230447a4a8a78f2105077e9b33047caa3adc19e3d93840b1d914baf91b3231239eb7cccaf3fb3f51c7232f75b534f7d1affb03b88dd41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b746acd4cba193a60c76692ceefbed436e57dc3f8068bcc991c4d2d722bef32fe7917d8f397f8b5d7ed403d9bd2696620625c460346498a09d650673b9f7ad6c930;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd094224cef4e0f4b360a0a26da9eed9f9ecf7937c2f19302bcb4918f4b3bc008402709fd4f1cce0739cd4ec3d70c87d5ee3f46d474030bed93c1fe476d45dfc1ff2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90b7fac6b767cfc763f5cfc4d3e1923a879dcdc1d24b7142140be91737a407addd49024d8d532214b3398d88a33dc8962578124e8295f977ac3f24fbc05546caa7fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d18943184a089a697aa3f5a66a83fcf8eb8a95449d2f68397f39823d6357054ead425badc555fbe019275ad8f4cbd59ec2a3603396c6aa8362080e27e79e85afe204;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10cbd12aedb87ce41b5b966c4ef526997774e28c121c1ecf690f7d01648cd14db53485370514ca21d4ed50f62a8cd96de221886885a2df29fb29f155d182d3d6c46f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53e3e656dd22c14c13828c96f45e5dd743b834f0d95cf58d706c949a91aa4d579eaef05b760c54e90ab39ac15d00cfc58b2e6a458d6b9982dfb03c69cd90d131f8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a489986b27f2a177207b534a9d9eb3d95c2c2a1805082fe129c71b73423fc5eac0156f8e28fe39948e7202863c14a164fd423fa2519a58c30b95900a76ba34c8d87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h184bb25085096ea63466bb9d0d4245f8a78fc1b5aa0598c9ef9ea7ad8036e0859a361aa7ac06bfdd78d19f1c978e12c709ba3ace014224964072363b5bb630051f303;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3bcb984aad8bbe42855090e99a5135c72efbda1675ade364e48e06f630a43509ba86471a21a805496440b7a51002b29eee3e01a0834f77e3d97572a140ef94c0b886;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc39970cd550407bee6172ed3b3a6530a2e356f85ace9b950862cb2d083ef829e064372ac283e7442995d6e1749f1fd47d48d9280a6328a983f02b1f1342922ab074;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e300aa61b7d2f02849a2ee874e91ac10be82362d2a2c058d08a0facb4df87895caa9a2ff52c393e7a72c9cf26f0a00f8a40c3fa43ae3211de40a5cf1756eee01c63;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19408244b7e46278ce73a28328a4652582867dc6aa388f537a1fa56a8aa126927fbc91c1af094dcae271a0b6808eca1c9a5aeb96a5e64068a08bc373ab237559b4b07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e4440cdf3478df042e724646cf9df8953fc9a4fde3be5fc04bcb038a2c3e9a08eb461219f4945f0667973d5c4b9051914b777d81293cc83e6099cf2fad17e988750a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h509185958af6fcdb18e721f1925a585e25006e0c6c83718c707d96e92250cc00d2ab631089d0578dcca9f631101422c7a6343636b9e77e5f1ca12f967082d5b4593a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba2693606ccff494e57224cbb29509f23c49a31c78d2ceafe1993e0dcd02e4c0257ae8c14c4588b50c1d7c0e3ef52e658fa1619e2882355d19bf87809fb8f54ef26b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h164a61e2a7237ecac668d9a949cbfd55472947d28bf45dcf3f812f44a3d07a72c697b43bc74ee1229038d31f55efdfb7ee9e2e4eddc09b9fd662bf789a339cae417a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ec0cd75fff11e63c6810329bbb525e4a3eb1ff0a7345b467f559f25c1ad45932066e3424eb052dbbce5333c590699439ab7923505df18df38501762983bef1af2ba0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h20a21f748ae191a7c9507c731033a9cb4d4ac89023913ff2eee732079d85a70ec7fdad7ba5de04bc7991998c94f16ab564aa8b0d6e0cc5ce96ccddb262989bd4b531;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h857d95a932435e27e627bbe553df92d48d735cd3ff9fa66a4bb94e8f2e26eaeb54d3283194602741177233fce0224eacdde107842faa19b27e42a1ebf5c5d02fbe64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha3ebd4a26188f106f847e438471bf53faf1630900716a8bc42c8da0b962fc09993bd04fb1649a444613c5ba288322610bf7e7d86a06e7808ba973c8564704183ab01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10470f38ba054232f482539e5a30cab4e5535d1d310841b73bf0cd2caae97ab5751ca628d64ff8ceac775d6687f15f8dcf20eed9a9e53058b95e29156fe32db89aca0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73343e129448e6bf0cae91d126967f17d819161489622b42543fc8adaf60110a538b65ae3fbde5ffd39ca9744940272f31fa911951dc91fc696a033f158a534c9889;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1836bb0ab5f18fbe4f975375ecc2b3fc3dfd1cb934ba63dafd68266e18b86507d967b0a91810eac6c72505bcfa1aa33ad3a01e10cf07847516f0e08ef6b8d755047d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e6bd430be689ef9f893e6b64368cf622743ad348b9458c438b944df6a8c5ffa9420e39e36761e98f578f94c2f0468d1f41ee54c1e22a9c6315d69b34964822a28bcc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1460425cd10253bb314291bc8a13cd509d0593a964d5487530f3a33faed191ac2ac2dc0d59613dee9672c4e45f687ba611472cd9d6c9c4fbcc7ed05d66e9ebb50c5fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c435a40921a21f62ab9c396e885aa61d81bccc31ca1137b1afed5477d83746e3fe59af9bb169862145eacb0b8d4841e9c07dfb95b1a9fe267461411af3ddc846a45a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa4f930243addaf517e74589f763982eddb569e824441a0a189b0e22207115b7932c4d131d2c283c7d5bd0842e28fe192301d1879339beeeab0884e1bc195be8cc95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a74f07b6f1983615250226e258bfa83e31cccbdda9427c71be916201f44c6f18c9d476e6577118a2388d6d8c45438f060539d9a097280cb0a748d5848b7f0b80a742;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdfd6dcad44c8008a3d53631f5d9cb791ecfc51364f75f9ba93c77a67882240b8fce357d54b201e8077fd3919c028315179d23296540ff8ebcf3f22db71f4007c6bf7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e24d83d0e5559ca779a8900c053b4657c65b88024ac864592227b314559b1dbefc965208a6e99c4c085279c5ce62753514f5d726988407de71bac9a70fd23ca5ad9f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5909c6179bbe4dd15e3f0a87ce90d359c8527c3ff736fba21d380139a4f7a5a70dc0b5c7c5aa6d9a70617361aa73d3e0eefacee98b70343a0cb0557386b260f7304f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf6e54ec9e85efef588a27cb3adbcb073100adc3bc363919f7d1b68f5164d920caff28992a901642a47fcaa6a7494f04f29385bce3e275ae53e37d73aef266b728775;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h595f7806014103f357a1eb5a0cd6dca1172036b54c44cc3eb077d86d46d5e704e95c089172a9fb4cded5b9772cbbecbd0221db7e6dd16989a7dc4a4d9b816b52f30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha669f19ad7b9925f9af44b1958e8f82a24b6cafda68c3d6b0c1334eed211ecc62e80ffe9b71d9fb74824644733a95f7cf7779164636c33b6bbd9e5d6db7a4ead59e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he7712d2af2261f371495dd36c95eab527f5bf3cc4202e5d7da5c69be4906f8e28351f4de2255811823ce47beca008a232cdb31859019a65bf541c4a9c05b1e96c1ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1459df8c16b57643fd7f0c2d12bb85f0f28a75b074f1d17ac67e2d8b7bdba0f0401c0666380b3ce8151208880f29f5cec1edd1416d90c7ada2c003a97722b5e374961;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdff12d9efdec27a5c14a1ede62ac248e4086aa5dafbc23a54aa378ef2e7cdeb61ff0cc928ccaf59d44c6de77b302dde87ac8f3f328861f276758e5a639ce5f840be1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9872496e91e5cb72f7ac8d11369120a52541024523a7a61739374ac304a541f3a25f032d7c64fa81a6a8289ae5bec5e25172fc43a8fbe82dbd9a3f4c0d56b6530077;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea35ee3803141df505645dfdce76f877ea0d9cd9ff31b9c73622466637353164abc49c9c73884e0c442f3b20fe7db9163449ea7ae5be9d3b68e41bed934c5c87b7cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hda017b8417f9c9d8408ecf827f84a8386b6e768a1c94b24179381cd8ab355a7c7f3b647b96980766c547dcfb676c784fd320b42457aa77fcdd73ec9933c56f9ab921;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h638512051806f60c10a2658f8dc26e919d0176628547bc74d70e4aecc5962fddd032350d12c1c113eaf372ce3c0471e7324d244aebf1bdc8ca3bdf4d20499a9db2c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd8b444a092788b9b811c765a3f228b53a696b53915e1fa3f4d1ca91ed149877fe0eb7940b2863745f0809edd2a939eb0f09ec7faed5361d3b318e8f4308d96de8ac6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e45425042766dd9f3916edd6985d2f1786ad541dedf4fdc0365556f2c1e3e7bee34c3e84aec468276ff67570446c4ddeee215b50190b3e1b89b5c94bf17e94db27a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7da276b7fe9ca5959f0826b8804f538939c17376959fd440351378b79b27431d97fe9ab073e5711efbb3ef2279e378f1966365fb410c2b7aba513ad4efa8967c97ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c902f8703053be7b2de087ab3ec0a68238afcbae3ace5fce115279bacf36b3ff5bab928fe65b54bf41c1bdeb6f94b713195ebebdf086cd5125231788469a9eecf74b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e58d9ddb50bdd619399604a015c6de318c578883ba8945dd589a228df0da4a9f7059d044e724e2ea88896e3291bba51bf3e40c141fc7ddd2a792505504fd08917e4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed22ea56e5432b8dfb2f539c35bc33d0a1f1124190eddd59b10b54e25bf890c0eacad1f1149e9f24492e8ff3c8dc8432cee2646da8c280b6ecdd7b877468888786a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h183edb0e7e16b613cb3b389a8b6dd02e923aa734823b749e5bcdae9444921c321384010e2f2cfc4ff690fb82b08e66011bfb3c2b35bc95df2ad19193c32e913058d46;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17d8bdf02ba9fdee2162d9c3e7303fa118e155e90ce01bc4132a91366dadc25dcaf1d4c44a084b406345d00c4db3ba356a00707eb86c077c935f6df7b3f1d075cc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc96b1ac3d729705bda5a44866251a72049c35ec723b0a9f9f2551c9be2ead63ac3152b48a1c441b13cc917b7a835fa607615cefb8290ae82bb7b3c86314951ebf4f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h144460de74ed28e08ef101152f5928ea3d1f7df647093e27e5f6f62c28356d4bec3b968f00ec3ff39039e0b721bd9428168274d2b94018b0c960a0a2bf105e7edefc6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c898c315cceb9e3c69447c5e8cf1854ecafa7ae0e78f421239af35ee7cc6c5cce8cf96458356be7f2db0883a817cf6d3a3fc06e2262a3f153a5e8df2cec1b05db62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h128a12e4d8d66256411280cb924a04fc3e6d0cf4a9725f3c213b416543d0acaefb86d3546b247b26aa01dc3b7e5dc7947c515da6a36996439a1d8b89c50a67f3e2bfb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c51e47070a6aa87b3617d910fa1ce34572fd7d965dff0517a6c58f6ea06913e039363e1cd402b8fff4e53db2817fa3e6b8e4f57b450e28aea787e5a84084418b21d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c80eeae8e7ce3d1fd5203854e6fefe4e6ddca58af7f67e2d4bc4212aac341c145c6eb0678fba0b2de5a35f82e883868069ed009b42d7f6d2bd79e38d0fd997e4a575;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h148e12493335642898b58209bf7d8c07641b0c547dcfaa465a1c190252788853b92b1d48385b547ed0d921dccf055ae199cd1334737d4546b8736807ec84849d08c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb16379af5010d93959e1b264912bfb12e8e68b56310b2e4d6b6682a129ce8772dc059386223488002d5d5da426f325102c6cc1775a3ffcc371c2c26836da65b1748;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a46951302f6b8b05867b9c531fe90a4b9261f9f29c2f0c96737b2a4f45c1c7bf9f472f64baa965ebea96954577cb121970df12554967f7aae649050e8d1579786ff2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h329f2f781458bb89c322770c2e6338b97eb884f90abe17371749bb94742c3325cacf9ddb9be79a7fd8b959b57208e65db4564e57962875994f42e7031d27bcd0b481;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9c52448757b087c1991222692fd3b33454b0c8d037c8c43389cb0723b3e52e0ca16dcfc2943467c6bd0270481eb33ca674d5b687dc9e122c5bd68eab60280e59f8c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h81b8cefa4c0724dc9738cf86c673c12ecd635d292669a987ed57e3eb22a8299c30d2a9eb76780fd5caedc5efd32e44e2744b0e3ca2e41f648f49a097740c79c2dd7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dd7f8f48b48179a6fedc3eaf23130ce71e0793c5977b91eabb4df8fb345e5abea15db344d212d37a4a039e330af8ec244dede7fa4a159a9f0c8f2599fbdf5b56e693;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ca19ca44c1f72edda2fe55e5409625c56080dd7f69145012b416f927be188697a1080d0cbcaf79686058e06faa7b4291f95ae34185c306fca5a3715b5379567d2dfb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h59b282b9b2af36e7ba99fd68093524f59a2b8a75d5b029e1e2352bc3e4ae0aebf69455b772a3637f782173baa2ae708c4b5ed2a32450fba55988240e469938937119;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h408c3c70187386496d3fd162de4d84b58fe382fbcd10f620aa80b90de545b073bc2cfcd4e49079d5a49e9c183065022f7359f46fe4294145be8b072a2ed3ebe9514f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h173ac42402334a04d2af654521d1137b8708c319da4c0241bc42b62f3cf8d7c24d9df289d2898d053ac1042d87f0c88213e34099cb09cc7be5d27f6687c27a23cfe9c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he1f82a209da3080fecb3c147cb38c690472ac335e228cd9d08a421f158255acca617b36830d2cdb749cada1b0d952d3c946e69ef7474b7558226f7fce519d228bd8f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90939d4aeb7e8b2fe1deffc38a2800b2dbd9452548f9baf602ed6aa74dbd5f1cdaac7f6dc011a4c83861e6ae8fa2f658ea4690af044a02b242a663fa87cec047d2bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15266d851ec15344dbdadccb1e2664ab565ecc2231b14fa6106b03cfd2fa1000a5fae08071fe214b99f4705de346f5b6510bfbf068b9edd683d53caba7866af8d06fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1715c980e3e00d7cef422662f4e4dd930417035ecf4da70405cb67f972a61c5b9b30294679c83d5d9e9394413381d60aa0e19be6203d088dcebc0ce2f44a783be5a47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5bbc642c623160bcb7a30751eaa89ba9284bd9bb44424d5e226311b8883430c481252daaaf0c1f7230c5d2aeecef9239cc538199889dbed2f623a9c21c325df1395d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f26416d065e6c09e84b19581660919f28a17c302d1b71dece9bbc60e1cfb18b708835c388290ff9a811a5e2808482c05db2e78e8dc9a8bd2c20007bced8b0c7263cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff4db2aec985a9f3b550c968ba4c1c8e800761aafe6101e40600714dee379fd7715acc3ae3adc0a3801259e68593da57033e6feb10504bc07804158278d25e4f6dfd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a9fdfb25595c615c2d57b21700fcc5938e2306c9b784cf30db6769526ddbd02927ee401b8daee5af07f667b71657e2979f2ce5a6b532306d670fae3d540233fc958;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b5f51e9f39e5cc82218d4e109b80901b4f0575a3a970d64d48ef155cb0583d484a78f59fccf9505cf619e76854b76a814a7e05959f5cf37d2af021b1399e7ec4fa68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he0d944545f3d7430a78fac4754a80169ab6cf8135ee0ddd23a1f43f924d07b89698ce2c216e26b31792e2f8882eb69f1ba480fe275f3ebc479ec4570e80be92f7895;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h65f6e70e1b849891fd9f0448b71228fd476abebbcfb67434da8be31d3de7135659f5176293649e2219897304b414c527e279b044f2ca63aa49b84542b70f84342636;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bd364ee8896bde471e5863e4d69164a9a9ed4121fd763a2b4a1bb468d4954bc2cef6f6a024404042d5daa28ca495a1800c276ad9ee692f323d066638c91dc4759a6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h178dbb71116e034df60f897c120c58854e324d0755a66aa5323b8c2a13082c7561ea065ad4d4b92670d1b2ddd4b48f8b9ebd49b0b743e71c0e5acd8901aa82e30a548;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h111771ef84fb28c914d7c4e671d8fae2061bd287557a843ed3f5d3a41eef3c8a194e62f34852de9d3d599142751ea94881ff87d6990ad5f2358065ff7a9c2a7065498;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h386ec8498add3178d055504c8b70ddbbbfca84bd9b0a7a0f82077096b19a79c5b16d56ffd83901eb295523c5050f9884b75f713d5bb477400c01707c9a5893ad1b3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cfd4ec48194a7bd22516e0d1956bd072c6f63d59137e4a2b3455fd06898ad4d8ddeac250f1663f4fabe8ee5c1ed442a7256f9ce044df3e1a96d35a625909080b73af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1efc3a9a5507cde9ba6442640c28480ffebdcd0126d96c22dcb6e47cb78b6c1f1f736d8ecad0e9ab22685482e19fcb70b23244e5a00a48e19fa21ab290fa84e8c091c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b6c21c8e53623b739baf549cbf4a9e3716dadf2f115ecefb31f7ade7922d95dc291611ce673d9048348f7fcff5453c9611c1e7ad54ac85e8c352906aeb1eecced80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b1308b7f09748ed3b6a9b9c4bfccfe1e8ec67a04c830e0c8b1d0e9e4952a7bb25ed85b8b5c7c2fd80d2b0eb5141afd225314c4c8f15c14ab8ece2df8b08054f1919;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb0233e3024bd2560d12ecb81f442830b953f634c494d54913df126e76356d6f3aac4b56fe6a8811250268a85341c27d27443dbb5fb42dcd04e1cc9fe906c83021b3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h72f08cab525871715efe317211371a43a35e8e4064631c48536be3a558a73c6d838755f1d31841decf90100b2d22cbcedacfa4852736b9e04bbb2321392dbb40153c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c190cd8e1f88b25ca5404d9c3e2ff026cec3e5f220cf031cf6de6ae27dcc2fd2b8c0130594806adf3d3f0403ce1ec7735dd746d43c531692e2a28871c45b2054eedd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d11f333a11890d6f2ea43b9612a2e7750046a2aaff82c2330a5aa595a8e78ee778941b4d78a501b8af53890f8c14cf1442d6c782d37862314e335d2b67a2d0b6085b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af3c229eed6e59252768e83218f47595f1bd40a1c8586b11e32853bae29a87fffbe5a0d23361d32825d1752b67f52b1b1128a474777f3cc420df16626b2014421be0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc995730ef753323341ff107117de68b820d9c9330064fddabda24af889cfee024b2b935afb093fe9469c8582ebf196a3ad9e6a3e272bd5659e143c2ab53a681772da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3aaab8184c2db42bf93436f496bb1f364ad6e713e8820cb4f3de9a4f194553d180af8a2c659d90f9b1b97c6eb8d00bff32d9c91cec58cc54059323eab97e8dbb0e87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f98844dd101777919c629f36b1e6e8a460802bec0457442bd69180c8a1e7f81717f919c7b737a0f4d15b461ff6112a81876f9bfe4202e17ebc0beaaf98fbc9b2010;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba8980e4b1e7737c950d6dfb75939f9f6ce6125742b2e171d734d4a254ed145d6b17cd8ed44e4a7c91ffd963d57fd0d5d7ecf58fc5006f2d309e8219238465aed416;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7647c3852165adaaa681f2bf1b3a18e358d07b3cfe94bdfc7d007cf41e1c4822712f12862483c8f03efd164a05bc44282757d22fd185b00807ebeefd7d5460d861a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b46fb595ce2e11152162c9c9a0c6b46f4ee38a8ab276c7076c81c75be60964af074ee42e994605e442858ad3404f2ee6fc672363acd3dd5515d4f656136838fcc913;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1beca7f8655db1cde0432a6cc7d8145081c16a425ac5f25820104fc355bd6cc84f54ca6fac847c819b58a5f4b3d2fecc584328f5fb46c262ddcd27a699c88e52c1461;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h195ec86816ecaaa39187baf5123518587c9c6c26ba53a8063046fde7c0b24d027f748a7976f225c61a11396f64b8f3645c3729579ca10f054f6d6a701f5b402d50d5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h46eb69b96bd5f3a85960878f20975efe5d61363dcb4c83df61bd76fd76fa0c5e4ea3e0b6483d1f8faf4b6170648e90015fd205ff108d2620d2107d6f36e844ea3eb1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ea51a99605931d7f2b08b036b23b8e12db44d71ecca86f719f4b79f2a045235c9165088eae717131a8c7605ec737d3a4061aa993ed0f12f440b1a611a2f2068bc74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9797fc82d431225c5b34aaa83d93594469172d0d54fd1ba76aa29308c409e6ca3093dc6fed2bd2d509d299ab4da0c8175831f584b9286751365a53b62856c47f49e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f935019fc5b3aae91aaff4a66a42cb8950860657d30086efc1d6d3d1ab456b3f3f67fd9b8f48da6a7aeec23f76c01bc7dfec2cabd627a4b4aaa2e1c258589633c05d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h141a3ef459f1514b96115e254ec4cfcef090e39a50ced3d2a8b2a2bf157e186fef0911bece7228c8ce959dd513241510db7a669bc8a5a02d41c520fd60eb53ecb03e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h42cad25563c56f4961b5b667e201666007d6d8995f706386a62d9438a3a17630dc410fa9a3a0f6104a546ed88123b2659bb1d59dbcf7581e170f100edec21ad3b6d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h937288cc0718d3626150e4caaa7e679585dac957abe9a326409d8239130a24d189c9d0ebf8084794e98d89922eb743dd01e358c92354b339eaad893690a5a00f264a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h169a72a4a9d6b691622a0993ec97a6ad47f39d90e3690e323f2dbd1925a3534e394fc049fb02c2f90ea10294a5bcf291c9ba023e909b82717188cf516f78f2566a521;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haf8dadd90c21f70241979142f7aac840777fdb615f41440b439aaf177c1c36a05ae9e7e7a3f2d197ad06c9104865a43acc9d692a5ebe2a80c28e0af8ef51bc487296;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1382958e9e5aecc5dd93d9706603a7e1bcedb8d0534825e9e536fc10171aa9bfd6a94959e50f867b28095c3384f328e4cbc73fce08a78894600cb1f0ef7756137997a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8331cc9d1ef0e7dc6c65648a3ee6595007974bb83c2b14c6e8696d5d5f39b04e632725e07c4d18cc889e3707914bd826c52d805405283a8d00a1645a4fce40da3cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb6ea4d81b969a9855767206abc187ef1801082657cf4adfd29edb7df658c865a946a375d8c27158ea13f114a856879c95c00851288a11b89040c85a4686706caa06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fac81696fab62da5a19e7d626b29278e557d6711c4e82a8714a8300c4abb8be8576274ee17914ef5913cec7e8794613de0eb5220a38a08827b053705c1cb3426e4fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c24cf3aaacf6bd940c172183ca36c3d74441c0809493e2f8ead737f9d0d5b184fd590c23e1c8b6df50c4b5fb3b3c3941355411c3cbc5860f5fd1440be9615701bfed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ec24ebe5c07720f1d0f2ddafeff9318ba149680c9c451a6d9b6c94240d8bf7307fc0b9a0d9daf4c1d71d139fe9cfe8522994b73aade64c8c555357799b388bf9ce1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1096f0ffe24c3da8da513f46647f872db44d4406871c5f5862ce95120bbbdfd320761be7a53dc200bccaf142827fb300a707db80774bd8a600978ca9f18632d7795a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1971992682d9aa8814600920bee10d4fac758ac3bbd8ec88322e0a6bdcf5fb582e412de0844cd40cbfc975be92a9a4fab4c8428cb776ba41764cec1eff96d9312126;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd5712373b6f01a9413bfa2808bac6e065d8bb4293d5deccc921e9882eaf316468be58b7168a9d5bdbe012b45ff6d7f6fc7a66ab29be02fcaf87bf022597a37da46cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d8a07832cc2ac284c346709970d77f407ee03e176cd8d6e88b8be1bd7d24677f8ff39190feb69f9e70cea074ba37f0c45b253c8024a1f066b4359e6f7018b4c7b1a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdf4966fb88924c586ef325f57bd4931d029da32d64804ff59aa6777aadd151adf13591142a68c70133e4c11b10bc0a94f5e36d340625a3bcf639c8742041bcb00761;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1855736812f3add4b404d2c5b9c77c0f76b3ddffbff89466f504085411231fbf1206ca8a6219ae61d15498b9a4d5984d9979f1091c8c076c41484b549a8e8c69dd16c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5579d7d4f63b0361e7a289f9d55c88e012f1dcc3543f71ea7ec7a042c1f8bd5dcca140fb4774f5e75dbf12153defde5e35c779679c42ba79caec9f1443af52358906;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19369c0535dea3bef294ea8e60071d6fc9f19ba4617509312173ac8bd3b457439abf078faf3d72470feb04742b29a9cf7625ae10403b971b61d15e00189faa0cb3c92;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hedc52dbfa69db26b819e8fd0eb1d012afdf09b0f378abd3c5414cf7455301ae81642391033f7f0f6deb6c76a63f405cd60c8ff314308034adab214eb4f44f2326f8f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19e5e1d3084d646dea1a21a5f2093e7bd232270762b13c2f3e122862120e87e1ec611884d231559bc945d12d07d954523c10245c94effb481bf8aaabaac01519a9e90;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10670455e7b5d2c269d6cdc453fb8d1bb564b3d7a9055e9ed9bfe694555a442d4466559b623b836a05db9cb53238acb7155a5528abfa82d10cee0f636d764e860eba2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c503e821b595bee73e1b88661eeb1f1f480ff435dbc9ff317b85a624744fcf98144dbd684f7ebe2cd24c2b14813008450c433177248ae8831a0873d6a992a779e65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16745836e0b2c9478da75aba1b3eb820574782a837ad638fa4f86722836055c8a15fc022c904c89f499c16ec1349d8aa3e95f9e1aab82ac4550f6d1035008e63d1a02;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h148de488cb3917bdd147539486dfdb0f044b724582f4479f9cd802451db494311c02b30b5ea4cde8271a3c1e7590a08fb53c1bfd2ee3207cb0367f86006944a51b6c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a11663b60ee41cfed65b5ed225369854b03e52145d6c661e5ff521fb5430407fa9cf586fb8f6c8cb26e38633becb6519dcc624bdddb946ae64ba0d90aae9de3e5675;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d059680bd7e5f73e8fc79c9a8378dfcfbe8882ae5161239af3c7777dbaed5ae2ea550776ce1a9efc7bb8acb490efccac37c8f216d6c333dab06828d245f2c1ac6398;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97bd40d8417631679bed07e495391be25d1785edd931f4fef3cf6fe69fd2b7050b48713dc27eabf210b518d88cc9326dcf956906b2842a4653296036c39d5df635c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2303d67751d93d6b1ad23ae921dbdde00f8a34a8f3583ac58a9c7120ee7c710724d027ce433523bd3de4f025e0c795ee5a159bba29816c95d7fe2c55ca4bac8f5ff2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d31308e7fe1a1e57de2348846c4805d2adf6cef76156c6bec919314f2d2504122d9c503733a86449efa7db28e8aa39e79ab1f6d91c30514e41268f16ae5d6cc8dba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h128edc20e176b2ef8adfe5aa5858eaba22ee9863460783c164f23201c76d4434007655c57dc03be2d2eb75ec80c1e1dc122084a360765cb1ecca329e7ce31fb840655;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bcbac95749ae2722dc8e50fa832cea48ea078e524cc44e01b92f3525328288ee6cb6db0a543c5acec6b36fe6cedcc0dc452456e81c3dc6db4841e64059fc2355e5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc83714ed06c98333292b0f15f9b2e7d63898a8888c5b8636bfe93140e333042b09465c6a9d19351f5ba00be4b772e066130f8a461e3d044d9ef4d174feaeb98b3f1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h38574b204c0bbe23fa1a2182578064d85e60deba9307b3ef74afe4cd2e3974dbad8852d67380c8b6c800c67c98a2258f8c3a64d1c60d5efb8e4ee5f637c26b06b251;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8bafdd75b12b559fec54e9d8c5fcbeb1640769d27923d4e05c5a16c5019712eec081a1b2f51c9f193a78d59d37365410d2a8714b498e90122b09f41bcdf3b4360c2b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1884cb3e68cf9d5b619c9e7a6595d47ba7493758a786dcdffcb4f8635411164bfe7faf25d79da165f222f3256d9f712b2ae0bc3e84e0a8365bab5a65a39ddad8e270f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1988d728c6e04138fca9918c5d3098f5a7d473a4e5717d43c9ff2633311e565702180b87468fa774041b5d22232178dfd380beeefd4559d41a94957dae755492ef1bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h299d955b2abbdd3f437a3e6b515ee407b8896875f59fbc27e3d15d55319bb492a344a9ad114a8fc180d949a76edf6b61f4c4de632ec1a10808dd6ee521bbbee4d639;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1384d61d97a6db0e67fed5766ecb4640a5471f12459c1bd20d1d4519fd6e5c8b3367754c636b87daf5e3589fb21192a6a07b8d357aec83f610c698d444137406a8434;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d730211d6a03ee441b448accd0131c23f4eddabc57c7655de4094798a4a529c4ca856e5e5287c580f4c4423dbb5db19a78ef9a3fef92fb788fc6523076cea40550f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c988f443b01fae39167d694f0e04f13ecec67acdfac852f922d399bce37d8da9806e60e6baa4bbabc2a0d991b1d9546f5a31f20b88f2620c56c8c68a714274e5557;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16930567835d506279dc1f98b277d47277aed0e029e385925c7d6bff1cc639080925e915842401923b742cfd6bc7c3f0f77bb7360ec5aa3a0b4bb2aa25cf70e5c207a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dbbbfb2528f3381c45d223b4c1c4aa331d159a55c6dd2fc3821a48c60a5814982e88c9ab6802bebe86bc835e5701348d53e5c6f9bfeab426220f82c2cc5cbf0a63f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb2ad8e655316c27d1206330c9806ac930e24dee99828f241ebaa7f9b928a429ccac1b8d570eb0a804a84629c23d9c02d0bae9e46369d4a4bdec437b24fd01c12e738;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3f36ff315d57df0e9e7ff49d81bff97b58b7512a02902161c035120d36e00eb5ec99c44f445337c81d7fd8f9fe5c7fe2d1475f74885495299017407fe2db689861a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1012236ee778449c685d0281a1a6a7241ee0faf21ddc14e2c69d42ea5000a4baea95f9d36ac450cbb52d19e1e62e7089192d7ee884a431208363d4665e86a6330ffff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193d370a4bb5516699d16297e0d209123251722006ffcb21e4362b3b495077e694649762e6e07c521c0ea1d4cff39559c367d2d92e78e2d2d84b29313300ea3938636;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a74bbdec7f03643806967e96eae1294b0621906de64059d40135d7ad763cd2d2c360beda96836d369a1011e6ce044b9e6fcbf0d821c990cce56a5f2c567b38f6edf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h65ef9ef4bb494be8b90dfbb26790d6de81a295e6f438de02695ffe971af6ab2201bf313842f2f70e2aa765ab5cea3c9060dbcddf074d1a7bd98800715dfe426e40ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h46c162e9f7b78f9dc42d6ea36d5ab5e51d9106b6b83dc5796b834080cf89de37df57adcefa34890b9a95be36ba96ccf50e4c2a3ee9df7d65c8614f756d3a7a7851f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12d9dc6197221fd7b79b35caebc1dc104b5fa13327fef590281239fe2a9f23097d484be95b0b5d2ed1a7c37a38ea5a7578ae5037246ac4b824b90407fcbb39b7c09d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1088a70a7fe803cd7409965590cb59e76e9e9d6ee0a1db6058865505db6a1d64b41e79412b271e9625e179772fd7878283451deb0e269ad5809c51327aeaf5d30c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e198b56d020052bcc54317f69219567a46238aa3931b4b698cc3b9d7b8ede18fe8744810e374dbc2602dc1f0a24a50ce2daaf8f0aa0f0da54c344874b2cb6fa51154;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h140880d2cc4be3d3db349b9deeb59badf4cf3abcf2a18a4a60cec55ef6d6fb29a4aa79a6d2283e81ad4a5cb2ae12587ae4a43ceecb77f4d4fd2ba6f073bf75eba8600;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff529d2e1936ebe5e8172b270159cc4a528f5a160ee048ed9b0b2af74a6f0e3f8dd9fb947bc4b7803c5ce127dd1ccd3bef3f563c8106d0f54aface6e9a404925fa46;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18736176064379513c941fdc4421b4b4e480476e5acffd6c42578abd67ad709e15cdd585a298a93d7e1d62dc6f9aa2af6d07dd1be66b41f2578c9a05015e30bca3036;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h52023358d69954b01a6a8e5a35ab7635e6b0765995b493f87452aa68129c02adbfb4e3a34eb51d37bbef0c7201d2087c29fab98fad02e463a3fbfe35e4547389a33b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h197b865aedd9c4c2083e00bf640d268248f316f87d3b67d69f22e2b704debd84e85069c999ccd5721f49692299412e3c426a76ad89c761ecef51391cd7bf61bf035d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa89b9ea9a3875d901fb0198cc07ca3257365fc989e6e9a86020df03d6a490891d78a8045bea56fbd371fe1d96225c1a05aed4049e4bdc1fc087b58760b6a70c6fc1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138991edfa051d55b54b9358e38216a344f50c0ecf9ed8f6fbe2a354d7bb0272c7e4f50b6bc540f6707da9b1ba09ef2831243758ca5d6b525214b941b024fb6e2b535;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d3258e082d414cbca07efa9f6357c8ecde7da864599249b38b94bdbe544fd81674f44ab840a1ce3fdb25ab699c6bb89269462f9a8881288ae8218993c90cf4bdcbb7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0da74b3b48db19c44e60de62527b7446197964568e665f6b5c8ac16ec137afb3d5490dfc97f0201683d11f921b48bb146dfba75e8fbbe3547b9b016c9551c14ea4f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ac3b71d3fc5fe150154dfac8873e477a41efc57fc21a3f03c33f8607de80775b1c47cc81b6e46c76ead89e2dbb2870cb719f127c8a4e6c72bd75240ddee6e5c24e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cfedfe172c4b34a5905f0482e5b9f8eb49aa2fba617d2fddd85da94f0cb1d45617d60ba30c3d35709ec4cdc6d8b7228979c2ad9bdb0843b55baa218c93d6880774b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haf252b8d9ef237796c45f4aa3628a0f0255567852dbb5f2548fde10f7e2887a95445d97bbd22c6a0157737c6939144d855f236de9c7e7835073ab73c6cea59c1b845;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ae959c65d559bac05eb2689030a49671ccc3674fbe5c241cb6880bb5b5cf9c3c086b6a354b4682b64d4963c995bb6125a4b688484956d7f13f3ccbfa86d7d293821;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1539ad9505602677bb8a6b13f61950fd5bf607a49211695ba68679650f1efa6a865ed5094684e8823680527e16b86a6f04c8645591627e8ad9a3a720cead4c83a9065;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19895f1b12c5da5ed8726c15dc65711650da653a3a353ad662854498cb343a8f2e30f2ac8ae59643f0aaed41c6498492f9a6e8bba6912280d8cf873b4a0d3aa70e5ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha9ad38b0c77cac8ff3fa83b2cfaaff28e873fce33e9864f987795d80aed1c6869c969233651a460204608a1c5dc0f1a9a6adca53f9868ea41d50eeeeece85236def9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1119fbf3c01e28c1d2f0359b70a97a6d9aeb0297e5f0757b009b607b5471cd3760007d617cfdb6e5fc4c94a531e6f36fe168fa344aabb7c8a80ce1ffa989a4dfc4ac5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c759291b9922ead7e274476ad1fe089d71bdeabbe7ede57d2a9a60ae15a0b8552da5e748cb285cfec1fd0d42bc84d2ba672a434be297eddba6ee5c558b8582b2099;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17411ad60acedf770f8191a3eb3010594fa843b8f7976fd8be45874472d2349a1d925008185d0a5af7da83016e8e1c9686641d88413fe0667d5391afcdbf087a1fbd5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb336cd57fb04fe23e588a72055a1c646539382de7e8410b739ccad5606be07422406b91776d1e8e479c3efd0e169f9624f4b4d2e17fea84c52b8758f4911bbe240c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h64f7a3d7fe3ce2a0d831118c46cf07e242178ec2238d9f6235d15baec91763c91051298f816af522df9cead5737d49e7fdcd8277b76305c7cd5ed1e41450318e146b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb73cd0414614c80f92d1d376c330beacc702c149843c029cc4e06557f9e471e32c3865902036a5b5fb5f0778afdb40224f19ef420f921cc84fad14279a5a0966a905;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d4789d589af8e63645389f25e764a9c532134d12921323f938932ff97d5934ec6ae836985bb6ade7020f9278405a5e904c2d3bf29ba1ffb3fb8629b7f94f6c1eece1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fd9b82da7a44ec72c94703c0d99726dcb0d05f2971c28120549142e345e156d61f5106ec0bee82529b596fda1b31e018d7f2c73ccfc843e8bca3d60a0c7e3ff2a8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171c0e3a832a9d89e6e446dec349406c4b20afb066cdf34f3131201a6dca16a3141e53bcf4a477e21a927ab124ecd90ae3ca4dcdf3cb2058d977dfe88cd642b66ef2b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11046336dc8f4bc5e3436fd99f41feb0c486234c8ca57e8f2c70b618e4207c3f0416199c6f3e91597d9c4ba31b9088b1a144a9b581d0117e485312618b6c3824e0c68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1151e0d70b92a12f2b90f5e5ed87abb041947dcd8c511bcb5e4ae06585235d04b449e1ebe8c986ddcb280e5cfa2d83f7160852a4066e7caab9a4031e697adf1bc6c14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3e25059ac9acd37fef09e5654884100fb4fc5b5e60a639af1dd1bf12be7408833e380d2b03f28e7e598cf40edcc6b1c40c7271b873573183b36c2cc9264778caa42;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b9d3377e7a3b836c929f44927e4619f812c28f6b7ff1139c8953154c3a7d5a78ee8a56b0acaff539b506fea9c4d847ba4e3f9a9df69827561c13712c616f812d62ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16346a23fb538bb416a5f12a65b8907fb8871275e889ed69c63ae189edda0d7a5b59ad26124432b71276d982879760781a100ea96d280b4a546d791adedef30571b15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hadaf4aae0396e1d4e1b3e6a27c03070777c0865a9f23f9cd6ebb4d8beb3ecbc73bb274d159aae7cc597c0012fde6ecf0f898893601a3f57e0a2fa84ce41107385943;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ddddbcc13684b3c7641f45e1d4a6fef4e3e2ed442392877f158c66606dc0e0f415b6ff37ead6b169e2b6b2475e2eb3805174e167641abc20387604769804b5f9ffd5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf17fa6e35fd4d63b8dd16bfa1bb07f7e904f92bcf715f6ef59d0cb7fd2e170915806e5f6094ad9a68d1ed477c07ed645d36586e8986ed72753e5ffc7d8d948e9939b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbece19c34f760a80bed007833523c197705f7171a4cb0255d89da43d3ff6d94ef0e92bcdc3ba809fd314527c3c66ea0969a421ae80c11fc719665dfb73f3a55f9f3a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2dddf1d59230734c827a02b77b7531492fd0c11859ec28696f6d822577ff92f4ad1316e60e25a549d294379f10ab5077e7e12a865f3c11343c23b916c45ac0fdf0f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb6cb2662a228703ad7bb01df32c1aa459fd0a3139f374cfb00098bd2b0993271a0efddddadec5549aa6b2adcb128bf73a515c1f0f65afb1d2fb8e5647c01844335dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8da94f188b5397da70b73bff1a478a0f84a11f66b6ffeaa326dd6963f839d1ce420341b21fefd19801cd4ad91e1fdd3d89cc309968fcdca093c5f125bcc66852e551;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1487a21d5daaa7fd1ca29f86c45dbfcb18273e787a67a2fa7ccff34f026f07298ccb11c7afa9f15728f4741788e0d0a91c8e654f6c00f4e2641227d0eb8afd46036;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80bad15cb19274afdb9da3a8ebd7f943d22a6ddca45fcdc82b8547d548cc67aa1424e5afb43b7574f7611215eac0b7cb49efe2a564478cc33bb9395749221a13736a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18135f1a26159c2b029fef5ded5b1e67271c66560310f71fd899c5442b3d7e58b53f92b83b372a3c033e3154c5126f419ea78c63de4755a6209fdb13dfa152e150c66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb28c9b380825b1a5b776f95fb8cbc1ba2343dca377ea3d1f24057220245e5a781f501aa31b48a82e439ce2e184413d7bc0f25b2083e9536d7d71288ed77970d7413b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16bb89a64a8f30c5235dc047e23e1d799dffbf7c489ed2837abb4aef9ad7a1b9b4458fcae56b260f273c89f5926cc648f13e50320aca7144285c6e31da28ec5274f81;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad06018e23efb3a7d598992f04ae350544d6299507f93bb6d46071acf7b95ac5ea45910b9557b6daa94f89708b611fe604ab7ffe872d6ab20c65f7095ee2cf855e5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13368cde347da80e97e4f4111f5971a559a6e9b0073ce966dd9cb3568cfb38f38c26ffcdd112508d5914794279593a09994a16a10915bcbde8d7bd7843fef577e9467;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1766b8511d5a1b0c1f69be21f2544eb746b6cae26a4cdbd7f93120188bd4c6afe0dc2cb20b35ca83c6346c5690d63fe817acc0f893db4e3ba918831e32ce70b819527;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f63b9e7d84ad795a3e6afadbcff77aea018be5949c9e0fc34ec36748248576818eb99cedc15f33c4773e14b3a264147ca95a0ffe54a3aad021dcd40dc85d4fbcb83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3857233c4765fde41c6e748191b56f56892932961734b1f89e235d4466637e4e16790805bb9275a2f40de94ee1bd57b0b78c30e007dca20623442a99bac6aa5c5357;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0f6583cb057276d1f8cda10b959112bb5db53477ab59772c5afce310fd7d85f1b5df6d12fbdd9f6e6abd9af82a8dff5f2b9838fa54e074c120ea47e325cc6178b04;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1216418e9c5f3fc37fcdd7233ed160acc25d5e9e59e57a01f3acebbac039b68e9d9eb3794c98da39484fabe9d9e954fe22c9a16e6d1c52685dff81e9b17d6b84e4115;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6adb6bde5ce0bacea09ccb93cc080bb9c153aa114afb7ab356e807226f14732f343602a58006e76914ff38b19a0691642d435939d0a8c12ec86acdff15473c5c135b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a906dd8aa5906e1401265e3aba5cbf4353e64347e07add96a53410050bdf0decd17bf3e6e6c2e3d0f27403c4f2bbf9a943f7eaeb7e5d5a728a40c062a7d82702cb8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h75efd6d0475418e41f64f102d80a67da99b641c94bb1b80ac1eb60679f287aac933cef8942f8c4bf5471094de581cdd05ee19441252f127b20972da7e585ef397ba5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d2f2f4bc4f542c262c77b9ee9bd71396f3e45c15ab9da940e722819d827200d7f3b3eca0bdeb87666d8f9eaf1c1c758ff097254ea4480948f30092d03c0dc22e257b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha033da84ccc82120718d268bdd807f3a128ca07557bcace5d2328ccc4cf370188a07b5cfd3a4e1ca35dc6a6bcfcaaa3011231c9b166e0ed3bb92e839462b7bea91b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc9d4e4f6b56289877f1493877c6aae1e68eae2e6a5fa85e02b94eca774f4a3db617afdc074105dece702ed6ee49e22b57c2ecd0fd50da907e201c25c857df3e5406;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a653de80b20a1779308fc12f4ef980edc84c5305da0a2159b342a7f10197c5a324c74037e9446323901d27ccf4aa5bada012567178e3552d2d3c059cf14192dc7a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e79d20ccdad3c315b5a2a4a6a0d3d6379c1d46734d2c8f8ebc1217c8a92751c5f32fa2787fef38f745354a04cd9c1aa06cc668fd8685b37c405d095056639b39697;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60576d5b97de116d106ca13b543d00897872ec972d14c8316855309548209984982136f504c98749e1d625a8a34e5328d878339fdff439722e65c8d38d08732ad448;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12716538b21a18010ff606ce6928a764fdfd2e70142ed73971df7166e81a5b3af59aa1b4cb04105b32d8dc31a28a750833a5175e5171435d7bcdaff2d5df02e48d202;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e6e4e84387c11093d395faf2b3383a087521a8277dc8b9b02d0e371eff6948d1c802d61201c2f1cdf9cd442b7d003e47e1ed8181cb5fc1b58db14aac372efa88f8d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12e7282c03a7f15f2081248e465c7e51d2c179bab89d86fa4d5eb51c160e9ef5997ed6b1e2e4ac48816a10075efa5618b7e86eac1bb97fc568ce163f70e0020d6b129;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5aafcc9fb353bb3d68ee3edd12c1c32057326989dc6ff5b5996b87a28c474520f3aea323352bcefe5cbc8663ce3e740133bfcfb164ced586b7bd1eef88f69f9db484;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hec69b92541c44f7b090c78e2415a62e43e5054eba2209f1ba8b6a2664cdd344a5f22cda38a197fd1b34daf71e50a731f70b3d6a17ef26c6334b3ce235036bcaf01ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb5b6161e708b0c78e7887177cff551317ddac2c24fe79a35f26adb9aa65520c3096ad05f5e9ca6e6bcb63d45e2207f4bc734a4d9728bfdee49626d6cbb18bf21f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h188deca6c7b2507c6f3da97feafd8ecc8db98045bdccfcbd183be498653a38a9645af4e0f0a967146066e10834e7afe2fe36a58dd65cd030198a471e554d1884acfa8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcea9d2374b0589b308cf71ed7293a83846293c9b8d644d2d1b8c5cb546ced8b40d77abbcf4cc1ef4871545ceb26e5a377757446a19139e986ffb4cefef23dd9612f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha2b4cd167c6ff43b5d59b397302951f75102c1e00355323c06a620da00f1e3ee48c637b43ed712e8252af6effba738ccd9ae261f0863f222a0ee5c9b2d088a26a2c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfbe30fd4d21640a84b5f644b391bc0ce9d5b8354e8c51795b22d690b151f8ac003441727653dadeca84a39935323c7c2fd7d9873cad02138d31d2f50c56a5cb78ccb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3eb645af477f6c38b5238ef27b83c4d70bf157749b8c782f10c6e64503a9e8db54a15110a41c60daad5db12447f957fb269c55fdc35794d961f647b7592716c58a50;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heaab512fd4568f62fa2394ed34815a429d50b5185a0d3f942a9cd6f7b522b4643be53138ea1b944fa63fff0e8a871daf4f85dd7b9341e21bead4a944c41c9b5e3588;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d2c9a52bbb38cb5d4c965e00a82ac5daddfc2b075e4f9a194166cf76e0cf5021eba10a78af7ae8b6a86feff3cdba843798e8a327ac698de2f93a242ed2eaef2f5d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h858374c47184158d55084ab3b93589dcb9e9412245ac101c2548084db5b6feea68a4b6f59d3fe986a4e2ec7dffb138818e4caa73e589bab6415396a7ad12bdea8dbe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1102880fdfa264972ce0233f32bbf95b2a5d863f21850932b8776bf2226b1956ac1a0619e86da4e44b36fc9907d6b133e70b0c9b8d135f57ea367d2267e921af879ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a45bfd9f82cc19ba26b39f26f8adf8e4f4b4723fff2ff37d067580adeda593da9584293b0b5a84e9c07ac0b6ac662fe94e4bbadf25170a4ff43806283e0c71f7ad94;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8662b3fc66a981daa52945f4b232e67fdb6d8a48c19a155245f1709910b467757d255d1f393fa125d9eab0e647f227d5f38e544ef90c6b2347ff456077087e147032;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19f65d1d3eb0c5d82f21af6d276adfd27e3153f81023c86e81317607a75a0e983fe28a7c65e7132b9c931c658b7c54624b9882fb021c603473ff907b333e32b2c75e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16915f2ee6b92b1dd0c61e3b289f1b44f9efc41ea3a22032f6e979f55c2f0cd32d05746ecdb88bf00dd40257b45de07ed0fce1f0ef903e80d4a492d158305c04e9039;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1462cbf20042faf125407b98d8c688b02e978a5bb41ab5530adfcf5b2d161198260d1adbe909b4b05934d94137ee57f8777d5a53f4317a4bad79cc973ac34e0321986;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a83d9eaf912c96d471e42afbcec882bb0a6c08614e229187aec3fdb8580c1b72ec8370f7d19a9e7528993521171f0f2807de6c27582482252e9a18b0f2255efc3b8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f18d8d89b6382496bedea6e70fb75bea65ded0c858fa18686253b017cc4b6319c77602c9df21bd04f9151fe116aec33fb553dbe6d52b3a2d01ab8ae56b359341651;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h55cfa1b6cb2a6dcd67d674532847d433c670eae00a8f161387ed6d2d1579b2f28efdafb6fbce58847ca737a6258514ea5c30d01f9652774ee3c988dd3430f92831d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c342a47a8c8ce6612157a4966c3e505ee6ae1023e6969b63305596b04d0dfe8f9ecdcf231359263d2f8a71b2b7bc24a8064952f95f264863e2e8d1cae5f9ea138a25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7ed86a2939610753af0e94360d822eafcd222374fea7debb36d8561f7abb50160bff11b17f86d75bc120a9d5aeb7738199035c0debfc4665d30c0384dd5e42aa049;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120c03bcd20ca4eea0e90588d3b15faa1b84eed612250b7f9e4d74ea5cb51103947ae8a89325a7df609390b26781a76f5dbd80deda7589c3b26c6198be0ae0df28538;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d1f9c0afe7c1bd4e9a934393de425949f9fb29374c82b6e752fdb78f90ef9ff0fe810cb1553f7d98c3c70cd343be142894ce38b883b7095795716417f5d49c7a8d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14e77b68f29696786850361fc38608893085fe8cb374ece36aeadb7c04f26a706085e0c8e32f9ef6ac3255b6adc0ffdccbd676a3e7add0b413acc3cbf3ab9aa6ad2d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13daa00dafd1f53ba8352baf5842726cc723301350ca75b6d2e78fb7e33467ec092ca6051bec19bf11450b854d037945e0635478bd3abc15a47d85b7829d61f1faa22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18139e24cb140dbb7e655752d69534ababcf389a069cf2a3ff36ea9ea64ee7817f2b0ff3adc813a33709c526f1e1fd42545de830b5fe0e063dee8cb6af442cd10ba5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198ea15be6576ec300d2052cc731b79cb1ba5ae95c8d0ecb46ec293811ff3739b5ad8514f3e9ca041b55d1b237d45db507160a329c6ff82b875ec9b02efcf2ffb373;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11928e5e1b8648ff732b4e64bbb8d169552cd3795d04e352a460cc687366b0904594fef2bf8adcd2d9794189cf197f321752241cb96fadbf9745c8bcae5d8d04a4d3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h68f8025c93f1aea6a67c014ea238fc2458d2bc00d5f6834f4e617c57bda1d29af47bfc76e5239f351a5fa82f171d559030dbe9de48cfdaf1deebcf17289781bf1c2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h201953c19769ffd5ab981bb8d3f3f8969631b4a189b18ce4e2234dc8522901685168f0366a85183f8efff26f03dc41e7dceac86ffe18c81e0575564bb9c907fd6b40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd501dc4465360ab7c4f57b32f20458cf34d6c3bf6488094da49b16c11b630eba188a2968a401d388f76846c5889c92e1ef95be7af3a2563465869110c9a47a23d4ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h140f5e2da9a694b11355bd72b943e59ed1d1afb715c481f712980d829b21336bc10f4c67d6d4559a230430e14507a5d43759b48f5eda7603e1e9b93b22135368a0811;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2fb958bbc90191ef79250b40e719e1240b28927eb194d5ab59b765dee0242f4339e2fe3044410239506d613a6885a24f9877f636e6b483cbbbab58b1c49674558aa1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hee287e2872b0a15e92d7e992c2a00615c4a1d73b1305e4315f36be851b3846c954f83d09cae34b70c9b162fa754a6d8afc70a556c2a1ef81244876f4aee6dabe103;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19401d0c624297f7c443c2a416ccdd53439d9f6c9a87fea8b7160a81b122066f593972a8ef18083526e6a58f9cfb91ad69b5a3fc966eb919966bdb59cc5676ee45791;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16846ff5abe0ffbfc61355364c90cfee435b94be55be7db4310daaef9585dce95741d0dc74884df87c32287d04ef8abe107090b8b371a6a0a8f4f49083ef62cd4365;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h41864f026140732c738a76fbe03caf9b3f5875bb214f4153867a2585968969002a89b3eb299db85ab10f3b19bfda52724fe4d808b9918226f300799e3df7590ed831;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d59b4aa6b0678296885af2b207bf383c1889818d564142d18b6a369f66b895a04640b61770d4d237e04cbba55579af02728638c4a5ae348914da6452063948e5c3f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e8bad9d03625fa57bc7877bc187fafd6eac321a93d6f8f84c8ec74bc45d963a390b55977ee6c278f53df3bc7cf34c58d9a58b9ccc4ca2aca9a45435d72b59ffd6313;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121045eca383b3ddb6832bda81f54fbafcf318716c423eccfd527b1d542456cee00a7832836034859c07e2da7dd5b95acdc751e0d6734772f575393083b9d2c6156ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f2d945525873cd1ba1dc7c1896b898b9e28202f4f9bdfd6487bbef61b91826bc4c73eabe7bc6ad48de140113ccd12ebce22f13e32d78c79d74a3e9092bd78b5b9d2c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h176ca1265b9dcdc9dc7f178005f8f5fee483eb83eeceadd7f6afd275b250e10871b8bd34b75726312a0da8ae5c1292a458a77a940a0f6c9ccbddf0cdc4677e076df94;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d037722cfbe4e79cbe623d4b08f01e647582306a596694985ce638955ca69d980721523c32143d60a739cf890b26e8d6dc24eb3d170231f5ebc263291f173172802b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac096ce2fd27ac249b38ce7ab8f1656422ae98baed0fe041f4bac869d25893dd10571d61296f441b2383b70b7e3276eae032eb9e06f37fa34138024734d395d58f1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a7a213a3c4e79eb680e6697505623edd05a7fe9cb0891e5608e0786fab90deae266828adb403fbf2d960f128e45dfa759a99d9b986a98abe7802ab40a177417e4bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16914dacfceefa4df7edcdc80d67339726eb2630cd2e480f53c2a3d1c2084b9897876d30a3f55479b3227ac299deb6f70f782b52879ef56625ba545f86767f261b0f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h76fff87e65c927ca55f0b8ea39bfebc6cb7e64efbdea78b3af20fef4b542eeab2fd9f76c0fc7f4a63e9e2076af36734ec39b6024e473781f228ca2e42f3c89d792d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d5906a293bc373f3081ea9cf8b8c0bd3d9fba9ccdd645ca11041f483c189859d32a464c0b41911b96ea17d2ce73957c5acbac22988714bf67182a6e6974f9481c3e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a79255401d299f4a941a9cf98bf6ccb06168c6166d89cb549c02239871a32446bf23ed6ff04947202a71431a144ac02da4030ccfcdf40191d426b80f886d9a3b576d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14c1935ff647f46bee9fa718fbead61337b6da6835a5332bae388e777229d53214d6b6f4326230e05ccb1ea2153e3bad6bb79af96577282ea19d8fd3d0a2e5d6cf8f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf5b9e8c1cd459aa0178d5cd98cacba78bd52c3634d3cc07ac19b94348bf9d1abf76efaa527641cb317ecdd8917d38f39094eab71318e3c1e59c490554a9b119b38ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5022f722440ec9c4e13807c251183e3f80b219f067b155e01d329d1df99b43f1dcd84a3a6e109171c515b98bf04423fdef2863d1a7fadd37e14207dfe02fa1ac60f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a0f9bae95150530084317b57e51814a0582cc186ce3ac980a34c0f4256a54dec7cab468c9ad4034e1d2a9d0c7496b67b79e11a9212dfffc607edfd69a11a96fc8c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h321943672e36a9d0adbbed1f0f89984b91416fa4ae678ebff01e02ebb030e76b8da6bea10c487a164059bcf5492409fb7f63fc0da8fc494243a83f949ff4ffaacade;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h87e73bc1f3b7348cdb577461fb0bee58ef560af7e9140b48d1859aa1aa3f861c7cce04cbaf1abb255c7731cc2fb1873d6726c1fabe468038762aa264b00c99f53d4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17210d5f81e05b71be37b8bb2787bbc26a53250c6e79b4930ec6ccf0a7f8fff9e2a6a1e51e56debc16533a8f1b4992c597411e58d9e0129f65ce9a36f393c743a742e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c8970e1f03e070db2855291bb8291b0ae6175bf8c7967e29dd6a9333aeb5818503141d7c135e7d576bb4ef818640db5b7ab060e82b4fcf6d663841688f7287f5175;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1831ef4bae4aa8d2e4f993fc305f129566f4d9a92b10903d33e55c8b2954368816b319d501c6dd6e7782aa3b3977f121101fb0a5c88aaf78e1bfea6c4a15956e84c23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180702dccd6975602bdd6f732ab2ac7ddb545ba48e07ce71a62813dc0ac9ae61d5463e826e54b49d8f4e057fcbcb6f2c949a5b5ae3c7cb2cf7427ef85dec0bb10e378;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h130b8782e21e95bf09e9300fdff2158f3348416de9715e272fd012d4b77ba6df9e3edf0e396eb7b1ab0cd7020d6c52cb25a5995189325ed929a3087f4480e3bd20f01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d32558985f5f8a0f2f6541c3c80f6df7e2484ec99366f707560ce3cd5c7db03cbebe8724f19f71ecc56db26295fc7709103f3c4d262259db038837e9b0eba4a2f849;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf2a31855f073e5c156b073b24ee1e412271d393b3d7996811d4ca89ca18e1fa7e47c191b0c4cf95d22931d081687a1a5059ec454c1ff94a6f6b281465fd26855235d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101c60bd27717113657f1104f8802c7991819d20db66e93fffac95ef067c482e96d1caa28320c61d796ff87f21bb01744e35772b1731fd63926208914553cd3e54ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f56e0494c1a573ca13227ff55fe70b368d8066f4a33cf8d03e99908d6848cbdfc9d4548118b4bf2642bc7e9f382a11c0720b60ec38a2aebe92b0f22e9416b3d1a3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h877558268d826edc54e3fcee62ca9196e7c5578a09e87c879a3c1faed376801cedcda0f2735ed748e7bb56d7305981402d5fe83ca679d990be10ead322d405dfe26b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h998affa6a3a8a36f851311385cf6e07e82acd764c3714096858b7987e2439cf2564c997cf0534759e44862a549fac456ce957621be2097cc8e7f9ed6d70dbbb8759b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1db63874b2c2771e69325a525cdc93b5c1e1a90fc78619d7be0047105007a70686d1baf9da19babe81f9edffd41c23d373b018c98d46e819f2d33457c106c3e65c616;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c156d03f6b67519f6814f593a90316fdeb10e1cfbf8107d425d4d37e3ea6c9643aae8d234a902307d5722c42a94ebf90aa0bd51ca65a0bb58185c4247ae450a9fe23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14154d0501bf1925c20876e0e2d11da6b415a562162d331cfa3330390864615e82a611c74e5c58d323e5457cb21fc2a99289c73ee18937bee4c8b9b01560c36acedf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17220c9967649220c5cf2f4a9aa13646f31cac85b559959185e5526737681aba029c9881031c76860f7b991ddc379007051ff4d209ef7d7ee278ba332785c3b22bdae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71c3f79c1748d7b29ff1815f7cfb7920d0175dff5dc03e4fcf43ef519a18533ffef0fc19f78a5fdee7a738d915f98c7bce55b308e4b4e2c7bb71834ece54cb77b65d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18eec386fd1288d8d1b5c8b480a6281fbf7a4a679d7cde0ceaef8010e7abac43ca72269f25d594724ec36de3a2349ad090bab670cf4a0ae0dcd761e7f961b95fe5a78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f11a4e0aa2080aa61314c6606b6dac5cca4e5cd41a21353917135ada06a6ed399ac82b079a05368f0300c2197db51dd27a782d04a246ef7b611bcd3392a2f01731b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf008a5ee77c2e69f3ac6c2f5f94e7cc8000d71042faddd897a4ba713410064e2d7c1c76637971f2c7866dd91e7a5d7993bec928ec4ba5e42e8808deae3fdf35d1f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4f18b010ab06b55c7d8f14122281ae7a391f5ba2a59bf9b8c4309cba0ae0e90dacad7c2c5c0d0dfc66578fd73a8b36dcb9d4c0a1fc18620a4eb76d50fbd71c504b64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7baa68c9a8afe1defcca26f3ae85966faa0cfdcf8aa558059e210cfc4986743184929b36f85b6b080e737caa345ff89ef6402c00e21025a2e557d65c602377c05f4b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h114f651bbe1d773250d7ed3461764b77266ac182c8a877736b86342ffae06e6a68fce7b6640828ab3a207640c31a9d4b5bf673e6b1414d003e231c722613b5323905d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9891824a6f914874c50c08a76759174504c01f0f99c5c7554ef1671208310fa68dc823fae99c561c544ea6d85a30cc9eb630344fb253de664981fc0c75ba6372c50;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1299cd09679bb376d269f266c033232983512b6676b2213fae4c79c677efd7f28abd378a092d2a2aa0038d94d3c2aec80b6d3888a3562923ccecb8b2c24ff05bc8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h99bcb5c12210b6f03c7cd0917043181237af38640480c95d4000c32abaa630cd932e0de4efbcac468f744ab40881bffe6cfc311f66f68f9fe964083233b748afd44f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf68c5a61f63a02b1386e5aa2beebcf27b49882900b3db1f50eab1d1b4c306b213d998b8b30a4cff38891ae5aa90a30b22b2423da2f798eaa8c39058548ebf0faa8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d784dce4e3e6fb96e890e8fa6596ecfd18d49632359b4023e8d9b7fe72d607b4cc2ddb4a7e7dcf0d88957081398461d437c175602dd9ef46aa369ed071d4e958692;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f959dbdda305b3a40d75ea69b80f9d757c75c12d10e07cff129ff52b620fcb23b9529d82e633f0339a2fba8883b0e545818f4a4750ef40fca9f3e5e387a2c174c475;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af29a09e7003853963efaa72e6ed712e698da4646e1668da99f23e0eae32e4d5cd02ff849a4e6b7e511f3556e49f8745d3ec69416dbd89e83076bb78c3df30ba13f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10aa7e0d2cdc5ad1e4a730b1274229e3a250e79238e5738e9460eeeaf4b5c663f8c1e66fea4dadfd0d2c629b32668f524d443e83a5fd34e16ea34b6d7733cc456ca7a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1034f1f1421ce63126be3196a22c3cec8c0eed3d974659c8d9998b0979becc4068254f14c47e91274b2204dc9bfb60ddae03c31ccb37c6cbd4c1d308d485904eeccd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h29f817159009f1bcdb6843e83026e1d4ca0a9a53db7cb537a5c16b63fb4bb71079d0d2af86734102cba8456a375c859fd5db26e14cc076ac9b954962138288d10304;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab4f900743c96b339dc447d962bec150a062c2d9c42306587c046339aeff45bd83eb4e109a48e6aba6bb925cbf862fe9688a03669817ecf453f14222ffc785dff927;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a8206bd8e3fba74c3ac2c6dd2550cb8cbaff8cdf5fca12253c275b8bde3a655cdc1e132282d50804f30849f3e4221318252f0b74bee16a3b537b4d902f07da88529;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c3f1587c82ee07b9b22aaee6e4a59fbb2c8dd78a2a4be8f36ebccd5d003afd293a34b0bc9cf24a5a63e16cae479e63db5c39780c6a71c0213ae892992ca32a8f2c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19f8b1dc7cee95aa9817067b2ba67f94f48ee6beadd7daf033f5966e0265c8729795c55ebfbbac35ba7fdd67c896ace62a2800c821b1b0dde7a26ad07d7ba418b4449;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da6e13a04c7a1dff1f07563613c35281f38fab876969187d70cda8c7e7540bc79cc178002e8ca1694395267fae7a83d279888345c6712f9e89371af9320bab73b5c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffb24987f3adcafbbabb1ab82607ef7d34d23971eb0bef1b163109ee5c5e61c051dad6a04f0bb335f0923cf663a895b6a3954ec1bbb4d0dbb184cf5a2d8f7b128d05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb20909a33fe944b3b12dda9dd36179ca576e2bc66eced7178077933bc642e3305ce421500574e8cfb16d485a88398dd25342882a1b62657935d65711f416c27caea6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12440f8a3bbe4508fa9ef9d35391072006fcebf1865b20dc7a0c411cd11887b27e565eb0758bca1ad00f3f1804c7980e1d26263133e3e06ca179e25a04c218809ced0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c0b2d4364288c86a2464c7371d03782381c7b2a07110a61016899890d9a83fde3bfa07daa9c04e2e1d22902858c65c9958358ef3591d7f7f0ad0f80a2e9b8ca2d7ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b702465795dabaaa30b75e7f70c9785cc93260dde7f448c7ff0fcd57ce7c2f4fe841b357031d7b3679bf27c99134fd0fe72aa686553ca345f302df39de27d4e2bd10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14f81cac96a846d6dd11155968bc7988180a217b91cbbac2d7a96abf40b0a1afbce119d0822fb30e6fb5811a0c3b66ff4e8d0dc05a722f2a45841a3a889907e604a5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e37d70132e3d76922c3362dc2258bb8427fe15c6be5149c4e523b28274ff9677093fed5aaa3e5cfb1ad5f58036f9c5170699252218b6c19e64c51f1e3d228eba5d38;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91f9ce1f1d6eb5f96cc10c6831bdf0ae18ed52a3321d2196fbc6bac39d3131222fa488281fe2fca940ca2fad7df01201554784b5a21c4cc4947e3349c67abad41058;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bca06568f1892784637239e8a158e66de6651823e396df734d29b71f3d72fd860409e5fb5646f3b0315af7169e9d2c0a02bb619283c1a066dcf82999b01d6c5bade;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h819b8816d77d15ad1a1dc0c29961562f2ba53ac8c83d32dd684719c02a1c56d844d32f9fc5005c0b31543afff6698398cc6f90cae1439bdf6c2fbee115f3ed32b08b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b6405aca68f0a8e6f24863feb476c0d6bda0ba07dffe71754d1691e58c4cbc514f1d3cf20c5d95760cb291fcc650aea53f2ca954bcd3c867d530e88d576db8693b56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d76f0930e2146e41a0ee55bb144f8ceee892c9a47cc9882a248ceb45093a392fa5325ced0b6685b9c5e1aaf51d5afc2ce6015f7758c630ff590a7ac22cacc71c72c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b26574de070f0b4e362922e34c1d579a71fb9ca73e0ed41b91db339d18b1f9cbf0ea471d301e58f4d70bbf3f5274fc4904c6431248015e5591d82ea28e712deb0211;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9ef158db55f1b5ebec17e4b59bfeb8a51d6c3f8865290aa8e1bced182baa8f7a4532a58383feede642baf9add8157446f4011fa51b3578f7faa4f81c1c1dc0f15ab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb8f6db4b33bb844baf14f00907de4403f102ba7fa8bd2f9fedda6bfc313eb8854a673fdaf900a72b7a348bbbc57e7da2b3ad7075467e718b71422c8e8c7a76d30d0a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h181fe453e5fd9d703e85717bcda96c7df4a69604827a2c7dda8d7e5aa22de38a66b17aebe01a7bd265fc49ec6bb165bc2e06d080fd9ab99de4d2ca40b9d82949a1bee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b6080579c1eca0c745dc9fd5dec0112b304bb82cd2254c800a7212d3a4ca1d4ddf87bcaad7dbb927560088fb30189a5910dd4771fae96052ad990663f716e4c4a795;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha47b805d750cf8991fe028b2c8bf8f29598d13c4b338c15086bf2140b4e170138b09f8d3e365fbfdcb2f2cefa55895d2fc0f12f3dfb9304dcf9ef266983977af11f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd4a7cc8b36e2b25ef7359da9a2ad8452867f36fb005da8a4940020fb917daba0c96a910f25c5f071d4e62a88c6be73d35ec7506212a713e83896d26e6030d34c6c9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d8988b39776936e5e0eacec3e8645b398144c767dbd0bcea42a230a8c06142e0a12852eb5cd59ef29d54def1204998858152843287dd44491dd3551e23d03e4601b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c363c2d3d223a55734faf4a52546ce175b15028f9a32a7d1de430505bafc1a7a30ced60685b6ea0f6504243446e1e76303bdc8b1a69692bd346aa88e19019b4b5d9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108c19a121d6693755c32c9879c4e35f04c372667fd21c477d7d6cd2d77081b07ea1725853007b8649227518b38d3fc25408e5e7d86c1820b424435f11016f936c60d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b8ce20f4e6d3775d27d9b9ef68a9a21e43bf8d3278c0e0fcd34e745172fba8188dc053c128ca28c2d07a69cacd5bbba661f8c6d98c1cfca172a0ff50abdbf22215e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17832aaf13ffcf67a82f16e27474c80fe16015c49dbc12f8525c1a75a27e83b3a1d8c480db3d62e57b744658d0b4af4518acba46bf33b7fccb283c80337287b3b06f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13515ee5fc400b04d7a1b6effbebce9e980e64932f8c226a5b697a682f89a375447ae18c0e34471a4a77c93d1e0c6a4f8db749d03e89e6680359b0fa4caa57f7ee1bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d663c7dcb8a53487683fdb46743b1a1f4488cd9cfb9769b4bd6929b747b8ff438e1a577f5f0d7052870ff2487374021c8dfae1b1f88aba87584818d514d9d0f519a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fda7e00d17786e916fb3531bb5e2cf0027e74f4fb8fdb839b1b8f194ac27475855edcca6501831e9363d1a5830617d5b3aef37dc8ff3625916fc59bdba53711f7e84;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbed58c589f4a29646367f07419c250f21191716d703f1db3921bc653d3373fa94f055e97c179f8d717ad2bcd9402f5b235c9541ff1c83d6f5f7fe57ee1c2c20ca143;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1abe255fafccdfa980dd22dcae6823d382631d2439992ee5856d6258da7f58ae9f1c909db93bc9ecfb433e30275a7a0786a744a2c9da4138c6cec49c0ee0c4246511f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a7a4f56904009c361d23dd11e428b48808f4da91cec26a72dbfa7ef511f1a4f7b2bd3a83ba320198e93a588d1948252b7ec5f32b1d92a6fe27bd9d7e7f9c351dc06d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b07515a8150ac799a3fb1d024184581580b430a0d2c0df0f920b6823e3c7b4a60aa98a6310a00c726ea18194475810f7c37a66719819aa45a9439797032de0bf790;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h164eda11f37fa044e087fa4817869ed5a7e524a669953d498dccb4fe5cafbdfff6451b5dc94cd4fc7db2fb79fe8ccce1b9f6d83b3796200244b0470315275d6cc32c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9cc7df11a0f3ae9905a6cec443e823f69c86be4e485bec943ace5d626ea5c0fef9bca70691ce5ccd2a46b593290ff66eec72f67f58e4372672f511d1e54ae6b0c9c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c63c64c50145333bcd81821eadd04cd465cef99c8e87d6a07ed61eaa5c131ab4bff7216a110e0fe4929f97023fd8e0635ccb988b0da003f4e12e58648a1759523732;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h567947d09261f3bc7cb9a57c9afb04c01fb038783cd222292ae0070a4adb989a76a343740486e990bca9e8ab9aa2cf4f8092dd90d777788118e7f3c88d8537799839;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc326ae3f492832d9415a88d9ac37bf40581a4fe848a7e55b227d83d29ec105a4557eb1b5c0d6eaebb75d6dadfda7d71bec7683070add673e900a028f4ab5397e2a2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb592d18dd23c398d147c002f8f11bf530a83951b93ed8aa9c6e79b0b925c7f3b619abb417ad787d125a7bb97cbe24670e7c8af63df2e94fef7325fe8fe03ec611dbc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c241141f304c84b19b9ea783a290063c13a574133b26c65af2e7c386ee526e489b36d8fcba61f7c5a5534094eb03e728d8640fcc8d56a340ee784a5162704e75f43c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb1238c5ffa2f38efca4a426768dc9128aff403984ed96ee43b76c1464e8ca6d00dd076345ff44671e21a22c7867e5a49d3536a8d61685684fedf241f22e1042a4d18;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f7e3b9bdd91424fdaff7f21a8b14cb4025578d3313a285f2f4679e178d67c7bba31183404ee25d3eac0573e192a0d33240a834a2de1bd073decfd176d52378397e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4bbbf60d7ffdaed8d126ea7ce937b33dbd863df52bde3c01566a659f4a18c69ad944f967120e9faa573551cf2ee69f8a00443f79b1275a7355f5772a3210e77437a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aae4bbae446a6edb098819ee33c0899f5e05da15b93c432af0e4c7ffce5cfd8c60f74f7c6211154526437e77f1e3443b3c485d370169f0d4e08802ff20996a41420;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a5d15bf6c85afd12838a1a75a96485eaf373e27a9023bc6b417d8670b6140e7e0fb8d7b90755c6d089f8e995abc3286b43a59d7ac868f93c5f98ca5d723334659464;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6755808ef46944e1cfa648ab371d22cba74d2f653bf592b92f1232bb14f18a9eae0a1791bf2cca0b27aa9b0a83dc3d02f0b9037d677ea93d8f3e180bdcacd3f23018;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c39cbc51e4415fbc2acc8b5cb1d5e287201a42e1f7c692bebd61021c5baea39e022075b2e29a3aa8b594b34ccf60ce934d1b996dadab6a3001092d3a7819560c71ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha36d73274fd3d0c7e79f74f74ee5b8566df8e8aa2c714b07d618f38ab6e4ffc10be8a0bb82fb92f169bfb963c24778583772921e1c650dd0ee3c041a272634a20827;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a3821a712b81e11eaa679f2f880c02234f22cf42c2fc2fd5a0c3bdbbfb1beba0ad9fb56d7aec668dc483f2f19746fdc12f2e6c243e2a65987aa5598901c74f0c1ad4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3972ef882377ef8a302e6aaf1e80ffbf3f90816946beeaad31d8917838d603c1a1f3dda0830db82582792385804420f134208094defeb288d58e26c71d66f9817cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h830e44d4247bce472018fae5752ab0f49889e8d3c55f2478ed82ffa90e96d530e44b48be4fbd2cef4e3359ddfaafc975acdbb6860d0578a5fe4e9f8d663de5b12773;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h72999b24ae46c1cd0c87e6bfb8eb4dde8e995837404da524c1ac9bb299f819f17fb73f0cab9109ad921e7c2ddefeb96c7b7e1993ec29f85d049237dd4bef726dc05e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b4bfc99af88b20d6a4862a2553e05d3d75f3a68928a09f9f44d63c2fd5b54d404fc02a8d49989b462e297cc41becae340ba61d95026c829b94968e772c72a436db02;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e2d50163d800dd60aab39e4e367d54f11975b8ceb1a74990adf9d52f484632e64d8c3deaebc54ebd232d946b4b4480de0e151ab39ae232d3962ada96adee2d7ede6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc019a26aa1f156dbe4d056f827fee826f36679275f78e765f645590400d5b63caa949c4b21ac8884be84b01c553045d46a348eb55244b39192bd798daf642535094;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haef43e163248f3669ccc8743712253eacc4d5d32a24ea3ec749804e9417c8d1f655a13ba811c21577336ce0a95eed41a306ffd94d06d09b7c62a0352d7c72cf7bc5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h95a623f438cff87a649bf7d238c387b04b0600a45ac1b37112b3488ca423a26214a807eb303ea53073cd3ad5f089b746ac117929fab62ff84a2bbd974c7053ef8eb1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17297fa21431266e7412ede6edd990d3bbfb5b917cbc5f45af692114853b2e0cb7fef773b272e12187f316e8c3b2106f5f67a14ba536640089d6945bf1129c704e8ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h626bc46cca56e44806b398e85f633315f95da47f65364306c108b1f63ee055a3e3580edbe70d59075d66c1687545849b933aee345883d8aeaf34eb5263673c1a4270;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6977a19d0b8171faa9e6849a1950df685fa2f20996e7f073c4df37814e047b24d676904622c4008f93b1e7e6661b19f68c58dd76115d09a1121e64a9081af49fef73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c18fab4f2fc97376f669e41df4d9805f61a0da5e554318d1da1f9c40a58ba9c6586b76b14338eecd0d8eb5de6192e373e273a3c4ba93380b74d885b05c6c816b6427;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h106d405d4d70e5a4631b7470bf18a2584d856a13a58c9fd0a5b15534b0003698e73c7f7e6918c461f0d920948e45c4d39e80de6945f9aa8f5bf2f1e03034740ab170c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1938bc71c10d710af437c4e59d43bf4852624991b74b4c7ad9f263ed2f479b62ea3d77ddf7d05dabfc859829d738846b05e69a0610f52fa34c26b67883477e049f40b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0c730f9b8074985561e23746be0761736fe301a79237031c26781e332903e2bcffa6d5916132789dd2459ee7f4dc01be7133d5c15341d18377d2c2c3a18a3a61873;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha91ea2b9aacbc1f3c97159981382b08e0ec269fea45e8722d2ab625b029451212f4c0d2ba14ae2087862fefb75865ca875203cd3dd9265ab808f93f27548a471c810;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61341d604fc16414362f12938aad5fee5f6e2cf814e82a2f5173629ebd6987649c3a1fa416495bb1d81aef1ffdaa5ba5cdccd4f70fff0487ea840090c1227356350d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f56be82442448845a20ab52116b9aca99ddae4c03c1ac7aa0eff30e28bc2398032487049ce51ff11cab42649eb93ef1b692da94dd0968fdd1bc84a4e1df39afa356;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4360aa8bc97fe73de1c3e8829821127634bcc459b218dbe27a25bd3b9dca86df0f7cad1a92d9a7ac01bfdbb304be29d3d339cf05560f67ab56d78bd0aff6aba8f498;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc883b15f4a154a7c210eccfd1319313889edd3ad0097aa3b0971d4a85ba80f7b21fcec983cd1a9cb6eb42afa30d205caf128125e4165e1607134b0bf6527f7b810d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b99efb1d390dc99ae34bd7e185b5534c0abee004be3e697c4949b6759b845038cb40ac91ffcab6456d550ddf9595235ab8f37ffb1262023dc062d982bfce25a43e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb52045e7ad8c1fce9d421b3a3a8ca13b84856d9d0cb31555379d3334dfc2404c0b3b544ebc7901a4cc91995bf097b277922860a5a6c9cae8f7f6e4a364defe5d3349;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4393a31963c13f34504cb953c4ba08c8fb8bc187d730593f375dced21977fdf7b37b2c70b281a744f4fbb2a935ced39b6f4ed1cdfd8355d5579851a453f78747265;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b245b576367586cfcbfff491a87296c91aa4d4936fcc531081115ec52bcbca72842814f02c641b2c91d12c17d73328609086be77aa339fbc8bcc9e4104c1b5783bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h94ae8cbf7b9fc7827350a4e896ef6e41e59853fac8f2426b2542e2448bda0c1201b31f732cc2e0efab463feea7d810d9464f885fc682faf4e81c3e2d333c87bfd67f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h235c44c48fdc2af9846d9270e47ccd26ca0e856b0011d92ac8b5b525eafe06fe3827b6e4c85ea3716c6650a9ed442847278d11f6481c150656467351e8ec911ba570;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h126decf08b1a607d9350a7c44066d3c7d26c8aba6c51ef24d756b1d32f86dc5a50b1e929d3d5c1382bb09c0e64443ed374065ecbf1cd04b6c0a618ac4029470c7d205;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b00917f6f87f933a8dc842bf9ea573823d0f96479a727116f71ef50c38cc73982072003f8bc4bac9bd945da81bbcd9ffa61c4e5b909a663da996b532f48f6b64619e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7765fa7ef02a6cf758af31c1ee09ccf25339f896ce90bb4c2f754791d4177ff03a67d670bfeec64582b0bcb66743cc2c18e4a62bad43df80fe05ff3436e707de43e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h25f546591ca8c34e5adb8311745cd58642e30651910e93313bfc617ad4d808fa20a28243e8da227a41dff5c27fe97772b2b5ec3d317a3d9adbe05f4c315286e68033;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19fd144c36ac3d3b3763344da6116a7b3b706606cd9c4d22f55e60b4d0817fba16edd20a686b7bd28e84ed80da676c922789d4e1e10d5af7ce2f445133903c2d0dcc6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1de623ea835ecf56f9e4ead2845b78173fdf057a61d35395dec0f12dda7b745ea2b3f3cc931b5d02c6e46ce232269b3b17f74fad8fc641fb418a07c00834e4b3927c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b575eb99aa9cdd3003f3f39d41990b532669963a4f522b9913a3fa5c38b769e0b226d7571c5e18433c156275b8aff241aeb9bdac6fcedb6c352e8149abab6e759a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d51e6c7f267f076f770cbee655a216a76c79632ccec64319b745ad748024dd2c3b2e0024e9e07e7534d5461184b2fe525d9b99c5301601b4de057cfb0199e534309;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12dccc6a98d47f407fc01983b4fb2459a3dc89b735f3cb8c4399ecddcab944b2507bf5b3223ed32ddf2f756c43b4fb5117570023e96987d427ebb0763cd27cf709cf7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha01c59a7abfac126e9b458a3bd8f46047ae28146887da04e8fde405e78f4fd9c66bbbabf5321b66e130d80fca08d363a9eac6003661bfa0c15ea5ebec6369a72743c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103eebf6f49e4084d6319f088f32d0e1ad313ef035fff8a2a8a6c2f8d55827f096e370537ecd106a034d43de0cebb4391aa17fdce5ede536db116a86e6ef31959d9bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1498612f0f4ee83bf7b36c9817a641bb432038b8fb0f68678f4d4490b259e4466361add5972bafdb47f419e430d217582a9166083c0e2643de6c03168d505299a5202;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121c8c0e1a1a2709acf93f8f33d1455b388a68b9778073002b3636be670d1dd42cd32b77d4195d1e22c80814a5d3a9541cf970c50a276de7135b943439c1ca43251f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc4e7d49860b388af6164ef8304d7bc4654dc57875cb3c1d2a9e22d35d1db491d94015550c280a99a8c8fe720d02cd66850b87fbe524a3282f24398febc4236ad468e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h192aa6a10c975df92f3a6298011f87f66553f75922575f5bd3c45ff22baebb1b1f7143e4a3935e4b2e4408200772c76f7ea3ec4f430535452444bff99d6adf8eca01b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1848b1bc2f01d93a67d07b5b6e115d55e184b6b0b4e331bdc61659b3d715652d785af2649178fe1ed8b7c023162010cdeebf6d92cd29da9f1a272324cb79dfc8ef938;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1641c92fa2b314cc1a7dd9f9f13b1372cfff745a59d4b821b0504d1faa6943e54ec4fd597d8ecf666b896797f45911ca781391901bdf4f772c83b8b0cd5d27de7087a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18805b433d4f8eb66ff7a5da4960f8c46704a3ab3880764aceb983c54d226379547d2f829307cc7bf47801044116ced6d1a3d946bf8aca1008be1cbb66f6d2f331081;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h170d54bf29edffe96aaae0611af495425c64c5ff9ef1b8a418c6a4b506f622b3fea1d4bd2dd878409983cc2824f2ba059219192ca620971e31d8b3596c402025a9b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a4a1937f55626ad228492d8f747f35d5c7b9fe94a46a4a83e4b9ac1620ef8b29a4f52b933e310b07b2a1cc63d0e4c781b5fcfdf9542d1d53c7d505c6f9256e7232b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb41e47d58b07829024f176f22e3546ffb983c24e93f1e98d6e9c926b68a2a6aeb1693d667ef8afbe0f72374f126691149057b96b4a7285c4d150f709a8038573b562;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h111e14e84a15b5c1cd3346a02dd81c6b72749662711bd7e5dd12e4540021f92a7758b1af32a3cff9c214c8624d0c05a4c8180186f785740a23718295df7bb7480da3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc9061e07cb5c14c79c22769a287eb0d77847bd02e4f9b2639d7b9cbb59fc58cc10bc12fd352e4c77fe1017fd9f41b301c34d5a45b3854ae780d82647f953960d2df9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8e5cc64adde86abd61866f25f9c7a3d3982a03a6f67976ce2002e4daca47adfa87dfb235077eb7b25401c61da998a9ae68935170abd779fefd7f0f8148f6d069b37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h134fe8532216217ff506721b7aef6cc9d69c23f2f825fb1763cd5f3a84eae499e4b52661532e955fd08225ff87f64c6ed873e1553f42a2a00f22466f9ecaf0ca20c89;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4b2f624bd069421918208bb53202b7b0916ada0d7aa4405a269d1e89831aa4eaae4f472358a36cab11f6338ddb66aa1c535b978db32bf179810b9b941f6215e878cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h163b6216fb4d3994c43ff2ab008c206bd30b0155532a939c0ade8744322f73bc219145bab64af8743dc0b49752e5f4ad154ae3a24f3183b92f4d7361dd92a69f17fb0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d6a282325b66ec55431ab42ca5254c4f6aed973c2821e4456b83916a7ae7c48da813774663fa78db6ca19f6790b6f3607d3126d6ed7c5d4fe9177ec7a17d4cd106d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b1013ef4223ec0dcbf8edcc3c569793b4b479aed5a7153f49f960cbf4f87fbd3f81a9fd33608482315ac71105063ed1936ce6ceba71b4a5f1b0cb2241b0b62bf6da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f2f50d1606088ecdaf15bd96e06628556f4bb4f23db6273d2934f76be4bab118e2e1620355424f015fd61f9938b7527a0762992433212ac8ccd29c67e07a5d3ef655;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha95190a24e0ae00d925323dd6f8900e8f743e14b1558613ef639f4c7d765bb74584bcf428a48074d44d8d8c680029e02b90ffd4c8d30a41616b6fc4a89c0e3155d4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14c2492f8acf1b6332730bde22cd6dee71d70da762104abc202aa107f592c32d0d08a179fec2b1ca9b6ee90c06b592656f005fb4c288c8ac0e590a16724a251f6ec7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbdb35c24bd57ef617342df19a08a9d29fab3bf22e7fc9b6ce50cfd3607dcfc859878ca1fbd47f8fe446a1bf0349dd737b59a5d396c4151121344acb30a16e939b1e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he06aeb4aef727698699ed0f586342dede0914262d9f1a2d097f918f890e853b4fbf1567733a47e498d537450beef5b46a0c2e46da0bc4aa2fe088d627f596eeaefc4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2fff492b31d77eaf5e5d3523669d403aa315b077ecf9c5781f5711babff8e264d4d53a1f55816a520b464ce4c3ad6321f73ba13c511c22db1d344e7eccd491cf4b13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7b018596d7a0e5e57fbf0f151727a1db9061197b45d5be907d82bf3e14abd281ff6b257524a3a2a76b9d2747ed71a6dcf8adf978559653d93fa8b795c33dadc56f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c22360df0eb18dccbea15e30f415cd4ba6e391c178a47184703d91fefcbd4365ec806396bf156d1a7713cfa93807b065f184c1be85899c0b4c2fde4d1286f58b4143;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h114a2e8610024014b7bf6ed791572f4e2131990dec7865f7f17ddc5d70af0d7064668a865ac49c4f1bd1874407195172294a35566ccd46175d0f3ba45ef42784ec16c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he027eb09e0b0c4fd402e49c6b878c874e2149c8b7fe556a6359f86c83eb54f8695edc24325238548241123a8f9289141402cec09688b8ae6c8aae2ed1974f19a3495;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha233ecf9fb20e8a70a6035fd383114575803477766a5ffb9a5fba719f1cab1116501d4d89e005c43fe6a3511c9a1c77a0f62af692785a87e780753b19c0fd4592ea3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0d7d0acbd815a5d8bc9a410bcb54c236c0c9895af93330cd5298487a485161567de6820f5342abbef37e05b82de4a5048108e1aed668c7039e0c23e3cbf149d7418;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6eaf922034c4984dd0699a486673d810ad8feccc502855286d3375566ca5cb2a3dbc0aa8f66d152b185f3da31110058ef135163999092285cd6f4ab6cdc3ef974418;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b6b8dae780e191b269b878abd6e4c3d9ec1a094fd9de96e2c3f45fd8d48e68f52b03581242c8e84fe08113015fe9750aef74a938737d198eedb022e2c14e73f56a9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc37b4ef0e495adae534ff10ba8314e4e9f55ab2582cdec6677c74787e7e155a155f95ad0ce96fef9c54d5401b80fa980d32bcbceaab56e459170b434754bf756ea7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f780407f05bf28f0c4c8beb63bf4b686c3232308249770b76205f494e5efe2ac1cbc1c9569077f0f06b3fd8de36208143e530972fc04a62ae610d69624a8efa407b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7085b2d62c3e93793473817d5e8c9eed599a1c01916e3493d9dc3141a96e68c3ed434a1fea66a2be8a44e5bcc3ce155e00400e5a2a7847583fbdd0c89d57d2d5cbc1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc5c2df27e816d95a9f8a624e7692a5c3b87f35afff6322fac9666af12de1eede95566bf48fcb85c8d439e5b0cbdd3c083889ad6cb90e0e4392f48f617e8f8945e7aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a285c3a8b2ac7307a6fca06adcefd5462f5833e803c09371db34022e336f451a30eeba1fb1498da2b886953f6cb9903dab8851387b2c2748182df4b3c2deda493c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12757a46c956a6cd92aafd76f3fc5487e95b761658f286a446bbe4af546c121ac94fb338737204bc69cde229d1a17bde56ee5f951e90d66b590cf031b84077700f2d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h187fc8568ef6622fb56726d59cb9976143cc00a4350f481d097fc37af9a06df268dd8ac21fbe22c611ba2f35c2be5fcc708cdb3a7e3ce071675ea578933857d2aabbc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a6722f068c48beae4da81cfce7d3e92d5c1eddae24ab1ea862169d311466b2c877f6f9fc16a6ae6d128b70a3cc452bdfdc163d1d3ce451ac65b290a65cfe10c77c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h82427d84fb20bf8b6fbfe671325e69547b21318026279c7caf04a27ea39c025a599c464a44190a5a5c7a1fbeff1779f45cd2102f829dde8906847469acaadbe34c66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f4c040392834c10132e0d44c326c0c77d48f4f71f8771bef99e9f59d8519a56f21ee32284bdf8e862824f4aba127dfbc3d559d329a7f573dae8cb41fe97c238f7436;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24192aaa57247838a8a5685e1ee32cca060b314e370c1bb6010427f17d0cdd645bc7e81f8566f558797e62e82d4bdcd1496a48c8eaa215c6b30b8a36a51b5bc7e3d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e03adbf6b6d31e3d68d5779f5a1fe57fc1e8ee31e2f8f78f776d6ecd74728eda7a78b55d8f26782d040e9670c3a791141fae7d641d71f3d2543a8c7d35ae2b70b61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a7e49dd36a5ef9ea791fdafe27096840fb35fc0c0042f0419247035b029dcfdaa309a5d6ea3412392b6c15459ad33436584edb39fae1c24e3fd4ef6c479b295a532a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbca51c0420c509d13590c7bcf36ac277598a1d9cbb0538c2c3309376a6dbcf0e5e14dc859cd3cfb6d3088851c2e13db1cd2891f236aa01242c4e9899a479c953b23d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he262f5a937f23168ccd3b1d18063755d64060872f628cb25e6f976d9588c54ed407f3a12d36407359b0e216dbf2410a4f3315014bbb91c56f374992ae7cbd8d50f06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4edde2ae54a9ab7db06d846ffa7e8c226998d8016e65500f1b787d92e78b286acfc98afde13671fd508b22cef1c4448bd36aa2904cc3fca5923f0f8749d2c7b4069a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d9e9e170f71aa52a42323598f080032449e6cca87dea3a1e9827e6b440e67ddcbf5df0d4de3d9a080ddfd458ad0b404f844d7304f88fd71afb131602f1ea1086626;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h573e79097f376fe04c3d40b8b24cd788e136b837b216be8b0e0bd4acb8de1f61c1b6603fc21acd7ba4805f28a10e05670d5202a378ba43f2cedcf85f4778bf57adaf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h51319c761cae0c81c13c29ae9d03f1163f4db8f16f56808be1267b92cb4112c8637ea6ac7563e6fb20778109eb9a1aaf28ad3495c1327b11089b090254edcf2cbe6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a2716696a7aeb12b0f1e64abcfdf00ef09fffae979e09bb6b590f2dc0beb446cf80ded07de82d159d7046a0495b692b6fcbef856b03930cf92a9a3c1a41a81d82a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h140cbf694be9ff2e2939624123cfc1afb41e10dbb7b2310c650c3aa7f0025b833659043436f8d7a35f2c8a010cf8e1fe7d96b7625e4d321a8a84d89a94b163a7db25e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f37bb7cfd1fc910571bbbfb44b26a32df6d1074a4fcd09d07c976531b4e2400dfc6b52f578f77573c114195e77cf1c15b818100ed25b374db9d440ba24d04064bd9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8be1e1e4b8f16715c301904d69262b7aa68cf332a41521b078cf61046620f22bff253603d110525b72612cb3460e56b063b9c2d2d0e9c06a56dcf6ca05b12f16d2c;
        #1
        $finish();
    end
endmodule
